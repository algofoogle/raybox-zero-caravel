VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 589.605 BY 600.325 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 14.320 589.605 14.920 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 357.040 589.605 357.640 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 257.080 589.605 257.680 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 85.720 589.605 86.320 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 100.000 589.605 100.600 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 114.280 589.605 114.880 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 128.560 589.605 129.160 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 142.840 589.605 143.440 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 157.120 589.605 157.720 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 171.400 589.605 172.000 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 185.680 589.605 186.280 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 199.960 589.605 200.560 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 214.240 589.605 214.840 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 228.520 589.605 229.120 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 242.800 589.605 243.400 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 271.360 589.605 271.960 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 285.640 589.605 286.240 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 299.920 589.605 300.520 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 314.200 589.605 314.800 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 328.480 589.605 329.080 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 342.760 589.605 343.360 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 371.320 589.605 371.920 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 385.600 589.605 386.200 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 399.880 589.605 400.480 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 414.160 589.605 414.760 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 428.440 589.605 429.040 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 442.720 589.605 443.320 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 457.000 589.605 457.600 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 471.280 589.605 471.880 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 485.560 589.605 486.160 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 499.840 589.605 500.440 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 514.120 589.605 514.720 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 528.400 589.605 529.000 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 542.680 589.605 543.280 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 556.960 589.605 557.560 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 571.240 589.605 571.840 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 28.600 589.605 29.200 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 42.880 589.605 43.480 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 57.160 589.605 57.760 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 71.440 589.605 72.040 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 585.605 585.520 589.605 586.120 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 596.325 7.730 600.325 ;
    END
  END i_spare_1
  PIN i_test_wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END i_test_wb_clk_i
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 596.325 55.570 600.325 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 596.325 43.610 600.325 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 596.325 31.650 600.325 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 596.325 19.690 600.325 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 596.325 127.330 600.325 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 596.325 115.370 600.325 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 596.325 103.410 600.325 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 596.325 91.450 600.325 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 596.325 79.490 600.325 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 596.325 67.530 600.325 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 596.325 199.090 600.325 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 596.325 175.170 600.325 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 596.325 163.210 600.325 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 596.325 151.250 600.325 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 596.325 139.290 600.325 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 596.325 187.130 600.325 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 596.325 581.810 600.325 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 596.325 462.210 600.325 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 596.325 450.250 600.325 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 596.325 438.290 600.325 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 596.325 426.330 600.325 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 596.325 414.370 600.325 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 596.325 402.410 600.325 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 596.325 569.850 600.325 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 596.325 557.890 600.325 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 596.325 545.930 600.325 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 596.325 533.970 600.325 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 596.325 522.010 600.325 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 596.325 510.050 600.325 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 596.325 498.090 600.325 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 596.325 486.130 600.325 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 596.325 474.170 600.325 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 596.325 390.450 600.325 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 596.325 270.850 600.325 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 596.325 258.890 600.325 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 596.325 246.930 600.325 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 596.325 234.970 600.325 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 596.325 223.010 600.325 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 596.325 211.050 600.325 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 596.325 378.490 600.325 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 596.325 366.530 600.325 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 596.325 354.570 600.325 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 596.325 342.610 600.325 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 596.325 330.650 600.325 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 596.325 318.690 600.325 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 596.325 306.730 600.325 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 596.325 294.770 600.325 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 596.325 282.810 600.325 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 583.930 586.215 ;
        RECT 5.330 577.945 583.930 580.775 ;
        RECT 5.330 572.505 583.930 575.335 ;
        RECT 5.330 567.065 583.930 569.895 ;
        RECT 5.330 561.625 583.930 564.455 ;
        RECT 5.330 556.185 583.930 559.015 ;
        RECT 5.330 550.745 583.930 553.575 ;
        RECT 5.330 545.305 583.930 548.135 ;
        RECT 5.330 539.865 583.930 542.695 ;
        RECT 5.330 534.425 583.930 537.255 ;
        RECT 5.330 528.985 583.930 531.815 ;
        RECT 5.330 523.545 583.930 526.375 ;
        RECT 5.330 518.105 583.930 520.935 ;
        RECT 5.330 512.665 583.930 515.495 ;
        RECT 5.330 507.225 583.930 510.055 ;
        RECT 5.330 501.785 583.930 504.615 ;
        RECT 5.330 496.345 583.930 499.175 ;
        RECT 5.330 490.905 583.930 493.735 ;
        RECT 5.330 485.465 583.930 488.295 ;
        RECT 5.330 480.025 583.930 482.855 ;
        RECT 5.330 474.585 583.930 477.415 ;
        RECT 5.330 469.145 583.930 471.975 ;
        RECT 5.330 463.705 583.930 466.535 ;
        RECT 5.330 458.265 583.930 461.095 ;
        RECT 5.330 452.825 583.930 455.655 ;
        RECT 5.330 447.385 583.930 450.215 ;
        RECT 5.330 441.945 583.930 444.775 ;
        RECT 5.330 436.505 583.930 439.335 ;
        RECT 5.330 431.065 583.930 433.895 ;
        RECT 5.330 425.625 583.930 428.455 ;
        RECT 5.330 420.185 583.930 423.015 ;
        RECT 5.330 414.745 583.930 417.575 ;
        RECT 5.330 409.305 583.930 412.135 ;
        RECT 5.330 403.865 583.930 406.695 ;
        RECT 5.330 398.425 583.930 401.255 ;
        RECT 5.330 392.985 583.930 395.815 ;
        RECT 5.330 387.545 583.930 390.375 ;
        RECT 5.330 382.105 583.930 384.935 ;
        RECT 5.330 376.665 583.930 379.495 ;
        RECT 5.330 371.225 583.930 374.055 ;
        RECT 5.330 365.785 583.930 368.615 ;
        RECT 5.330 360.345 583.930 363.175 ;
        RECT 5.330 354.905 583.930 357.735 ;
        RECT 5.330 349.465 583.930 352.295 ;
        RECT 5.330 344.025 583.930 346.855 ;
        RECT 5.330 338.585 583.930 341.415 ;
        RECT 5.330 333.145 583.930 335.975 ;
        RECT 5.330 327.705 583.930 330.535 ;
        RECT 5.330 322.265 583.930 325.095 ;
        RECT 5.330 316.825 583.930 319.655 ;
        RECT 5.330 311.385 583.930 314.215 ;
        RECT 5.330 305.945 583.930 308.775 ;
        RECT 5.330 300.505 583.930 303.335 ;
        RECT 5.330 295.065 583.930 297.895 ;
        RECT 5.330 289.625 583.930 292.455 ;
        RECT 5.330 284.185 583.930 287.015 ;
        RECT 5.330 278.745 583.930 281.575 ;
        RECT 5.330 273.305 583.930 276.135 ;
        RECT 5.330 267.865 583.930 270.695 ;
        RECT 5.330 262.425 583.930 265.255 ;
        RECT 5.330 256.985 583.930 259.815 ;
        RECT 5.330 251.545 583.930 254.375 ;
        RECT 5.330 246.105 583.930 248.935 ;
        RECT 5.330 240.665 583.930 243.495 ;
        RECT 5.330 235.225 583.930 238.055 ;
        RECT 5.330 229.785 583.930 232.615 ;
        RECT 5.330 224.345 583.930 227.175 ;
        RECT 5.330 218.905 583.930 221.735 ;
        RECT 5.330 213.465 583.930 216.295 ;
        RECT 5.330 208.025 583.930 210.855 ;
        RECT 5.330 202.585 583.930 205.415 ;
        RECT 5.330 197.145 583.930 199.975 ;
        RECT 5.330 191.705 583.930 194.535 ;
        RECT 5.330 186.265 583.930 189.095 ;
        RECT 5.330 180.825 583.930 183.655 ;
        RECT 5.330 175.385 583.930 178.215 ;
        RECT 5.330 169.945 583.930 172.775 ;
        RECT 5.330 164.505 583.930 167.335 ;
        RECT 5.330 159.065 583.930 161.895 ;
        RECT 5.330 153.625 583.930 156.455 ;
        RECT 5.330 148.185 583.930 151.015 ;
        RECT 5.330 142.745 583.930 145.575 ;
        RECT 5.330 137.305 583.930 140.135 ;
        RECT 5.330 131.865 583.930 134.695 ;
        RECT 5.330 126.425 583.930 129.255 ;
        RECT 5.330 120.985 583.930 123.815 ;
        RECT 5.330 115.545 583.930 118.375 ;
        RECT 5.330 110.105 583.930 112.935 ;
        RECT 5.330 104.665 583.930 107.495 ;
        RECT 5.330 99.225 583.930 102.055 ;
        RECT 5.330 93.785 583.930 96.615 ;
        RECT 5.330 88.345 583.930 91.175 ;
        RECT 5.330 82.905 583.930 85.735 ;
        RECT 5.330 77.465 583.930 80.295 ;
        RECT 5.330 72.025 583.930 74.855 ;
        RECT 5.330 66.585 583.930 69.415 ;
        RECT 5.330 61.145 583.930 63.975 ;
        RECT 5.330 55.705 583.930 58.535 ;
        RECT 5.330 50.265 583.930 53.095 ;
        RECT 5.330 44.825 583.930 47.655 ;
        RECT 5.330 39.385 583.930 42.215 ;
        RECT 5.330 33.945 583.930 36.775 ;
        RECT 5.330 28.505 583.930 31.335 ;
        RECT 5.330 23.065 583.930 25.895 ;
        RECT 5.330 17.625 583.930 20.455 ;
        RECT 5.330 12.185 583.930 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 583.740 587.605 ;
      LAYER met1 ;
        RECT 5.520 9.560 583.740 587.760 ;
      LAYER met2 ;
        RECT 8.010 596.045 19.130 596.325 ;
        RECT 19.970 596.045 31.090 596.325 ;
        RECT 31.930 596.045 43.050 596.325 ;
        RECT 43.890 596.045 55.010 596.325 ;
        RECT 55.850 596.045 66.970 596.325 ;
        RECT 67.810 596.045 78.930 596.325 ;
        RECT 79.770 596.045 90.890 596.325 ;
        RECT 91.730 596.045 102.850 596.325 ;
        RECT 103.690 596.045 114.810 596.325 ;
        RECT 115.650 596.045 126.770 596.325 ;
        RECT 127.610 596.045 138.730 596.325 ;
        RECT 139.570 596.045 150.690 596.325 ;
        RECT 151.530 596.045 162.650 596.325 ;
        RECT 163.490 596.045 174.610 596.325 ;
        RECT 175.450 596.045 186.570 596.325 ;
        RECT 187.410 596.045 198.530 596.325 ;
        RECT 199.370 596.045 210.490 596.325 ;
        RECT 211.330 596.045 222.450 596.325 ;
        RECT 223.290 596.045 234.410 596.325 ;
        RECT 235.250 596.045 246.370 596.325 ;
        RECT 247.210 596.045 258.330 596.325 ;
        RECT 259.170 596.045 270.290 596.325 ;
        RECT 271.130 596.045 282.250 596.325 ;
        RECT 283.090 596.045 294.210 596.325 ;
        RECT 295.050 596.045 306.170 596.325 ;
        RECT 307.010 596.045 318.130 596.325 ;
        RECT 318.970 596.045 330.090 596.325 ;
        RECT 330.930 596.045 342.050 596.325 ;
        RECT 342.890 596.045 354.010 596.325 ;
        RECT 354.850 596.045 365.970 596.325 ;
        RECT 366.810 596.045 377.930 596.325 ;
        RECT 378.770 596.045 389.890 596.325 ;
        RECT 390.730 596.045 401.850 596.325 ;
        RECT 402.690 596.045 413.810 596.325 ;
        RECT 414.650 596.045 425.770 596.325 ;
        RECT 426.610 596.045 437.730 596.325 ;
        RECT 438.570 596.045 449.690 596.325 ;
        RECT 450.530 596.045 461.650 596.325 ;
        RECT 462.490 596.045 473.610 596.325 ;
        RECT 474.450 596.045 485.570 596.325 ;
        RECT 486.410 596.045 497.530 596.325 ;
        RECT 498.370 596.045 509.490 596.325 ;
        RECT 510.330 596.045 521.450 596.325 ;
        RECT 522.290 596.045 533.410 596.325 ;
        RECT 534.250 596.045 545.370 596.325 ;
        RECT 546.210 596.045 557.330 596.325 ;
        RECT 558.170 596.045 569.290 596.325 ;
        RECT 570.130 596.045 581.250 596.325 ;
        RECT 582.090 596.045 583.180 596.325 ;
        RECT 7.920 4.280 583.180 596.045 ;
        RECT 7.920 4.000 14.530 4.280 ;
        RECT 15.370 4.000 29.250 4.280 ;
        RECT 30.090 4.000 43.970 4.280 ;
        RECT 44.810 4.000 58.690 4.280 ;
        RECT 59.530 4.000 73.410 4.280 ;
        RECT 74.250 4.000 88.130 4.280 ;
        RECT 88.970 4.000 102.850 4.280 ;
        RECT 103.690 4.000 117.570 4.280 ;
        RECT 118.410 4.000 132.290 4.280 ;
        RECT 133.130 4.000 147.010 4.280 ;
        RECT 147.850 4.000 161.730 4.280 ;
        RECT 162.570 4.000 176.450 4.280 ;
        RECT 177.290 4.000 191.170 4.280 ;
        RECT 192.010 4.000 205.890 4.280 ;
        RECT 206.730 4.000 220.610 4.280 ;
        RECT 221.450 4.000 235.330 4.280 ;
        RECT 236.170 4.000 250.050 4.280 ;
        RECT 250.890 4.000 264.770 4.280 ;
        RECT 265.610 4.000 279.490 4.280 ;
        RECT 280.330 4.000 294.210 4.280 ;
        RECT 295.050 4.000 308.930 4.280 ;
        RECT 309.770 4.000 323.650 4.280 ;
        RECT 324.490 4.000 338.370 4.280 ;
        RECT 339.210 4.000 353.090 4.280 ;
        RECT 353.930 4.000 367.810 4.280 ;
        RECT 368.650 4.000 382.530 4.280 ;
        RECT 383.370 4.000 397.250 4.280 ;
        RECT 398.090 4.000 411.970 4.280 ;
        RECT 412.810 4.000 426.690 4.280 ;
        RECT 427.530 4.000 441.410 4.280 ;
        RECT 442.250 4.000 456.130 4.280 ;
        RECT 456.970 4.000 470.850 4.280 ;
        RECT 471.690 4.000 485.570 4.280 ;
        RECT 486.410 4.000 500.290 4.280 ;
        RECT 501.130 4.000 515.010 4.280 ;
        RECT 515.850 4.000 529.730 4.280 ;
        RECT 530.570 4.000 544.450 4.280 ;
        RECT 545.290 4.000 559.170 4.280 ;
        RECT 560.010 4.000 573.890 4.280 ;
        RECT 574.730 4.000 583.180 4.280 ;
      LAYER met3 ;
        RECT 21.050 586.520 585.605 587.685 ;
        RECT 21.050 585.120 585.205 586.520 ;
        RECT 21.050 572.240 585.605 585.120 ;
        RECT 21.050 570.840 585.205 572.240 ;
        RECT 21.050 557.960 585.605 570.840 ;
        RECT 21.050 556.560 585.205 557.960 ;
        RECT 21.050 543.680 585.605 556.560 ;
        RECT 21.050 542.280 585.205 543.680 ;
        RECT 21.050 529.400 585.605 542.280 ;
        RECT 21.050 528.000 585.205 529.400 ;
        RECT 21.050 515.120 585.605 528.000 ;
        RECT 21.050 513.720 585.205 515.120 ;
        RECT 21.050 500.840 585.605 513.720 ;
        RECT 21.050 499.440 585.205 500.840 ;
        RECT 21.050 486.560 585.605 499.440 ;
        RECT 21.050 485.160 585.205 486.560 ;
        RECT 21.050 472.280 585.605 485.160 ;
        RECT 21.050 470.880 585.205 472.280 ;
        RECT 21.050 458.000 585.605 470.880 ;
        RECT 21.050 456.600 585.205 458.000 ;
        RECT 21.050 443.720 585.605 456.600 ;
        RECT 21.050 442.320 585.205 443.720 ;
        RECT 21.050 429.440 585.605 442.320 ;
        RECT 21.050 428.040 585.205 429.440 ;
        RECT 21.050 415.160 585.605 428.040 ;
        RECT 21.050 413.760 585.205 415.160 ;
        RECT 21.050 400.880 585.605 413.760 ;
        RECT 21.050 399.480 585.205 400.880 ;
        RECT 21.050 386.600 585.605 399.480 ;
        RECT 21.050 385.200 585.205 386.600 ;
        RECT 21.050 372.320 585.605 385.200 ;
        RECT 21.050 370.920 585.205 372.320 ;
        RECT 21.050 358.040 585.605 370.920 ;
        RECT 21.050 356.640 585.205 358.040 ;
        RECT 21.050 343.760 585.605 356.640 ;
        RECT 21.050 342.360 585.205 343.760 ;
        RECT 21.050 329.480 585.605 342.360 ;
        RECT 21.050 328.080 585.205 329.480 ;
        RECT 21.050 315.200 585.605 328.080 ;
        RECT 21.050 313.800 585.205 315.200 ;
        RECT 21.050 300.920 585.605 313.800 ;
        RECT 21.050 299.520 585.205 300.920 ;
        RECT 21.050 286.640 585.605 299.520 ;
        RECT 21.050 285.240 585.205 286.640 ;
        RECT 21.050 272.360 585.605 285.240 ;
        RECT 21.050 270.960 585.205 272.360 ;
        RECT 21.050 258.080 585.605 270.960 ;
        RECT 21.050 256.680 585.205 258.080 ;
        RECT 21.050 243.800 585.605 256.680 ;
        RECT 21.050 242.400 585.205 243.800 ;
        RECT 21.050 229.520 585.605 242.400 ;
        RECT 21.050 228.120 585.205 229.520 ;
        RECT 21.050 215.240 585.605 228.120 ;
        RECT 21.050 213.840 585.205 215.240 ;
        RECT 21.050 200.960 585.605 213.840 ;
        RECT 21.050 199.560 585.205 200.960 ;
        RECT 21.050 186.680 585.605 199.560 ;
        RECT 21.050 185.280 585.205 186.680 ;
        RECT 21.050 172.400 585.605 185.280 ;
        RECT 21.050 171.000 585.205 172.400 ;
        RECT 21.050 158.120 585.605 171.000 ;
        RECT 21.050 156.720 585.205 158.120 ;
        RECT 21.050 143.840 585.605 156.720 ;
        RECT 21.050 142.440 585.205 143.840 ;
        RECT 21.050 129.560 585.605 142.440 ;
        RECT 21.050 128.160 585.205 129.560 ;
        RECT 21.050 115.280 585.605 128.160 ;
        RECT 21.050 113.880 585.205 115.280 ;
        RECT 21.050 101.000 585.605 113.880 ;
        RECT 21.050 99.600 585.205 101.000 ;
        RECT 21.050 86.720 585.605 99.600 ;
        RECT 21.050 85.320 585.205 86.720 ;
        RECT 21.050 72.440 585.605 85.320 ;
        RECT 21.050 71.040 585.205 72.440 ;
        RECT 21.050 58.160 585.605 71.040 ;
        RECT 21.050 56.760 585.205 58.160 ;
        RECT 21.050 43.880 585.605 56.760 ;
        RECT 21.050 42.480 585.205 43.880 ;
        RECT 21.050 29.600 585.605 42.480 ;
        RECT 21.050 28.200 585.205 29.600 ;
        RECT 21.050 15.320 585.605 28.200 ;
        RECT 21.050 13.920 585.205 15.320 ;
        RECT 21.050 9.015 585.605 13.920 ;
      LAYER met4 ;
        RECT 74.815 10.240 97.440 585.305 ;
        RECT 99.840 10.240 174.240 585.305 ;
        RECT 176.640 10.240 251.040 585.305 ;
        RECT 253.440 10.240 327.840 585.305 ;
        RECT 330.240 10.240 404.640 585.305 ;
        RECT 407.040 10.240 481.440 585.305 ;
        RECT 483.840 10.240 523.185 585.305 ;
        RECT 74.815 9.015 523.185 10.240 ;
  END
END top_ew_algofoogle
END LIBRARY

