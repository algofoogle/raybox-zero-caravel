VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 590.535 BY 601.255 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 576.930 597.255 577.210 601.255 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 353.640 590.535 354.240 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 258.440 590.535 259.040 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 95.240 590.535 95.840 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 108.840 590.535 109.440 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 122.440 590.535 123.040 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 136.040 590.535 136.640 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 149.640 590.535 150.240 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 163.240 590.535 163.840 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 176.840 590.535 177.440 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 190.440 590.535 191.040 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 204.040 590.535 204.640 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 217.640 590.535 218.240 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 231.240 590.535 231.840 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 244.840 590.535 245.440 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 272.040 590.535 272.640 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 285.640 590.535 286.240 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 299.240 590.535 299.840 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 312.840 590.535 313.440 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 326.440 590.535 327.040 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 340.040 590.535 340.640 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 367.240 590.535 367.840 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 380.840 590.535 381.440 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 394.440 590.535 395.040 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 408.040 590.535 408.640 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 421.640 590.535 422.240 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 435.240 590.535 435.840 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 448.840 590.535 449.440 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 462.440 590.535 463.040 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 476.040 590.535 476.640 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 489.640 590.535 490.240 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 503.240 590.535 503.840 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 516.840 590.535 517.440 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 530.440 590.535 531.040 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 544.040 590.535 544.640 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 557.640 590.535 558.240 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 40.840 590.535 41.440 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 54.440 590.535 55.040 ;
    END
  END i_reg_mosi
  PIN i_reg_outs_enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 68.040 590.535 68.640 ;
    END
  END i_reg_outs_enb
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 586.535 81.640 590.535 82.240 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END i_reset_lock_b
  PIN i_spare_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 586.535 571.240 590.535 571.840 ;
    END
  END i_spare_0
  PIN i_spare_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 597.255 13.710 601.255 ;
    END
  END i_spare_1
  PIN i_test_uc2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 586.535 27.240 590.535 27.840 ;
    END
  END i_test_uc2
  PIN i_test_wci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END i_test_wci
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 59.430 597.255 59.710 601.255 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 597.255 48.210 601.255 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 36.430 597.255 36.710 601.255 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 597.255 25.210 601.255 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 128.430 597.255 128.710 601.255 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 116.930 597.255 117.210 601.255 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 105.430 597.255 105.710 601.255 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 93.930 597.255 94.210 601.255 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 82.430 597.255 82.710 601.255 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 70.930 597.255 71.210 601.255 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 197.430 597.255 197.710 601.255 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 174.430 597.255 174.710 601.255 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 162.930 597.255 163.210 601.255 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 597.255 151.710 601.255 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 139.930 597.255 140.210 601.255 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 185.930 597.255 186.210 601.255 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 597.255 565.710 601.255 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 597.255 450.710 601.255 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 597.255 439.210 601.255 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 597.255 427.710 601.255 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 597.255 416.210 601.255 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 597.255 404.710 601.255 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 597.255 393.210 601.255 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 597.255 554.210 601.255 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 597.255 542.710 601.255 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 597.255 531.210 601.255 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 597.255 519.710 601.255 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 597.255 508.210 601.255 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 597.255 496.710 601.255 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 597.255 485.210 601.255 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 597.255 473.710 601.255 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 597.255 462.210 601.255 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 590.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 590.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 590.480 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 597.255 381.710 601.255 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 597.255 266.710 601.255 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 597.255 255.210 601.255 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 597.255 243.710 601.255 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 597.255 232.210 601.255 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 597.255 220.710 601.255 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 597.255 209.210 601.255 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 597.255 370.210 601.255 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 597.255 358.710 601.255 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 597.255 347.210 601.255 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 597.255 335.710 601.255 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 597.255 324.210 601.255 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 597.255 312.710 601.255 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 597.255 301.210 601.255 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 597.255 289.710 601.255 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 597.255 278.210 601.255 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 588.825 584.850 590.430 ;
        RECT 5.330 583.385 584.850 586.215 ;
        RECT 5.330 577.945 584.850 580.775 ;
        RECT 5.330 572.505 584.850 575.335 ;
        RECT 5.330 567.065 584.850 569.895 ;
        RECT 5.330 561.625 584.850 564.455 ;
        RECT 5.330 556.185 584.850 559.015 ;
        RECT 5.330 550.745 584.850 553.575 ;
        RECT 5.330 545.305 584.850 548.135 ;
        RECT 5.330 539.865 584.850 542.695 ;
        RECT 5.330 534.425 584.850 537.255 ;
        RECT 5.330 528.985 584.850 531.815 ;
        RECT 5.330 523.545 584.850 526.375 ;
        RECT 5.330 518.105 584.850 520.935 ;
        RECT 5.330 512.665 584.850 515.495 ;
        RECT 5.330 507.225 584.850 510.055 ;
        RECT 5.330 501.785 584.850 504.615 ;
        RECT 5.330 496.345 584.850 499.175 ;
        RECT 5.330 490.905 584.850 493.735 ;
        RECT 5.330 485.465 584.850 488.295 ;
        RECT 5.330 480.025 584.850 482.855 ;
        RECT 5.330 474.585 584.850 477.415 ;
        RECT 5.330 469.145 584.850 471.975 ;
        RECT 5.330 463.705 584.850 466.535 ;
        RECT 5.330 458.265 584.850 461.095 ;
        RECT 5.330 452.825 584.850 455.655 ;
        RECT 5.330 447.385 584.850 450.215 ;
        RECT 5.330 441.945 584.850 444.775 ;
        RECT 5.330 436.505 584.850 439.335 ;
        RECT 5.330 431.065 584.850 433.895 ;
        RECT 5.330 425.625 584.850 428.455 ;
        RECT 5.330 420.185 584.850 423.015 ;
        RECT 5.330 414.745 584.850 417.575 ;
        RECT 5.330 409.305 584.850 412.135 ;
        RECT 5.330 403.865 584.850 406.695 ;
        RECT 5.330 398.425 584.850 401.255 ;
        RECT 5.330 392.985 584.850 395.815 ;
        RECT 5.330 387.545 584.850 390.375 ;
        RECT 5.330 382.105 584.850 384.935 ;
        RECT 5.330 376.665 584.850 379.495 ;
        RECT 5.330 371.225 584.850 374.055 ;
        RECT 5.330 365.785 584.850 368.615 ;
        RECT 5.330 360.345 584.850 363.175 ;
        RECT 5.330 354.905 584.850 357.735 ;
        RECT 5.330 349.465 584.850 352.295 ;
        RECT 5.330 344.025 584.850 346.855 ;
        RECT 5.330 338.585 584.850 341.415 ;
        RECT 5.330 333.145 584.850 335.975 ;
        RECT 5.330 327.705 584.850 330.535 ;
        RECT 5.330 322.265 584.850 325.095 ;
        RECT 5.330 316.825 584.850 319.655 ;
        RECT 5.330 311.385 584.850 314.215 ;
        RECT 5.330 305.945 584.850 308.775 ;
        RECT 5.330 300.505 584.850 303.335 ;
        RECT 5.330 295.065 584.850 297.895 ;
        RECT 5.330 289.625 584.850 292.455 ;
        RECT 5.330 284.185 584.850 287.015 ;
        RECT 5.330 278.745 584.850 281.575 ;
        RECT 5.330 273.305 584.850 276.135 ;
        RECT 5.330 267.865 584.850 270.695 ;
        RECT 5.330 262.425 584.850 265.255 ;
        RECT 5.330 256.985 584.850 259.815 ;
        RECT 5.330 251.545 584.850 254.375 ;
        RECT 5.330 246.105 584.850 248.935 ;
        RECT 5.330 240.665 584.850 243.495 ;
        RECT 5.330 235.225 584.850 238.055 ;
        RECT 5.330 229.785 584.850 232.615 ;
        RECT 5.330 224.345 584.850 227.175 ;
        RECT 5.330 218.905 584.850 221.735 ;
        RECT 5.330 213.465 584.850 216.295 ;
        RECT 5.330 208.025 584.850 210.855 ;
        RECT 5.330 202.585 584.850 205.415 ;
        RECT 5.330 197.145 584.850 199.975 ;
        RECT 5.330 191.705 584.850 194.535 ;
        RECT 5.330 186.265 584.850 189.095 ;
        RECT 5.330 180.825 584.850 183.655 ;
        RECT 5.330 175.385 584.850 178.215 ;
        RECT 5.330 169.945 584.850 172.775 ;
        RECT 5.330 164.505 584.850 167.335 ;
        RECT 5.330 159.065 584.850 161.895 ;
        RECT 5.330 153.625 584.850 156.455 ;
        RECT 5.330 148.185 584.850 151.015 ;
        RECT 5.330 142.745 584.850 145.575 ;
        RECT 5.330 137.305 584.850 140.135 ;
        RECT 5.330 131.865 584.850 134.695 ;
        RECT 5.330 126.425 584.850 129.255 ;
        RECT 5.330 120.985 584.850 123.815 ;
        RECT 5.330 115.545 584.850 118.375 ;
        RECT 5.330 110.105 584.850 112.935 ;
        RECT 5.330 104.665 584.850 107.495 ;
        RECT 5.330 99.225 584.850 102.055 ;
        RECT 5.330 93.785 584.850 96.615 ;
        RECT 5.330 88.345 584.850 91.175 ;
        RECT 5.330 82.905 584.850 85.735 ;
        RECT 5.330 77.465 584.850 80.295 ;
        RECT 5.330 72.025 584.850 74.855 ;
        RECT 5.330 66.585 584.850 69.415 ;
        RECT 5.330 61.145 584.850 63.975 ;
        RECT 5.330 55.705 584.850 58.535 ;
        RECT 5.330 50.265 584.850 53.095 ;
        RECT 5.330 44.825 584.850 47.655 ;
        RECT 5.330 39.385 584.850 42.215 ;
        RECT 5.330 33.945 584.850 36.775 ;
        RECT 5.330 28.505 584.850 31.335 ;
        RECT 5.330 23.065 584.850 25.895 ;
        RECT 5.330 17.625 584.850 20.455 ;
        RECT 5.330 12.185 584.850 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 584.660 590.325 ;
      LAYER met1 ;
        RECT 5.520 10.640 585.970 597.000 ;
      LAYER met2 ;
        RECT 15.280 596.975 24.650 597.450 ;
        RECT 25.490 596.975 36.150 597.450 ;
        RECT 36.990 596.975 47.650 597.450 ;
        RECT 48.490 596.975 59.150 597.450 ;
        RECT 59.990 596.975 70.650 597.450 ;
        RECT 71.490 596.975 82.150 597.450 ;
        RECT 82.990 596.975 93.650 597.450 ;
        RECT 94.490 596.975 105.150 597.450 ;
        RECT 105.990 596.975 116.650 597.450 ;
        RECT 117.490 596.975 128.150 597.450 ;
        RECT 128.990 596.975 139.650 597.450 ;
        RECT 140.490 596.975 151.150 597.450 ;
        RECT 151.990 596.975 162.650 597.450 ;
        RECT 163.490 596.975 174.150 597.450 ;
        RECT 174.990 596.975 185.650 597.450 ;
        RECT 186.490 596.975 197.150 597.450 ;
        RECT 197.990 596.975 208.650 597.450 ;
        RECT 209.490 596.975 220.150 597.450 ;
        RECT 220.990 596.975 231.650 597.450 ;
        RECT 232.490 596.975 243.150 597.450 ;
        RECT 243.990 596.975 254.650 597.450 ;
        RECT 255.490 596.975 266.150 597.450 ;
        RECT 266.990 596.975 277.650 597.450 ;
        RECT 278.490 596.975 289.150 597.450 ;
        RECT 289.990 596.975 300.650 597.450 ;
        RECT 301.490 596.975 312.150 597.450 ;
        RECT 312.990 596.975 323.650 597.450 ;
        RECT 324.490 596.975 335.150 597.450 ;
        RECT 335.990 596.975 346.650 597.450 ;
        RECT 347.490 596.975 358.150 597.450 ;
        RECT 358.990 596.975 369.650 597.450 ;
        RECT 370.490 596.975 381.150 597.450 ;
        RECT 381.990 596.975 392.650 597.450 ;
        RECT 393.490 596.975 404.150 597.450 ;
        RECT 404.990 596.975 415.650 597.450 ;
        RECT 416.490 596.975 427.150 597.450 ;
        RECT 427.990 596.975 438.650 597.450 ;
        RECT 439.490 596.975 450.150 597.450 ;
        RECT 450.990 596.975 461.650 597.450 ;
        RECT 462.490 596.975 473.150 597.450 ;
        RECT 473.990 596.975 484.650 597.450 ;
        RECT 485.490 596.975 496.150 597.450 ;
        RECT 496.990 596.975 507.650 597.450 ;
        RECT 508.490 596.975 519.150 597.450 ;
        RECT 519.990 596.975 530.650 597.450 ;
        RECT 531.490 596.975 542.150 597.450 ;
        RECT 542.990 596.975 553.650 597.450 ;
        RECT 554.490 596.975 565.150 597.450 ;
        RECT 565.990 596.975 576.650 597.450 ;
        RECT 577.490 596.975 585.940 597.450 ;
        RECT 15.280 4.280 585.940 596.975 ;
        RECT 15.830 3.670 29.710 4.280 ;
        RECT 30.550 3.670 44.430 4.280 ;
        RECT 45.270 3.670 59.150 4.280 ;
        RECT 59.990 3.670 73.870 4.280 ;
        RECT 74.710 3.670 88.590 4.280 ;
        RECT 89.430 3.670 103.310 4.280 ;
        RECT 104.150 3.670 118.030 4.280 ;
        RECT 118.870 3.670 132.750 4.280 ;
        RECT 133.590 3.670 147.470 4.280 ;
        RECT 148.310 3.670 162.190 4.280 ;
        RECT 163.030 3.670 176.910 4.280 ;
        RECT 177.750 3.670 191.630 4.280 ;
        RECT 192.470 3.670 206.350 4.280 ;
        RECT 207.190 3.670 221.070 4.280 ;
        RECT 221.910 3.670 235.790 4.280 ;
        RECT 236.630 3.670 250.510 4.280 ;
        RECT 251.350 3.670 265.230 4.280 ;
        RECT 266.070 3.670 279.950 4.280 ;
        RECT 280.790 3.670 294.670 4.280 ;
        RECT 295.510 3.670 309.390 4.280 ;
        RECT 310.230 3.670 324.110 4.280 ;
        RECT 324.950 3.670 338.830 4.280 ;
        RECT 339.670 3.670 353.550 4.280 ;
        RECT 354.390 3.670 368.270 4.280 ;
        RECT 369.110 3.670 382.990 4.280 ;
        RECT 383.830 3.670 397.710 4.280 ;
        RECT 398.550 3.670 412.430 4.280 ;
        RECT 413.270 3.670 427.150 4.280 ;
        RECT 427.990 3.670 441.870 4.280 ;
        RECT 442.710 3.670 456.590 4.280 ;
        RECT 457.430 3.670 471.310 4.280 ;
        RECT 472.150 3.670 486.030 4.280 ;
        RECT 486.870 3.670 500.750 4.280 ;
        RECT 501.590 3.670 515.470 4.280 ;
        RECT 516.310 3.670 530.190 4.280 ;
        RECT 531.030 3.670 544.910 4.280 ;
        RECT 545.750 3.670 559.630 4.280 ;
        RECT 560.470 3.670 574.350 4.280 ;
        RECT 575.190 3.670 585.940 4.280 ;
      LAYER met3 ;
        RECT 21.050 572.240 586.535 591.425 ;
        RECT 21.050 570.840 586.135 572.240 ;
        RECT 21.050 558.640 586.535 570.840 ;
        RECT 21.050 557.240 586.135 558.640 ;
        RECT 21.050 545.040 586.535 557.240 ;
        RECT 21.050 543.640 586.135 545.040 ;
        RECT 21.050 531.440 586.535 543.640 ;
        RECT 21.050 530.040 586.135 531.440 ;
        RECT 21.050 517.840 586.535 530.040 ;
        RECT 21.050 516.440 586.135 517.840 ;
        RECT 21.050 504.240 586.535 516.440 ;
        RECT 21.050 502.840 586.135 504.240 ;
        RECT 21.050 490.640 586.535 502.840 ;
        RECT 21.050 489.240 586.135 490.640 ;
        RECT 21.050 477.040 586.535 489.240 ;
        RECT 21.050 475.640 586.135 477.040 ;
        RECT 21.050 463.440 586.535 475.640 ;
        RECT 21.050 462.040 586.135 463.440 ;
        RECT 21.050 449.840 586.535 462.040 ;
        RECT 21.050 448.440 586.135 449.840 ;
        RECT 21.050 436.240 586.535 448.440 ;
        RECT 21.050 434.840 586.135 436.240 ;
        RECT 21.050 422.640 586.535 434.840 ;
        RECT 21.050 421.240 586.135 422.640 ;
        RECT 21.050 409.040 586.535 421.240 ;
        RECT 21.050 407.640 586.135 409.040 ;
        RECT 21.050 395.440 586.535 407.640 ;
        RECT 21.050 394.040 586.135 395.440 ;
        RECT 21.050 381.840 586.535 394.040 ;
        RECT 21.050 380.440 586.135 381.840 ;
        RECT 21.050 368.240 586.535 380.440 ;
        RECT 21.050 366.840 586.135 368.240 ;
        RECT 21.050 354.640 586.535 366.840 ;
        RECT 21.050 353.240 586.135 354.640 ;
        RECT 21.050 341.040 586.535 353.240 ;
        RECT 21.050 339.640 586.135 341.040 ;
        RECT 21.050 327.440 586.535 339.640 ;
        RECT 21.050 326.040 586.135 327.440 ;
        RECT 21.050 313.840 586.535 326.040 ;
        RECT 21.050 312.440 586.135 313.840 ;
        RECT 21.050 300.240 586.535 312.440 ;
        RECT 21.050 298.840 586.135 300.240 ;
        RECT 21.050 286.640 586.535 298.840 ;
        RECT 21.050 285.240 586.135 286.640 ;
        RECT 21.050 273.040 586.535 285.240 ;
        RECT 21.050 271.640 586.135 273.040 ;
        RECT 21.050 259.440 586.535 271.640 ;
        RECT 21.050 258.040 586.135 259.440 ;
        RECT 21.050 245.840 586.535 258.040 ;
        RECT 21.050 244.440 586.135 245.840 ;
        RECT 21.050 232.240 586.535 244.440 ;
        RECT 21.050 230.840 586.135 232.240 ;
        RECT 21.050 218.640 586.535 230.840 ;
        RECT 21.050 217.240 586.135 218.640 ;
        RECT 21.050 205.040 586.535 217.240 ;
        RECT 21.050 203.640 586.135 205.040 ;
        RECT 21.050 191.440 586.535 203.640 ;
        RECT 21.050 190.040 586.135 191.440 ;
        RECT 21.050 177.840 586.535 190.040 ;
        RECT 21.050 176.440 586.135 177.840 ;
        RECT 21.050 164.240 586.535 176.440 ;
        RECT 21.050 162.840 586.135 164.240 ;
        RECT 21.050 150.640 586.535 162.840 ;
        RECT 21.050 149.240 586.135 150.640 ;
        RECT 21.050 137.040 586.535 149.240 ;
        RECT 21.050 135.640 586.135 137.040 ;
        RECT 21.050 123.440 586.535 135.640 ;
        RECT 21.050 122.040 586.135 123.440 ;
        RECT 21.050 109.840 586.535 122.040 ;
        RECT 21.050 108.440 586.135 109.840 ;
        RECT 21.050 96.240 586.535 108.440 ;
        RECT 21.050 94.840 586.135 96.240 ;
        RECT 21.050 82.640 586.535 94.840 ;
        RECT 21.050 81.240 586.135 82.640 ;
        RECT 21.050 69.040 586.535 81.240 ;
        RECT 21.050 67.640 586.135 69.040 ;
        RECT 21.050 55.440 586.535 67.640 ;
        RECT 21.050 54.040 586.135 55.440 ;
        RECT 21.050 41.840 586.535 54.040 ;
        RECT 21.050 40.440 586.135 41.840 ;
        RECT 21.050 28.240 586.535 40.440 ;
        RECT 21.050 26.840 586.135 28.240 ;
        RECT 21.050 10.715 586.535 26.840 ;
      LAYER met4 ;
        RECT 42.615 13.095 97.440 587.345 ;
        RECT 99.840 13.095 174.240 587.345 ;
        RECT 176.640 13.095 251.040 587.345 ;
        RECT 253.440 13.095 327.840 587.345 ;
        RECT 330.240 13.095 404.640 587.345 ;
        RECT 407.040 13.095 481.440 587.345 ;
        RECT 483.840 13.095 558.240 587.345 ;
        RECT 560.640 13.095 576.545 587.345 ;
  END
END top_ew_algofoogle
END LIBRARY

