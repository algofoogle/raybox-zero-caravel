// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_outs_enb,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_spare_0,
    i_spare_1,
    i_test_wb_clk_i,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_outs_enb;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_spare_0;
 input i_spare_1;
 input i_test_wb_clk_i;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire _00000_;
 wire _00001_;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire clknet_leaf_0_i_clk;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net77;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net78;
 wire net93;
 wire net94;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net111;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdx[5] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_mapdy[5] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.side_hot ;
 wire \rbzero.spi_registers.got_new_floor ;
 wire \rbzero.spi_registers.got_new_leak ;
 wire \rbzero.spi_registers.got_new_mapd ;
 wire \rbzero.spi_registers.got_new_other ;
 wire \rbzero.spi_registers.got_new_sky ;
 wire \rbzero.spi_registers.got_new_texadd[0] ;
 wire \rbzero.spi_registers.got_new_texadd[1] ;
 wire \rbzero.spi_registers.got_new_texadd[2] ;
 wire \rbzero.spi_registers.got_new_texadd[3] ;
 wire \rbzero.spi_registers.got_new_vinf ;
 wire \rbzero.spi_registers.got_new_vshift ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.new_floor[0] ;
 wire \rbzero.spi_registers.new_floor[1] ;
 wire \rbzero.spi_registers.new_floor[2] ;
 wire \rbzero.spi_registers.new_floor[3] ;
 wire \rbzero.spi_registers.new_floor[4] ;
 wire \rbzero.spi_registers.new_floor[5] ;
 wire \rbzero.spi_registers.new_leak[0] ;
 wire \rbzero.spi_registers.new_leak[1] ;
 wire \rbzero.spi_registers.new_leak[2] ;
 wire \rbzero.spi_registers.new_leak[3] ;
 wire \rbzero.spi_registers.new_leak[4] ;
 wire \rbzero.spi_registers.new_leak[5] ;
 wire \rbzero.spi_registers.new_mapd[0] ;
 wire \rbzero.spi_registers.new_mapd[10] ;
 wire \rbzero.spi_registers.new_mapd[11] ;
 wire \rbzero.spi_registers.new_mapd[12] ;
 wire \rbzero.spi_registers.new_mapd[13] ;
 wire \rbzero.spi_registers.new_mapd[14] ;
 wire \rbzero.spi_registers.new_mapd[15] ;
 wire \rbzero.spi_registers.new_mapd[1] ;
 wire \rbzero.spi_registers.new_mapd[2] ;
 wire \rbzero.spi_registers.new_mapd[3] ;
 wire \rbzero.spi_registers.new_mapd[4] ;
 wire \rbzero.spi_registers.new_mapd[5] ;
 wire \rbzero.spi_registers.new_mapd[6] ;
 wire \rbzero.spi_registers.new_mapd[7] ;
 wire \rbzero.spi_registers.new_mapd[8] ;
 wire \rbzero.spi_registers.new_mapd[9] ;
 wire \rbzero.spi_registers.new_other[0] ;
 wire \rbzero.spi_registers.new_other[10] ;
 wire \rbzero.spi_registers.new_other[1] ;
 wire \rbzero.spi_registers.new_other[2] ;
 wire \rbzero.spi_registers.new_other[3] ;
 wire \rbzero.spi_registers.new_other[4] ;
 wire \rbzero.spi_registers.new_other[6] ;
 wire \rbzero.spi_registers.new_other[7] ;
 wire \rbzero.spi_registers.new_other[8] ;
 wire \rbzero.spi_registers.new_other[9] ;
 wire \rbzero.spi_registers.new_sky[0] ;
 wire \rbzero.spi_registers.new_sky[1] ;
 wire \rbzero.spi_registers.new_sky[2] ;
 wire \rbzero.spi_registers.new_sky[3] ;
 wire \rbzero.spi_registers.new_sky[4] ;
 wire \rbzero.spi_registers.new_sky[5] ;
 wire \rbzero.spi_registers.new_texadd[0][0] ;
 wire \rbzero.spi_registers.new_texadd[0][10] ;
 wire \rbzero.spi_registers.new_texadd[0][11] ;
 wire \rbzero.spi_registers.new_texadd[0][12] ;
 wire \rbzero.spi_registers.new_texadd[0][13] ;
 wire \rbzero.spi_registers.new_texadd[0][14] ;
 wire \rbzero.spi_registers.new_texadd[0][15] ;
 wire \rbzero.spi_registers.new_texadd[0][16] ;
 wire \rbzero.spi_registers.new_texadd[0][17] ;
 wire \rbzero.spi_registers.new_texadd[0][18] ;
 wire \rbzero.spi_registers.new_texadd[0][19] ;
 wire \rbzero.spi_registers.new_texadd[0][1] ;
 wire \rbzero.spi_registers.new_texadd[0][20] ;
 wire \rbzero.spi_registers.new_texadd[0][21] ;
 wire \rbzero.spi_registers.new_texadd[0][22] ;
 wire \rbzero.spi_registers.new_texadd[0][23] ;
 wire \rbzero.spi_registers.new_texadd[0][2] ;
 wire \rbzero.spi_registers.new_texadd[0][3] ;
 wire \rbzero.spi_registers.new_texadd[0][4] ;
 wire \rbzero.spi_registers.new_texadd[0][5] ;
 wire \rbzero.spi_registers.new_texadd[0][6] ;
 wire \rbzero.spi_registers.new_texadd[0][7] ;
 wire \rbzero.spi_registers.new_texadd[0][8] ;
 wire \rbzero.spi_registers.new_texadd[0][9] ;
 wire \rbzero.spi_registers.new_texadd[1][0] ;
 wire \rbzero.spi_registers.new_texadd[1][10] ;
 wire \rbzero.spi_registers.new_texadd[1][11] ;
 wire \rbzero.spi_registers.new_texadd[1][12] ;
 wire \rbzero.spi_registers.new_texadd[1][13] ;
 wire \rbzero.spi_registers.new_texadd[1][14] ;
 wire \rbzero.spi_registers.new_texadd[1][15] ;
 wire \rbzero.spi_registers.new_texadd[1][16] ;
 wire \rbzero.spi_registers.new_texadd[1][17] ;
 wire \rbzero.spi_registers.new_texadd[1][18] ;
 wire \rbzero.spi_registers.new_texadd[1][19] ;
 wire \rbzero.spi_registers.new_texadd[1][1] ;
 wire \rbzero.spi_registers.new_texadd[1][20] ;
 wire \rbzero.spi_registers.new_texadd[1][21] ;
 wire \rbzero.spi_registers.new_texadd[1][22] ;
 wire \rbzero.spi_registers.new_texadd[1][23] ;
 wire \rbzero.spi_registers.new_texadd[1][2] ;
 wire \rbzero.spi_registers.new_texadd[1][3] ;
 wire \rbzero.spi_registers.new_texadd[1][4] ;
 wire \rbzero.spi_registers.new_texadd[1][5] ;
 wire \rbzero.spi_registers.new_texadd[1][6] ;
 wire \rbzero.spi_registers.new_texadd[1][7] ;
 wire \rbzero.spi_registers.new_texadd[1][8] ;
 wire \rbzero.spi_registers.new_texadd[1][9] ;
 wire \rbzero.spi_registers.new_texadd[2][0] ;
 wire \rbzero.spi_registers.new_texadd[2][10] ;
 wire \rbzero.spi_registers.new_texadd[2][11] ;
 wire \rbzero.spi_registers.new_texadd[2][12] ;
 wire \rbzero.spi_registers.new_texadd[2][13] ;
 wire \rbzero.spi_registers.new_texadd[2][14] ;
 wire \rbzero.spi_registers.new_texadd[2][15] ;
 wire \rbzero.spi_registers.new_texadd[2][16] ;
 wire \rbzero.spi_registers.new_texadd[2][17] ;
 wire \rbzero.spi_registers.new_texadd[2][18] ;
 wire \rbzero.spi_registers.new_texadd[2][19] ;
 wire \rbzero.spi_registers.new_texadd[2][1] ;
 wire \rbzero.spi_registers.new_texadd[2][20] ;
 wire \rbzero.spi_registers.new_texadd[2][21] ;
 wire \rbzero.spi_registers.new_texadd[2][22] ;
 wire \rbzero.spi_registers.new_texadd[2][23] ;
 wire \rbzero.spi_registers.new_texadd[2][2] ;
 wire \rbzero.spi_registers.new_texadd[2][3] ;
 wire \rbzero.spi_registers.new_texadd[2][4] ;
 wire \rbzero.spi_registers.new_texadd[2][5] ;
 wire \rbzero.spi_registers.new_texadd[2][6] ;
 wire \rbzero.spi_registers.new_texadd[2][7] ;
 wire \rbzero.spi_registers.new_texadd[2][8] ;
 wire \rbzero.spi_registers.new_texadd[2][9] ;
 wire \rbzero.spi_registers.new_texadd[3][0] ;
 wire \rbzero.spi_registers.new_texadd[3][10] ;
 wire \rbzero.spi_registers.new_texadd[3][11] ;
 wire \rbzero.spi_registers.new_texadd[3][12] ;
 wire \rbzero.spi_registers.new_texadd[3][13] ;
 wire \rbzero.spi_registers.new_texadd[3][14] ;
 wire \rbzero.spi_registers.new_texadd[3][15] ;
 wire \rbzero.spi_registers.new_texadd[3][16] ;
 wire \rbzero.spi_registers.new_texadd[3][17] ;
 wire \rbzero.spi_registers.new_texadd[3][18] ;
 wire \rbzero.spi_registers.new_texadd[3][19] ;
 wire \rbzero.spi_registers.new_texadd[3][1] ;
 wire \rbzero.spi_registers.new_texadd[3][20] ;
 wire \rbzero.spi_registers.new_texadd[3][21] ;
 wire \rbzero.spi_registers.new_texadd[3][22] ;
 wire \rbzero.spi_registers.new_texadd[3][23] ;
 wire \rbzero.spi_registers.new_texadd[3][2] ;
 wire \rbzero.spi_registers.new_texadd[3][3] ;
 wire \rbzero.spi_registers.new_texadd[3][4] ;
 wire \rbzero.spi_registers.new_texadd[3][5] ;
 wire \rbzero.spi_registers.new_texadd[3][6] ;
 wire \rbzero.spi_registers.new_texadd[3][7] ;
 wire \rbzero.spi_registers.new_texadd[3][8] ;
 wire \rbzero.spi_registers.new_texadd[3][9] ;
 wire \rbzero.spi_registers.new_vinf ;
 wire \rbzero.spi_registers.new_vshift[0] ;
 wire \rbzero.spi_registers.new_vshift[1] ;
 wire \rbzero.spi_registers.new_vshift[2] ;
 wire \rbzero.spi_registers.new_vshift[3] ;
 wire \rbzero.spi_registers.new_vshift[4] ;
 wire \rbzero.spi_registers.new_vshift[5] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[16] ;
 wire \rbzero.spi_registers.spi_buffer[17] ;
 wire \rbzero.spi_registers.spi_buffer[18] ;
 wire \rbzero.spi_registers.spi_buffer[19] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[20] ;
 wire \rbzero.spi_registers.spi_buffer[21] ;
 wire \rbzero.spi_registers.spi_buffer[22] ;
 wire \rbzero.spi_registers.spi_buffer[23] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.texadd0[0] ;
 wire \rbzero.spi_registers.texadd0[10] ;
 wire \rbzero.spi_registers.texadd0[11] ;
 wire \rbzero.spi_registers.texadd0[12] ;
 wire \rbzero.spi_registers.texadd0[13] ;
 wire \rbzero.spi_registers.texadd0[14] ;
 wire \rbzero.spi_registers.texadd0[15] ;
 wire \rbzero.spi_registers.texadd0[16] ;
 wire \rbzero.spi_registers.texadd0[17] ;
 wire \rbzero.spi_registers.texadd0[18] ;
 wire \rbzero.spi_registers.texadd0[19] ;
 wire \rbzero.spi_registers.texadd0[1] ;
 wire \rbzero.spi_registers.texadd0[20] ;
 wire \rbzero.spi_registers.texadd0[21] ;
 wire \rbzero.spi_registers.texadd0[22] ;
 wire \rbzero.spi_registers.texadd0[23] ;
 wire \rbzero.spi_registers.texadd0[2] ;
 wire \rbzero.spi_registers.texadd0[3] ;
 wire \rbzero.spi_registers.texadd0[4] ;
 wire \rbzero.spi_registers.texadd0[5] ;
 wire \rbzero.spi_registers.texadd0[6] ;
 wire \rbzero.spi_registers.texadd0[7] ;
 wire \rbzero.spi_registers.texadd0[8] ;
 wire \rbzero.spi_registers.texadd0[9] ;
 wire \rbzero.spi_registers.texadd1[0] ;
 wire \rbzero.spi_registers.texadd1[10] ;
 wire \rbzero.spi_registers.texadd1[11] ;
 wire \rbzero.spi_registers.texadd1[12] ;
 wire \rbzero.spi_registers.texadd1[13] ;
 wire \rbzero.spi_registers.texadd1[14] ;
 wire \rbzero.spi_registers.texadd1[15] ;
 wire \rbzero.spi_registers.texadd1[16] ;
 wire \rbzero.spi_registers.texadd1[17] ;
 wire \rbzero.spi_registers.texadd1[18] ;
 wire \rbzero.spi_registers.texadd1[19] ;
 wire \rbzero.spi_registers.texadd1[1] ;
 wire \rbzero.spi_registers.texadd1[20] ;
 wire \rbzero.spi_registers.texadd1[21] ;
 wire \rbzero.spi_registers.texadd1[22] ;
 wire \rbzero.spi_registers.texadd1[23] ;
 wire \rbzero.spi_registers.texadd1[2] ;
 wire \rbzero.spi_registers.texadd1[3] ;
 wire \rbzero.spi_registers.texadd1[4] ;
 wire \rbzero.spi_registers.texadd1[5] ;
 wire \rbzero.spi_registers.texadd1[6] ;
 wire \rbzero.spi_registers.texadd1[7] ;
 wire \rbzero.spi_registers.texadd1[8] ;
 wire \rbzero.spi_registers.texadd1[9] ;
 wire \rbzero.spi_registers.texadd2[0] ;
 wire \rbzero.spi_registers.texadd2[10] ;
 wire \rbzero.spi_registers.texadd2[11] ;
 wire \rbzero.spi_registers.texadd2[12] ;
 wire \rbzero.spi_registers.texadd2[13] ;
 wire \rbzero.spi_registers.texadd2[14] ;
 wire \rbzero.spi_registers.texadd2[15] ;
 wire \rbzero.spi_registers.texadd2[16] ;
 wire \rbzero.spi_registers.texadd2[17] ;
 wire \rbzero.spi_registers.texadd2[18] ;
 wire \rbzero.spi_registers.texadd2[19] ;
 wire \rbzero.spi_registers.texadd2[1] ;
 wire \rbzero.spi_registers.texadd2[20] ;
 wire \rbzero.spi_registers.texadd2[21] ;
 wire \rbzero.spi_registers.texadd2[22] ;
 wire \rbzero.spi_registers.texadd2[23] ;
 wire \rbzero.spi_registers.texadd2[2] ;
 wire \rbzero.spi_registers.texadd2[3] ;
 wire \rbzero.spi_registers.texadd2[4] ;
 wire \rbzero.spi_registers.texadd2[5] ;
 wire \rbzero.spi_registers.texadd2[6] ;
 wire \rbzero.spi_registers.texadd2[7] ;
 wire \rbzero.spi_registers.texadd2[8] ;
 wire \rbzero.spi_registers.texadd2[9] ;
 wire \rbzero.spi_registers.texadd3[0] ;
 wire \rbzero.spi_registers.texadd3[10] ;
 wire \rbzero.spi_registers.texadd3[11] ;
 wire \rbzero.spi_registers.texadd3[12] ;
 wire \rbzero.spi_registers.texadd3[13] ;
 wire \rbzero.spi_registers.texadd3[14] ;
 wire \rbzero.spi_registers.texadd3[15] ;
 wire \rbzero.spi_registers.texadd3[16] ;
 wire \rbzero.spi_registers.texadd3[17] ;
 wire \rbzero.spi_registers.texadd3[18] ;
 wire \rbzero.spi_registers.texadd3[19] ;
 wire \rbzero.spi_registers.texadd3[1] ;
 wire \rbzero.spi_registers.texadd3[20] ;
 wire \rbzero.spi_registers.texadd3[21] ;
 wire \rbzero.spi_registers.texadd3[22] ;
 wire \rbzero.spi_registers.texadd3[23] ;
 wire \rbzero.spi_registers.texadd3[2] ;
 wire \rbzero.spi_registers.texadd3[3] ;
 wire \rbzero.spi_registers.texadd3[4] ;
 wire \rbzero.spi_registers.texadd3[5] ;
 wire \rbzero.spi_registers.texadd3[6] ;
 wire \rbzero.spi_registers.texadd3[7] ;
 wire \rbzero.spi_registers.texadd3[8] ;
 wire \rbzero.spi_registers.texadd3[9] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.texu_hot[0] ;
 wire \rbzero.texu_hot[1] ;
 wire \rbzero.texu_hot[2] ;
 wire \rbzero.texu_hot[3] ;
 wire \rbzero.texu_hot[4] ;
 wire \rbzero.texu_hot[5] ;
 wire \rbzero.trace_state[0] ;
 wire \rbzero.trace_state[1] ;
 wire \rbzero.trace_state[2] ;
 wire \rbzero.trace_state[3] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_hot[0] ;
 wire \rbzero.wall_hot[1] ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \reg_gpout[0] ;
 wire \reg_gpout[1] ;
 wire \reg_gpout[2] ;
 wire \reg_gpout[3] ;
 wire \reg_gpout[4] ;
 wire \reg_gpout[5] ;
 wire reg_hsync;
 wire \reg_rgb[14] ;
 wire \reg_rgb[15] ;
 wire \reg_rgb[22] ;
 wire \reg_rgb[23] ;
 wire \reg_rgb[6] ;
 wire \reg_rgb[7] ;
 wire reg_vsync;
 wire net95;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net129;
 wire net75;
 wire net76;
 wire net127;
 wire net128;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_101_i_clk;
 wire clknet_leaf_102_i_clk;
 wire clknet_leaf_103_i_clk;
 wire clknet_leaf_104_i_clk;
 wire clknet_leaf_105_i_clk;
 wire clknet_leaf_106_i_clk;
 wire clknet_leaf_107_i_clk;
 wire clknet_leaf_108_i_clk;
 wire clknet_leaf_110_i_clk;
 wire clknet_leaf_111_i_clk;
 wire clknet_leaf_112_i_clk;
 wire clknet_leaf_113_i_clk;
 wire clknet_leaf_114_i_clk;
 wire clknet_leaf_115_i_clk;
 wire clknet_leaf_116_i_clk;
 wire clknet_leaf_117_i_clk;
 wire clknet_leaf_118_i_clk;
 wire clknet_leaf_119_i_clk;
 wire clknet_leaf_120_i_clk;
 wire clknet_leaf_121_i_clk;
 wire clknet_leaf_122_i_clk;
 wire clknet_leaf_123_i_clk;
 wire clknet_leaf_124_i_clk;
 wire clknet_leaf_125_i_clk;
 wire clknet_leaf_126_i_clk;
 wire clknet_leaf_127_i_clk;
 wire clknet_leaf_128_i_clk;
 wire clknet_leaf_129_i_clk;
 wire clknet_leaf_130_i_clk;
 wire clknet_leaf_131_i_clk;
 wire clknet_leaf_132_i_clk;
 wire clknet_leaf_133_i_clk;
 wire clknet_leaf_134_i_clk;
 wire clknet_leaf_135_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_0_1_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_1_1_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_2_1_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_2_3_1_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_4_0_0_i_clk;
 wire clknet_4_1_0_i_clk;
 wire clknet_4_2_0_i_clk;
 wire clknet_4_3_0_i_clk;
 wire clknet_4_4_0_i_clk;
 wire clknet_4_5_0_i_clk;
 wire clknet_4_6_0_i_clk;
 wire clknet_4_7_0_i_clk;
 wire clknet_4_8_0_i_clk;
 wire clknet_4_9_0_i_clk;
 wire clknet_4_10_0_i_clk;
 wire clknet_4_11_0_i_clk;
 wire clknet_4_12_0_i_clk;
 wire clknet_4_13_0_i_clk;
 wire clknet_4_14_0_i_clk;
 wire clknet_4_15_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_opt_2_0_i_clk;
 wire clknet_opt_3_0_i_clk;
 wire clknet_opt_3_1_i_clk;
 wire clknet_opt_4_0_i_clk;
 wire clknet_opt_5_0_i_clk;
 wire clknet_opt_6_0_i_clk;
 wire clknet_0__05775_;
 wire clknet_1_0__leaf__05775_;
 wire clknet_1_1__leaf__05775_;
 wire clknet_0__06050_;
 wire clknet_1_0__leaf__06050_;
 wire clknet_1_1__leaf__06050_;
 wire clknet_0__05825_;
 wire clknet_1_0__leaf__05825_;
 wire clknet_1_1__leaf__05825_;
 wire clknet_0__03869_;
 wire clknet_1_0__leaf__03869_;
 wire clknet_1_1__leaf__03869_;
 wire clknet_0__03868_;
 wire clknet_1_0__leaf__03868_;
 wire clknet_1_1__leaf__03868_;
 wire clknet_0__03857_;
 wire clknet_1_0__leaf__03857_;
 wire clknet_1_1__leaf__03857_;
 wire clknet_0__03867_;
 wire clknet_1_0__leaf__03867_;
 wire clknet_1_1__leaf__03867_;
 wire clknet_0__03866_;
 wire clknet_1_0__leaf__03866_;
 wire clknet_1_1__leaf__03866_;
 wire clknet_0__03865_;
 wire clknet_1_0__leaf__03865_;
 wire clknet_1_1__leaf__03865_;
 wire clknet_0__03864_;
 wire clknet_1_0__leaf__03864_;
 wire clknet_1_1__leaf__03864_;
 wire clknet_0__03863_;
 wire clknet_1_0__leaf__03863_;
 wire clknet_1_1__leaf__03863_;
 wire clknet_0__03862_;
 wire clknet_1_0__leaf__03862_;
 wire clknet_1_1__leaf__03862_;
 wire clknet_0__03861_;
 wire clknet_1_0__leaf__03861_;
 wire clknet_1_1__leaf__03861_;
 wire clknet_0__03860_;
 wire clknet_1_0__leaf__03860_;
 wire clknet_1_1__leaf__03860_;
 wire clknet_0__03859_;
 wire clknet_1_0__leaf__03859_;
 wire clknet_1_1__leaf__03859_;
 wire clknet_0__03858_;
 wire clknet_1_0__leaf__03858_;
 wire clknet_1_1__leaf__03858_;
 wire clknet_0__03846_;
 wire clknet_1_0__leaf__03846_;
 wire clknet_1_1__leaf__03846_;
 wire clknet_0__03856_;
 wire clknet_1_0__leaf__03856_;
 wire clknet_1_1__leaf__03856_;
 wire clknet_0__03855_;
 wire clknet_1_0__leaf__03855_;
 wire clknet_1_1__leaf__03855_;
 wire clknet_0__03854_;
 wire clknet_1_0__leaf__03854_;
 wire clknet_1_1__leaf__03854_;
 wire clknet_0__03853_;
 wire clknet_1_0__leaf__03853_;
 wire clknet_1_1__leaf__03853_;
 wire clknet_0__03852_;
 wire clknet_1_0__leaf__03852_;
 wire clknet_1_1__leaf__03852_;
 wire clknet_0__03851_;
 wire clknet_1_0__leaf__03851_;
 wire clknet_1_1__leaf__03851_;
 wire clknet_0__03850_;
 wire clknet_1_0__leaf__03850_;
 wire clknet_1_1__leaf__03850_;
 wire clknet_0__03849_;
 wire clknet_1_0__leaf__03849_;
 wire clknet_1_1__leaf__03849_;
 wire clknet_0__03848_;
 wire clknet_1_0__leaf__03848_;
 wire clknet_1_1__leaf__03848_;
 wire clknet_0__03847_;
 wire clknet_1_0__leaf__03847_;
 wire clknet_1_1__leaf__03847_;
 wire clknet_0__03510_;
 wire clknet_1_0__leaf__03510_;
 wire clknet_1_1__leaf__03510_;
 wire clknet_0__03845_;
 wire clknet_1_0__leaf__03845_;
 wire clknet_1_1__leaf__03845_;
 wire clknet_0__03844_;
 wire clknet_1_0__leaf__03844_;
 wire clknet_1_1__leaf__03844_;
 wire clknet_0__03843_;
 wire clknet_1_0__leaf__03843_;
 wire clknet_1_1__leaf__03843_;
 wire clknet_0__03842_;
 wire clknet_1_0__leaf__03842_;
 wire clknet_1_1__leaf__03842_;
 wire clknet_0__03841_;
 wire clknet_1_0__leaf__03841_;
 wire clknet_1_1__leaf__03841_;
 wire clknet_0__03840_;
 wire clknet_1_0__leaf__03840_;
 wire clknet_1_1__leaf__03840_;
 wire clknet_0__03839_;
 wire clknet_1_0__leaf__03839_;
 wire clknet_1_1__leaf__03839_;
 wire clknet_0__03838_;
 wire clknet_1_0__leaf__03838_;
 wire clknet_1_1__leaf__03838_;
 wire clknet_0__03837_;
 wire clknet_1_0__leaf__03837_;
 wire clknet_1_1__leaf__03837_;
 wire clknet_0__03511_;
 wire clknet_1_0__leaf__03511_;
 wire clknet_1_1__leaf__03511_;
 wire clknet_0__03503_;
 wire clknet_1_0__leaf__03503_;
 wire clknet_1_1__leaf__03503_;
 wire clknet_0__03509_;
 wire clknet_1_0__leaf__03509_;
 wire clknet_1_1__leaf__03509_;
 wire clknet_0__03508_;
 wire clknet_1_0__leaf__03508_;
 wire clknet_1_1__leaf__03508_;
 wire clknet_0__03507_;
 wire clknet_1_0__leaf__03507_;
 wire clknet_1_1__leaf__03507_;
 wire clknet_0__03506_;
 wire clknet_1_0__leaf__03506_;
 wire clknet_1_1__leaf__03506_;
 wire clknet_0__03505_;
 wire clknet_1_0__leaf__03505_;
 wire clknet_1_1__leaf__03505_;
 wire clknet_0__03504_;
 wire clknet_1_0__leaf__03504_;
 wire clknet_1_1__leaf__03504_;
 wire clknet_0__06001_;
 wire clknet_1_0__leaf__06001_;
 wire clknet_1_1__leaf__06001_;
 wire clknet_0__05942_;
 wire clknet_1_0__leaf__05942_;
 wire clknet_1_1__leaf__05942_;
 wire clknet_0__05887_;
 wire clknet_1_0__leaf__05887_;
 wire clknet_1_1__leaf__05887_;
 wire clknet_0__05832_;
 wire clknet_1_0__leaf__05832_;
 wire clknet_1_1__leaf__05832_;
 wire net74;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;

 sky130_fd_sc_hd__buf_4 _10448_ (.A(\gpout0.hpos[0] ),
    .X(_04029_));
 sky130_fd_sc_hd__buf_4 _10449_ (.A(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__buf_4 _10450_ (.A(\gpout0.hpos[7] ),
    .X(_04031_));
 sky130_fd_sc_hd__clkbuf_4 _10451_ (.A(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__clkbuf_4 _10452_ (.A(\gpout0.hpos[8] ),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_4 _10453_ (.A(\gpout0.hpos[9] ),
    .X(_04034_));
 sky130_fd_sc_hd__nor2b_2 _10454_ (.A(_04033_),
    .B_N(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__xor2_4 _10455_ (.A(net47),
    .B(net48),
    .X(_04036_));
 sky130_fd_sc_hd__and4_2 _10456_ (.A(_04030_),
    .B(_04032_),
    .C(_04035_),
    .D(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__buf_4 _10457_ (.A(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_4 _10458_ (.A(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(\rbzero.tex_r1[63] ),
    .A1(net50),
    .S(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_1 _10460_ (.A(_04040_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[63] ),
    .S(_04039_),
    .X(_04041_));
 sky130_fd_sc_hd__clkbuf_1 _10462_ (.A(_04041_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_04039_),
    .X(_04042_));
 sky130_fd_sc_hd__clkbuf_1 _10464_ (.A(_04042_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(_04039_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_1 _10466_ (.A(_04043_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_04039_),
    .X(_04044_));
 sky130_fd_sc_hd__clkbuf_1 _10468_ (.A(_04044_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_04039_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _10470_ (.A(_04045_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_04039_),
    .X(_04046_));
 sky130_fd_sc_hd__clkbuf_1 _10472_ (.A(_04046_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _10473_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(_04039_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_1 _10474_ (.A(_04047_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_04039_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_1 _10476_ (.A(_04048_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(_04039_),
    .X(_04049_));
 sky130_fd_sc_hd__clkbuf_1 _10478_ (.A(_04049_),
    .X(_01588_));
 sky130_fd_sc_hd__clkbuf_4 _10479_ (.A(_04038_),
    .X(_04050_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__clkbuf_1 _10481_ (.A(_04051_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _10482_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(_04050_),
    .X(_04052_));
 sky130_fd_sc_hd__clkbuf_1 _10483_ (.A(_04052_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_04050_),
    .X(_04053_));
 sky130_fd_sc_hd__clkbuf_1 _10485_ (.A(_04053_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _10486_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_04050_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_1 _10487_ (.A(_04054_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_04050_),
    .X(_04055_));
 sky130_fd_sc_hd__clkbuf_1 _10489_ (.A(_04055_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(_04050_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_1 _10491_ (.A(_04056_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_04050_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_1 _10493_ (.A(_04057_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(_04050_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _10495_ (.A(_04058_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_04050_),
    .X(_04059_));
 sky130_fd_sc_hd__clkbuf_1 _10497_ (.A(_04059_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(_04050_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _10499_ (.A(_04060_),
    .X(_01578_));
 sky130_fd_sc_hd__clkbuf_4 _10500_ (.A(_04038_),
    .X(_04061_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(_04062_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _10503_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(_04061_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _10504_ (.A(_04063_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_04061_),
    .X(_04064_));
 sky130_fd_sc_hd__clkbuf_1 _10506_ (.A(_04064_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(_04061_),
    .X(_04065_));
 sky130_fd_sc_hd__clkbuf_1 _10508_ (.A(_04065_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(\rbzero.tex_r1[39] ),
    .A1(net74),
    .S(_04061_),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _10510_ (.A(_04066_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(_04061_),
    .X(_04067_));
 sky130_fd_sc_hd__clkbuf_1 _10512_ (.A(_04067_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04061_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_1 _10514_ (.A(_04068_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_04061_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _10516_ (.A(_04069_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_04061_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_1 _10518_ (.A(_04070_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(_04061_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _10520_ (.A(_04071_),
    .X(_01568_));
 sky130_fd_sc_hd__clkbuf_4 _10521_ (.A(_04038_),
    .X(_04072_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__clkbuf_1 _10523_ (.A(_04073_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _10524_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(_04072_),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _10525_ (.A(_04074_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_04072_),
    .X(_04075_));
 sky130_fd_sc_hd__clkbuf_1 _10527_ (.A(_04075_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(_04072_),
    .X(_04076_));
 sky130_fd_sc_hd__clkbuf_1 _10529_ (.A(_04076_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_04072_),
    .X(_04077_));
 sky130_fd_sc_hd__clkbuf_1 _10531_ (.A(_04077_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(_04072_),
    .X(_04078_));
 sky130_fd_sc_hd__clkbuf_1 _10533_ (.A(_04078_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_04072_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _10535_ (.A(_04079_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _10536_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(_04072_),
    .X(_04080_));
 sky130_fd_sc_hd__clkbuf_1 _10537_ (.A(_04080_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_04072_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_1 _10539_ (.A(_04081_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _10540_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(_04072_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _10541_ (.A(_04082_),
    .X(_01558_));
 sky130_fd_sc_hd__clkbuf_4 _10542_ (.A(_04038_),
    .X(_04083_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__clkbuf_1 _10544_ (.A(_04084_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _10545_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(_04083_),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _10546_ (.A(_04085_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _10547_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_04083_),
    .X(_04086_));
 sky130_fd_sc_hd__clkbuf_1 _10548_ (.A(_04086_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _10549_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(_04083_),
    .X(_04087_));
 sky130_fd_sc_hd__clkbuf_1 _10550_ (.A(_04087_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_04083_),
    .X(_04088_));
 sky130_fd_sc_hd__clkbuf_1 _10552_ (.A(_04088_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(_04083_),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_1 _10554_ (.A(_04089_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_04083_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_1 _10556_ (.A(_04090_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _10557_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(_04083_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _10558_ (.A(_04091_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _10559_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_04083_),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _10560_ (.A(_04092_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _10561_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(_04083_),
    .X(_04093_));
 sky130_fd_sc_hd__clkbuf_1 _10562_ (.A(_04093_),
    .X(_01548_));
 sky130_fd_sc_hd__clkbuf_4 _10563_ (.A(_04038_),
    .X(_04094_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_04094_),
    .X(_04095_));
 sky130_fd_sc_hd__clkbuf_1 _10565_ (.A(_04095_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_04094_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _10567_ (.A(_04096_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_04094_),
    .X(_04097_));
 sky130_fd_sc_hd__clkbuf_1 _10569_ (.A(_04097_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(_04094_),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _10571_ (.A(_04098_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_04094_),
    .X(_04099_));
 sky130_fd_sc_hd__clkbuf_1 _10573_ (.A(_04099_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_04094_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _10575_ (.A(_04100_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04094_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_1 _10577_ (.A(_04101_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10578_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(_04094_),
    .X(_04102_));
 sky130_fd_sc_hd__clkbuf_1 _10579_ (.A(_04102_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10580_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04094_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _10581_ (.A(_04103_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(_04094_),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_1 _10583_ (.A(_04104_),
    .X(_01538_));
 sky130_fd_sc_hd__clkbuf_4 _10584_ (.A(_04038_),
    .X(_04105_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _10586_ (.A(_04106_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _10587_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_04105_),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _10588_ (.A(_04107_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_04105_),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_1 _10590_ (.A(_04108_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10591_ (.A0(\rbzero.tex_r1[0] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(_04105_),
    .X(_04109_));
 sky130_fd_sc_hd__clkbuf_1 _10592_ (.A(_04109_),
    .X(_01534_));
 sky130_fd_sc_hd__inv_2 _10593_ (.A(\gpout0.hpos[0] ),
    .Y(_04110_));
 sky130_fd_sc_hd__buf_4 _10594_ (.A(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__buf_6 _10595_ (.A(_04036_),
    .X(_04112_));
 sky130_fd_sc_hd__nand4_4 _10596_ (.A(_04111_),
    .B(_04032_),
    .C(_04035_),
    .D(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__buf_4 _10597_ (.A(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_4 _10598_ (.A(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(net50),
    .A1(\rbzero.tex_r0[63] ),
    .S(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _10600_ (.A(_04116_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04115_),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_04117_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_04115_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(_04118_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04115_),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_04119_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(_04115_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(_04120_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04115_),
    .X(_04121_));
 sky130_fd_sc_hd__clkbuf_1 _10610_ (.A(_04121_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(_04115_),
    .X(_04122_));
 sky130_fd_sc_hd__clkbuf_1 _10612_ (.A(_04122_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04115_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_04123_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(_04115_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _10616_ (.A(_04124_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10617_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04115_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _10618_ (.A(_04125_),
    .X(_01524_));
 sky130_fd_sc_hd__clkbuf_4 _10619_ (.A(_04114_),
    .X(_04126_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__clkbuf_1 _10621_ (.A(_04127_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04126_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_04128_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_04126_),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_04129_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_04126_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(_04130_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(_04126_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_04131_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04126_),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _10631_ (.A(_04132_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(_04126_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_04133_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04126_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _10635_ (.A(_04134_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_04126_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_1 _10637_ (.A(_04135_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04126_),
    .X(_04136_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_04136_),
    .X(_01514_));
 sky130_fd_sc_hd__clkbuf_4 _10640_ (.A(_04114_),
    .X(_04137_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__clkbuf_1 _10642_ (.A(_04138_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04137_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(_04139_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(_04137_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(_04140_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04137_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(_04141_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(_04137_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(_04142_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04137_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _10652_ (.A(_04143_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(_04137_),
    .X(_04144_));
 sky130_fd_sc_hd__clkbuf_1 _10654_ (.A(_04144_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04137_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _10656_ (.A(_04145_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(_04137_),
    .X(_04146_));
 sky130_fd_sc_hd__clkbuf_1 _10658_ (.A(_04146_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04137_),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _10660_ (.A(_04147_),
    .X(_01504_));
 sky130_fd_sc_hd__clkbuf_4 _10661_ (.A(_04114_),
    .X(_04148_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(_04149_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04148_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(_04150_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(_04148_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(_04151_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04148_),
    .X(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(_04152_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(_04148_),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(_04153_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04148_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _10673_ (.A(_04154_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_04148_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_04155_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04148_),
    .X(_04156_));
 sky130_fd_sc_hd__clkbuf_1 _10677_ (.A(_04156_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(_04148_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_04157_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04148_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_04158_),
    .X(_01494_));
 sky130_fd_sc_hd__clkbuf_4 _10682_ (.A(_04114_),
    .X(_04159_));
 sky130_fd_sc_hd__mux2_1 _10683_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _10684_ (.A(_04160_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04159_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _10686_ (.A(_04161_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(_04159_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10688_ (.A(_04162_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04159_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _10690_ (.A(_04163_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(_04159_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _10692_ (.A(_04164_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10693_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04159_),
    .X(_04165_));
 sky130_fd_sc_hd__clkbuf_1 _10694_ (.A(_04165_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(_04159_),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_1 _10696_ (.A(_04166_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04159_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _10698_ (.A(_04167_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(_04159_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(_04168_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04159_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _10702_ (.A(_04169_),
    .X(_01484_));
 sky130_fd_sc_hd__clkbuf_4 _10703_ (.A(_04114_),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _10705_ (.A(_04171_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04170_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(_04172_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(_04170_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(_04173_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04170_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(_04174_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_04170_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(_04175_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04170_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _10715_ (.A(_04176_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(_04170_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _10717_ (.A(_04177_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04170_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _10719_ (.A(_04178_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(_04170_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_04179_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04170_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _10723_ (.A(_04180_),
    .X(_01474_));
 sky130_fd_sc_hd__buf_4 _10724_ (.A(_04114_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(_04182_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_04181_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(_04183_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10729_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_04181_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(_04184_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10731_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04181_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_1 _10732_ (.A(_04185_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(\rbzero.tex_g1[63] ),
    .A1(net51),
    .S(_04105_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _10734_ (.A(_04186_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10735_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[63] ),
    .S(_04105_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _10736_ (.A(_04187_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_04105_),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _10738_ (.A(_04188_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10739_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(_04105_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _10740_ (.A(_04189_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04105_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _10742_ (.A(_04190_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_04105_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _10744_ (.A(_04191_),
    .X(_01464_));
 sky130_fd_sc_hd__clkbuf_4 _10745_ (.A(_04038_),
    .X(_04192_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _10747_ (.A(_04193_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(_04192_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _10749_ (.A(_04194_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_04192_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _10751_ (.A(_04195_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(_04192_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(_04196_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_04192_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _10755_ (.A(_04197_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(_04192_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _10757_ (.A(_04198_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04192_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_04199_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(_04192_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_04200_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04192_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_04201_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_04192_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_04202_),
    .X(_01454_));
 sky130_fd_sc_hd__buf_4 _10766_ (.A(_04037_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_4 _10767_ (.A(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_04205_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(_04204_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _10771_ (.A(_04206_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_04204_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _10773_ (.A(_04207_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(_04204_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _10775_ (.A(_04208_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_04204_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _10777_ (.A(_04209_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10778_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(_04204_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _10779_ (.A(_04210_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10780_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_04204_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10781_ (.A(_04211_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10782_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_04204_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _10783_ (.A(_04212_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _10784_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_04204_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _10785_ (.A(_04213_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10786_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(_04204_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _10787_ (.A(_04214_),
    .X(_01444_));
 sky130_fd_sc_hd__clkbuf_4 _10788_ (.A(_04203_),
    .X(_04215_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(_04216_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(_04215_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_04217_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_04215_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _10794_ (.A(_04218_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(_04215_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_04219_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_04215_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _10798_ (.A(_04220_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(_04215_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _10800_ (.A(_04221_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10801_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_04215_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _10802_ (.A(_04222_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(_04215_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _10804_ (.A(_04223_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10805_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_04215_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _10806_ (.A(_04224_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(_04215_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _10808_ (.A(_04225_),
    .X(_01434_));
 sky130_fd_sc_hd__clkbuf_4 _10809_ (.A(_04203_),
    .X(_04226_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(_04227_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(_04226_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(_04228_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_04226_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _10815_ (.A(_04229_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(_04226_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_04230_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04226_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _10819_ (.A(_04231_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10820_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(_04226_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _10821_ (.A(_04232_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10822_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_04226_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _10823_ (.A(_04233_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(_04226_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _10825_ (.A(_04234_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10826_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04226_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _10827_ (.A(_04235_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(_04226_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _10829_ (.A(_04236_),
    .X(_01424_));
 sky130_fd_sc_hd__clkbuf_4 _10830_ (.A(_04203_),
    .X(_04237_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(_04238_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(_04237_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_04239_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_04237_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(_04240_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(_04237_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(_04241_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_04237_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(_04242_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _10841_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(_04237_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _10842_ (.A(_04243_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_04237_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _10844_ (.A(_04244_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(_04237_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _10846_ (.A(_04245_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_04237_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _10848_ (.A(_04246_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(_04237_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_04247_),
    .X(_01414_));
 sky130_fd_sc_hd__buf_4 _10851_ (.A(_04203_),
    .X(_04248_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _10853_ (.A(_04249_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(_04248_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _10855_ (.A(_04250_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10856_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_04248_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _10857_ (.A(_04251_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10858_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(_04248_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _10859_ (.A(_04252_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10860_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_04248_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _10861_ (.A(_04253_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(_04248_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _10863_ (.A(_04254_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_04248_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _10865_ (.A(_04255_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(\rbzero.tex_g1[0] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_04248_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(_04256_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(net51),
    .A1(\rbzero.tex_g0[63] ),
    .S(_04181_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(_04257_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_04181_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _10871_ (.A(_04258_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(_04181_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_04259_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04181_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(_04260_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_04181_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(_04261_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04181_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_04262_),
    .X(_01400_));
 sky130_fd_sc_hd__clkbuf_4 _10880_ (.A(_04114_),
    .X(_04263_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _10882_ (.A(_04264_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_04263_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _10884_ (.A(_04265_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(_04263_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(_04266_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04263_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_04267_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(_04263_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_04268_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_04263_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_04269_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(_04263_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_04270_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_04263_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(_04271_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(_04263_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_04272_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04263_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_04273_),
    .X(_01390_));
 sky130_fd_sc_hd__buf_4 _10901_ (.A(_04113_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_4 _10902_ (.A(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_04276_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04275_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(_04277_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(_04275_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_04278_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_04275_),
    .X(_04279_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_04279_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(_04275_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_04280_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04275_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(_04281_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _10915_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_04275_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _10916_ (.A(_04282_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _10917_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04275_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _10918_ (.A(_04283_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _10919_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(_04275_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _10920_ (.A(_04284_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04275_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _10922_ (.A(_04285_),
    .X(_01380_));
 sky130_fd_sc_hd__clkbuf_4 _10923_ (.A(_04274_),
    .X(_04286_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_04287_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04286_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(_04288_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(_04286_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_04289_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04286_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _10931_ (.A(_04290_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(_04286_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _10933_ (.A(_04291_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _10934_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04286_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _10935_ (.A(_04292_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(_04286_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _10937_ (.A(_04293_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_04286_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _10939_ (.A(_04294_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _10940_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(_04286_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _10941_ (.A(_04295_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _10942_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04286_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _10943_ (.A(_04296_),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_4 _10944_ (.A(_04274_),
    .X(_04297_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(_04298_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_04297_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_04299_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(_04297_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_04300_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_04297_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _10952_ (.A(_04301_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _10953_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(_04297_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _10954_ (.A(_04302_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04297_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _10956_ (.A(_04303_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(_04297_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _10958_ (.A(_04304_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _10959_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04297_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _10960_ (.A(_04305_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(_04297_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _10962_ (.A(_04306_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _10963_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_04297_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _10964_ (.A(_04307_),
    .X(_01360_));
 sky130_fd_sc_hd__clkbuf_4 _10965_ (.A(_04274_),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _10967_ (.A(_04309_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04308_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_04310_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(_04308_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(_04311_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_04308_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(_04312_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(_04308_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _10975_ (.A(_04313_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _10976_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04308_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _10977_ (.A(_04314_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _10978_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_04308_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _10979_ (.A(_04315_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _10980_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_04308_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _10981_ (.A(_04316_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(_04308_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _10983_ (.A(_04317_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04308_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(_04318_),
    .X(_01350_));
 sky130_fd_sc_hd__buf_4 _10986_ (.A(_04274_),
    .X(_04319_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _10988_ (.A(_04320_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04319_),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_1 _10990_ (.A(_04321_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(_04319_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _10992_ (.A(_04322_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04319_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _10994_ (.A(_04323_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(_04319_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _10996_ (.A(_04324_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_04319_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _10998_ (.A(_04325_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_04319_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _11000_ (.A(_04326_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_04319_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _11002_ (.A(_04327_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\rbzero.tex_b1[63] ),
    .A1(net52),
    .S(_04248_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(_04328_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[63] ),
    .S(_04248_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_04329_),
    .X(_01340_));
 sky130_fd_sc_hd__clkbuf_4 _11007_ (.A(_04203_),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_1 _11008_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _11009_ (.A(_04331_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _11010_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(_04330_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_1 _11011_ (.A(_04332_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04330_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _11013_ (.A(_04333_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(_04330_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _11015_ (.A(_04334_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_04330_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _11017_ (.A(_04335_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(_04330_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _11019_ (.A(_04336_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_04330_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _11021_ (.A(_04337_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(_04330_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _11023_ (.A(_04338_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04330_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _11025_ (.A(_04339_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(_04330_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _11027_ (.A(_04340_),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_4 _11028_ (.A(_04203_),
    .X(_04341_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _11030_ (.A(_04342_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(_04341_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _11032_ (.A(_04343_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04341_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _11034_ (.A(_04344_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(_04341_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _11036_ (.A(_04345_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04341_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _11038_ (.A(_04346_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(_04341_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _11040_ (.A(_04347_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04341_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _11042_ (.A(_04348_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(_04341_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _11044_ (.A(_04349_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_04341_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _11046_ (.A(_04350_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(_04341_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_04351_),
    .X(_01320_));
 sky130_fd_sc_hd__clkbuf_4 _11049_ (.A(_04203_),
    .X(_04352_));
 sky130_fd_sc_hd__mux2_1 _11050_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _11051_ (.A(_04353_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(_04352_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _11053_ (.A(_04354_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_04352_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(_04355_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(_04352_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _11057_ (.A(_04356_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04352_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _11059_ (.A(_04357_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(_04352_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(_04358_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_04352_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(_04359_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(_04352_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(_04360_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_04352_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(_04361_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(_04352_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(_04362_),
    .X(_01310_));
 sky130_fd_sc_hd__clkbuf_4 _11070_ (.A(_04203_),
    .X(_04363_));
 sky130_fd_sc_hd__mux2_1 _11071_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _11072_ (.A(_04364_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(_04363_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _11074_ (.A(_04365_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_04363_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _11076_ (.A(_04366_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_04363_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _11078_ (.A(_04367_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_04363_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _11080_ (.A(_04368_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(_04363_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _11082_ (.A(_04369_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_04363_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_1 _11084_ (.A(_04370_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(_04363_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _11086_ (.A(_04371_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_04363_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _11088_ (.A(_04372_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_04363_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _11090_ (.A(_04373_),
    .X(_01300_));
 sky130_fd_sc_hd__clkbuf_4 _11091_ (.A(_04203_),
    .X(_04374_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _11093_ (.A(_04375_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(_04374_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(_04376_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04374_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(_04377_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(_04374_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(_04378_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_04374_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(_04379_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(_04374_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _11103_ (.A(_04380_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04374_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _11105_ (.A(_04381_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_04374_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _11107_ (.A(_04382_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04374_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _11109_ (.A(_04383_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(_04374_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _11111_ (.A(_04384_),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_4 _11112_ (.A(_04037_),
    .X(_04385_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _11114_ (.A(_04386_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(_04385_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(_04387_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04385_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(_04388_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_04385_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _11120_ (.A(_04389_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04385_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _11122_ (.A(_04390_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _11123_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(_04385_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _11124_ (.A(_04391_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04385_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _11126_ (.A(_04392_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_04385_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _11128_ (.A(_04393_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04385_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(_04394_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _11131_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_04385_),
    .X(_04395_));
 sky130_fd_sc_hd__clkbuf_1 _11132_ (.A(_04395_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _11133_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_04038_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _11134_ (.A(_04396_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _11135_ (.A0(\rbzero.tex_b1[0] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_04038_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _11136_ (.A(_04397_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _11137_ (.A0(net52),
    .A1(\rbzero.tex_b0[63] ),
    .S(_04319_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _11138_ (.A(_04398_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _11139_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_04319_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _11140_ (.A(_04399_),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_4 _11141_ (.A(_04274_),
    .X(_04400_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(_04401_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _11144_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_04400_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _11145_ (.A(_04402_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(_04400_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _11147_ (.A(_04403_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_04400_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _11149_ (.A(_04404_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(_04400_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _11151_ (.A(_04405_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_04400_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _11153_ (.A(_04406_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(_04400_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(_04407_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_04400_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _11157_ (.A(_04408_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _11158_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(_04400_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _11159_ (.A(_04409_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_04400_),
    .X(_04410_));
 sky130_fd_sc_hd__clkbuf_1 _11161_ (.A(_04410_),
    .X(_01074_));
 sky130_fd_sc_hd__clkbuf_4 _11162_ (.A(_04274_),
    .X(_04411_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(_04411_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(_04412_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04411_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _11166_ (.A(_04413_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(_04411_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _11168_ (.A(_04414_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_04411_),
    .X(_04415_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(_04415_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(_04411_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(_04416_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_04411_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _11174_ (.A(_04417_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_04411_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _11176_ (.A(_04418_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _11177_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_04411_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _11178_ (.A(_04419_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _11179_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_04411_),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_1 _11180_ (.A(_04420_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _11181_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_04411_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_1 _11182_ (.A(_04421_),
    .X(_01064_));
 sky130_fd_sc_hd__clkbuf_4 _11183_ (.A(_04274_),
    .X(_04422_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(_04423_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_04422_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _11187_ (.A(_04424_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(_04422_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(_04425_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_04422_),
    .X(_04426_));
 sky130_fd_sc_hd__clkbuf_1 _11191_ (.A(_04426_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(_04422_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _11193_ (.A(_04427_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04422_),
    .X(_04428_));
 sky130_fd_sc_hd__clkbuf_1 _11195_ (.A(_04428_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _11196_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_04422_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _11197_ (.A(_04429_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_04422_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _11199_ (.A(_04430_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(_04422_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _11201_ (.A(_04431_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _11202_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_04422_),
    .X(_04432_));
 sky130_fd_sc_hd__clkbuf_1 _11203_ (.A(_04432_),
    .X(_01054_));
 sky130_fd_sc_hd__clkbuf_4 _11204_ (.A(_04274_),
    .X(_04433_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__clkbuf_1 _11206_ (.A(_04434_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_04433_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(_04435_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(_04433_),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(_04436_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_04433_),
    .X(_04437_));
 sky130_fd_sc_hd__clkbuf_1 _11212_ (.A(_04437_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(_04433_),
    .X(_04438_));
 sky130_fd_sc_hd__clkbuf_1 _11214_ (.A(_04438_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _11215_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_04433_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _11216_ (.A(_04439_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(_04433_),
    .X(_04440_));
 sky130_fd_sc_hd__clkbuf_1 _11218_ (.A(_04440_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04433_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _11220_ (.A(_04441_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _11221_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(_04433_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _11222_ (.A(_04442_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _11223_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_04433_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _11224_ (.A(_04443_),
    .X(_01044_));
 sky130_fd_sc_hd__clkbuf_4 _11225_ (.A(_04274_),
    .X(_04444_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _11227_ (.A(_04445_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04444_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _11229_ (.A(_04446_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _11230_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(_04444_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _11231_ (.A(_04447_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_04444_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _11233_ (.A(_04448_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(_04444_),
    .X(_04449_));
 sky130_fd_sc_hd__clkbuf_1 _11235_ (.A(_04449_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04444_),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _11237_ (.A(_04450_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(_04444_),
    .X(_04451_));
 sky130_fd_sc_hd__clkbuf_1 _11239_ (.A(_04451_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_04444_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _11241_ (.A(_04452_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _11242_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_04444_),
    .X(_04453_));
 sky130_fd_sc_hd__clkbuf_1 _11243_ (.A(_04453_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_04444_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _11245_ (.A(_04454_),
    .X(_01034_));
 sky130_fd_sc_hd__clkbuf_4 _11246_ (.A(_04113_),
    .X(_04455_));
 sky130_fd_sc_hd__mux2_1 _11247_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _11248_ (.A(_04456_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_04455_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _11250_ (.A(_04457_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(_04455_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _11252_ (.A(_04458_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _11253_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_04455_),
    .X(_04459_));
 sky130_fd_sc_hd__clkbuf_1 _11254_ (.A(_04459_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(_04455_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _11256_ (.A(_04460_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _11257_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_04455_),
    .X(_04461_));
 sky130_fd_sc_hd__clkbuf_1 _11258_ (.A(_04461_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(_04455_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _11260_ (.A(_04462_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _11261_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04455_),
    .X(_04463_));
 sky130_fd_sc_hd__clkbuf_1 _11262_ (.A(_04463_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _11263_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(_04455_),
    .X(_04464_));
 sky130_fd_sc_hd__clkbuf_1 _11264_ (.A(_04464_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _11265_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_04455_),
    .X(_04465_));
 sky130_fd_sc_hd__clkbuf_1 _11266_ (.A(_04465_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _11267_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_04114_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_1 _11268_ (.A(_04466_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _11269_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04114_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _11270_ (.A(_04467_),
    .X(_01022_));
 sky130_fd_sc_hd__clkinv_4 _11271_ (.A(_04036_),
    .Y(_04468_));
 sky130_fd_sc_hd__buf_6 _11272_ (.A(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__buf_4 _11273_ (.A(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__buf_6 _11274_ (.A(_04470_),
    .X(net64));
 sky130_fd_sc_hd__buf_2 _11275_ (.A(\gpout0.hpos[3] ),
    .X(_04471_));
 sky130_fd_sc_hd__and3_1 _11276_ (.A(_04471_),
    .B(\gpout0.hpos[5] ),
    .C(\gpout0.hpos[4] ),
    .X(_04472_));
 sky130_fd_sc_hd__buf_2 _11277_ (.A(\gpout0.hpos[5] ),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_4 _11278_ (.A(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__inv_2 _11279_ (.A(\gpout0.hpos[3] ),
    .Y(_04475_));
 sky130_fd_sc_hd__buf_4 _11280_ (.A(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__clkinv_4 _11281_ (.A(\gpout0.hpos[4] ),
    .Y(_04477_));
 sky130_fd_sc_hd__nor2_2 _11282_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__buf_2 _11283_ (.A(\gpout0.hpos[6] ),
    .X(_04479_));
 sky130_fd_sc_hd__buf_4 _11284_ (.A(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__buf_2 _11285_ (.A(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__o21ai_1 _11286_ (.A1(_04474_),
    .A2(_04478_),
    .B1(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__or4b_1 _11287_ (.A(_04032_),
    .B(_04472_),
    .C(_04482_),
    .D_N(_04035_),
    .X(_04483_));
 sky130_fd_sc_hd__buf_6 _11288_ (.A(_04483_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 _11289_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_04484_));
 sky130_fd_sc_hd__buf_2 _11290_ (.A(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__buf_4 _11291_ (.A(\rbzero.trace_state[2] ),
    .X(_04486_));
 sky130_fd_sc_hd__or2_2 _11292_ (.A(\rbzero.trace_state[1] ),
    .B(\rbzero.trace_state[0] ),
    .X(_04487_));
 sky130_fd_sc_hd__clkinv_2 _11293_ (.A(\rbzero.vga_sync.vsync ),
    .Y(_04488_));
 sky130_fd_sc_hd__nand2_8 _11294_ (.A(_04488_),
    .B(_04036_),
    .Y(_04489_));
 sky130_fd_sc_hd__inv_2 _11295_ (.A(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__buf_4 _11296_ (.A(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__o31a_1 _11297_ (.A1(\rbzero.trace_state[3] ),
    .A2(_04486_),
    .A3(_04487_),
    .B1(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__buf_4 _11298_ (.A(\rbzero.trace_state[1] ),
    .X(_04493_));
 sky130_fd_sc_hd__buf_4 _11299_ (.A(\rbzero.trace_state[0] ),
    .X(_04494_));
 sky130_fd_sc_hd__buf_2 _11300_ (.A(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__nor2_1 _11301_ (.A(\rbzero.trace_state[3] ),
    .B(_04486_),
    .Y(_04496_));
 sky130_fd_sc_hd__and3_1 _11302_ (.A(_04493_),
    .B(_04495_),
    .C(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__and4bb_1 _11303_ (.A_N(_04486_),
    .B_N(_04493_),
    .C(_04495_),
    .D(\rbzero.trace_state[3] ),
    .X(_04498_));
 sky130_fd_sc_hd__nor2_1 _11304_ (.A(_04497_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__buf_4 _11305_ (.A(_04491_),
    .X(_04500_));
 sky130_fd_sc_hd__a32o_1 _11306_ (.A1(_04485_),
    .A2(_04492_),
    .A3(_04499_),
    .B1(_04497_),
    .B2(_04500_),
    .X(_00001_));
 sky130_fd_sc_hd__inv_2 _11307_ (.A(\gpout0.hpos[7] ),
    .Y(_04501_));
 sky130_fd_sc_hd__a21bo_2 _11308_ (.A1(_04501_),
    .A2(_04482_),
    .B1_N(_04035_),
    .X(net71));
 sky130_fd_sc_hd__buf_2 _11309_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_04502_));
 sky130_fd_sc_hd__buf_2 _11310_ (.A(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__buf_2 _11311_ (.A(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__a21bo_1 _11312_ (.A1(_04504_),
    .A2(_04499_),
    .B1_N(_04492_),
    .X(_00000_));
 sky130_fd_sc_hd__inv_2 _11313_ (.A(net72),
    .Y(_04505_));
 sky130_fd_sc_hd__clkbuf_4 _11314_ (.A(\gpout0.hpos[2] ),
    .X(_04506_));
 sky130_fd_sc_hd__buf_4 _11315_ (.A(\gpout0.hpos[1] ),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_4 _11316_ (.A(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__or2_1 _11317_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .X(_04509_));
 sky130_fd_sc_hd__or2_2 _11318_ (.A(\gpout0.hpos[2] ),
    .B(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__o21ai_1 _11319_ (.A1(_04506_),
    .A2(_04508_),
    .B1(_04030_),
    .Y(_04511_));
 sky130_fd_sc_hd__a22o_1 _11320_ (.A1(_04506_),
    .A2(_04508_),
    .B1(_04510_),
    .B2(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__buf_4 _11321_ (.A(_04471_),
    .X(_04513_));
 sky130_fd_sc_hd__clkinv_4 _11322_ (.A(\gpout0.hpos[6] ),
    .Y(_04514_));
 sky130_fd_sc_hd__clkinv_2 _11323_ (.A(\rbzero.wall_hot[1] ),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _11324_ (.A(_04515_),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04516_));
 sky130_fd_sc_hd__clkbuf_4 _11325_ (.A(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__buf_4 _11326_ (.A(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__inv_2 _11327_ (.A(\rbzero.wall_hot[0] ),
    .Y(_04519_));
 sky130_fd_sc_hd__nor2_1 _11328_ (.A(_04515_),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__clkbuf_4 _11329_ (.A(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_4 _11330_ (.A(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__nor2_1 _11331_ (.A(_04515_),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04523_));
 sky130_fd_sc_hd__clkbuf_4 _11332_ (.A(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__clkbuf_4 _11333_ (.A(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__clkbuf_4 _11334_ (.A(\rbzero.wall_hot[0] ),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_4 _11335_ (.A(_04515_),
    .X(_04527_));
 sky130_fd_sc_hd__o21a_1 _11336_ (.A1(\rbzero.spi_registers.texadd3[19] ),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__a221o_1 _11337_ (.A1(\rbzero.spi_registers.texadd2[19] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[19] ),
    .C1(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__o21a_1 _11338_ (.A1(\rbzero.spi_registers.texadd0[19] ),
    .A2(_04518_),
    .B1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__and3_1 _11339_ (.A(\rbzero.spi_registers.texadd2[14] ),
    .B(\rbzero.wall_hot[1] ),
    .C(_04526_),
    .X(_04531_));
 sky130_fd_sc_hd__a31o_1 _11340_ (.A1(\rbzero.spi_registers.texadd3[14] ),
    .A2(_04527_),
    .A3(_04519_),
    .B1(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__or2_1 _11341_ (.A(\rbzero.spi_registers.texadd3[13] ),
    .B(\rbzero.wall_hot[1] ),
    .X(_04533_));
 sky130_fd_sc_hd__o211a_1 _11342_ (.A1(\rbzero.spi_registers.texadd1[13] ),
    .A2(_04527_),
    .B1(_04519_),
    .C1(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_4 _11343_ (.A(\rbzero.side_hot ),
    .X(_04535_));
 sky130_fd_sc_hd__buf_4 _11344_ (.A(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__o21a_1 _11345_ (.A1(\rbzero.spi_registers.texadd3[12] ),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04537_));
 sky130_fd_sc_hd__a221o_1 _11346_ (.A1(\rbzero.spi_registers.texadd2[12] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[12] ),
    .C1(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__o21a_1 _11347_ (.A1(\rbzero.spi_registers.texadd0[12] ),
    .A2(_04517_),
    .B1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__and2_1 _11348_ (.A(_04536_),
    .B(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__nor2_1 _11349_ (.A(_04536_),
    .B(_04539_),
    .Y(_04541_));
 sky130_fd_sc_hd__or2_1 _11350_ (.A(_04540_),
    .B(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__o21a_1 _11351_ (.A1(\rbzero.spi_registers.texadd3[11] ),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04543_));
 sky130_fd_sc_hd__a221o_1 _11352_ (.A1(\rbzero.spi_registers.texadd2[11] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[11] ),
    .C1(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__o21a_1 _11353_ (.A1(\rbzero.spi_registers.texadd0[11] ),
    .A2(_04517_),
    .B1(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__xnor2_1 _11354_ (.A(\rbzero.texu_hot[5] ),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__o21a_1 _11355_ (.A1(\rbzero.spi_registers.texadd3[10] ),
    .A2(_04526_),
    .B1(_04515_),
    .X(_04547_));
 sky130_fd_sc_hd__a221o_1 _11356_ (.A1(\rbzero.spi_registers.texadd2[10] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[10] ),
    .C1(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__o21a_1 _11357_ (.A1(\rbzero.spi_registers.texadd0[10] ),
    .A2(_04517_),
    .B1(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__xnor2_1 _11358_ (.A(\rbzero.texu_hot[4] ),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__o21a_1 _11359_ (.A1(\rbzero.spi_registers.texadd3[9] ),
    .A2(\rbzero.wall_hot[0] ),
    .B1(_04515_),
    .X(_04551_));
 sky130_fd_sc_hd__a221o_1 _11360_ (.A1(\rbzero.spi_registers.texadd2[9] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[9] ),
    .C1(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__o21a_1 _11361_ (.A1(\rbzero.spi_registers.texadd0[9] ),
    .A2(_04517_),
    .B1(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__o21a_1 _11362_ (.A1(\rbzero.spi_registers.texadd3[8] ),
    .A2(\rbzero.wall_hot[0] ),
    .B1(_04515_),
    .X(_04554_));
 sky130_fd_sc_hd__a221o_1 _11363_ (.A1(\rbzero.spi_registers.texadd2[8] ),
    .A2(_04520_),
    .B1(_04523_),
    .B2(\rbzero.spi_registers.texadd1[8] ),
    .C1(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__o21a_1 _11364_ (.A1(\rbzero.spi_registers.texadd0[8] ),
    .A2(_04517_),
    .B1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__nand2_1 _11365_ (.A(\rbzero.texu_hot[2] ),
    .B(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__or2_1 _11366_ (.A(\rbzero.texu_hot[2] ),
    .B(_04556_),
    .X(_04558_));
 sky130_fd_sc_hd__and2_1 _11367_ (.A(_04557_),
    .B(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__o21a_1 _11368_ (.A1(\rbzero.spi_registers.texadd3[7] ),
    .A2(\rbzero.wall_hot[0] ),
    .B1(_04515_),
    .X(_04560_));
 sky130_fd_sc_hd__a221o_1 _11369_ (.A1(\rbzero.spi_registers.texadd2[7] ),
    .A2(_04520_),
    .B1(_04523_),
    .B2(\rbzero.spi_registers.texadd1[7] ),
    .C1(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__o21a_1 _11370_ (.A1(\rbzero.spi_registers.texadd0[7] ),
    .A2(_04516_),
    .B1(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__o21a_1 _11371_ (.A1(\rbzero.spi_registers.texadd3[6] ),
    .A2(\rbzero.wall_hot[0] ),
    .B1(_04515_),
    .X(_04563_));
 sky130_fd_sc_hd__a221o_1 _11372_ (.A1(\rbzero.spi_registers.texadd2[6] ),
    .A2(_04521_),
    .B1(_04523_),
    .B2(\rbzero.spi_registers.texadd1[6] ),
    .C1(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__or2_1 _11373_ (.A(\rbzero.spi_registers.texadd0[6] ),
    .B(_04516_),
    .X(_04565_));
 sky130_fd_sc_hd__nand3_1 _11374_ (.A(\rbzero.texu_hot[0] ),
    .B(_04564_),
    .C(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__xnor2_1 _11375_ (.A(\rbzero.texu_hot[1] ),
    .B(_04562_),
    .Y(_04567_));
 sky130_fd_sc_hd__nor2_1 _11376_ (.A(_04566_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__a21o_1 _11377_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_04562_),
    .B1(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__nand2_1 _11378_ (.A(_04559_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__xnor2_1 _11379_ (.A(\rbzero.texu_hot[3] ),
    .B(_04553_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21oi_1 _11380_ (.A1(_04557_),
    .A2(_04570_),
    .B1(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__a21o_1 _11381_ (.A1(\rbzero.texu_hot[3] ),
    .A2(_04553_),
    .B1(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__and2b_1 _11382_ (.A_N(_04550_),
    .B(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__a21oi_1 _11383_ (.A1(\rbzero.texu_hot[4] ),
    .A2(_04549_),
    .B1(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__nor2_1 _11384_ (.A(_04546_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__a21oi_2 _11385_ (.A1(\rbzero.texu_hot[5] ),
    .A2(_04545_),
    .B1(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__nor2_1 _11386_ (.A(_04542_),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__mux2_1 _11387_ (.A0(\rbzero.spi_registers.texadd0[13] ),
    .A1(\rbzero.spi_registers.texadd2[13] ),
    .S(\rbzero.wall_hot[1] ),
    .X(_04579_));
 sky130_fd_sc_hd__o21ba_1 _11388_ (.A1(_04519_),
    .A2(_04579_),
    .B1_N(_04534_),
    .X(_04580_));
 sky130_fd_sc_hd__o21a_1 _11389_ (.A1(_04540_),
    .A2(_04578_),
    .B1(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__or2_1 _11390_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_04517_),
    .X(_04582_));
 sky130_fd_sc_hd__inv_2 _11391_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .Y(_04583_));
 sky130_fd_sc_hd__a21oi_1 _11392_ (.A1(_04583_),
    .A2(_04524_),
    .B1(_04532_),
    .Y(_04584_));
 sky130_fd_sc_hd__o211a_1 _11393_ (.A1(_04534_),
    .A2(_04581_),
    .B1(_04582_),
    .C1(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__o21a_1 _11394_ (.A1(\rbzero.spi_registers.texadd3[15] ),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04586_));
 sky130_fd_sc_hd__a221o_1 _11395_ (.A1(\rbzero.spi_registers.texadd2[15] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[15] ),
    .C1(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__o21a_1 _11396_ (.A1(\rbzero.spi_registers.texadd0[15] ),
    .A2(_04517_),
    .B1(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__o21a_1 _11397_ (.A1(_04532_),
    .A2(_04585_),
    .B1(_04588_),
    .X(_04589_));
 sky130_fd_sc_hd__o21a_1 _11398_ (.A1(\rbzero.spi_registers.texadd3[16] ),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04590_));
 sky130_fd_sc_hd__a221o_1 _11399_ (.A1(\rbzero.spi_registers.texadd2[16] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[16] ),
    .C1(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__o21a_1 _11400_ (.A1(\rbzero.spi_registers.texadd0[16] ),
    .A2(_04517_),
    .B1(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__and2_1 _11401_ (.A(_04589_),
    .B(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__o21a_1 _11402_ (.A1(\rbzero.spi_registers.texadd3[17] ),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04594_));
 sky130_fd_sc_hd__a221o_1 _11403_ (.A1(\rbzero.spi_registers.texadd2[17] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[17] ),
    .C1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__o21a_1 _11404_ (.A1(\rbzero.spi_registers.texadd0[17] ),
    .A2(_04517_),
    .B1(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__nand2_1 _11405_ (.A(_04593_),
    .B(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__o21a_1 _11406_ (.A1(\rbzero.spi_registers.texadd3[18] ),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04598_));
 sky130_fd_sc_hd__a221o_1 _11407_ (.A1(\rbzero.spi_registers.texadd2[18] ),
    .A2(_04521_),
    .B1(_04524_),
    .B2(\rbzero.spi_registers.texadd1[18] ),
    .C1(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__o21ai_1 _11408_ (.A1(\rbzero.spi_registers.texadd0[18] ),
    .A2(_04518_),
    .B1(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__nor2_1 _11409_ (.A(_04597_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__and2_1 _11410_ (.A(_04530_),
    .B(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__clkbuf_4 _11411_ (.A(_04526_),
    .X(_04603_));
 sky130_fd_sc_hd__buf_4 _11412_ (.A(_04527_),
    .X(_04604_));
 sky130_fd_sc_hd__o21a_1 _11413_ (.A1(\rbzero.spi_registers.texadd3[20] ),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__a221o_1 _11414_ (.A1(\rbzero.spi_registers.texadd2[20] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[20] ),
    .C1(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__o21a_1 _11415_ (.A1(\rbzero.spi_registers.texadd0[20] ),
    .A2(_04518_),
    .B1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__nand2_1 _11416_ (.A(_04602_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__o21a_1 _11417_ (.A1(\rbzero.spi_registers.texadd3[21] ),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04609_));
 sky130_fd_sc_hd__a221o_1 _11418_ (.A1(\rbzero.spi_registers.texadd2[21] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[21] ),
    .C1(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__o21ai_1 _11419_ (.A1(\rbzero.spi_registers.texadd0[21] ),
    .A2(_04518_),
    .B1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nor2_1 _11420_ (.A(_04608_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__o21a_1 _11421_ (.A1(\rbzero.spi_registers.texadd3[22] ),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04613_));
 sky130_fd_sc_hd__a221o_1 _11422_ (.A1(\rbzero.spi_registers.texadd2[22] ),
    .A2(_04603_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[22] ),
    .C1(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__o21a_1 _11423_ (.A1(\rbzero.spi_registers.texadd0[22] ),
    .A2(_04518_),
    .B1(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__or3_1 _11424_ (.A(_04111_),
    .B(_04612_),
    .C(_04615_),
    .X(_04616_));
 sky130_fd_sc_hd__and3_1 _11425_ (.A(\rbzero.spi_registers.texadd1[23] ),
    .B(\rbzero.wall_hot[1] ),
    .C(_04519_),
    .X(_04617_));
 sky130_fd_sc_hd__nor2_1 _11426_ (.A(\rbzero.wall_hot[1] ),
    .B(_04519_),
    .Y(_04618_));
 sky130_fd_sc_hd__a221o_1 _11427_ (.A1(\rbzero.spi_registers.texadd3[23] ),
    .A2(_04604_),
    .B1(_04522_),
    .B2(\rbzero.spi_registers.texadd2[23] ),
    .C1(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__o22a_1 _11428_ (.A1(\rbzero.spi_registers.texadd0[23] ),
    .A2(_04518_),
    .B1(_04617_),
    .B2(_04619_),
    .X(_04620_));
 sky130_fd_sc_hd__nor2_1 _11429_ (.A(_04029_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__a21oi_1 _11430_ (.A1(_04612_),
    .A2(_04615_),
    .B1(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__and3_1 _11431_ (.A(_04612_),
    .B(_04615_),
    .C(_04621_),
    .X(_04623_));
 sky130_fd_sc_hd__a211oi_1 _11432_ (.A1(_04616_),
    .A2(_04622_),
    .B1(_04508_),
    .C1(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__nor2_1 _11433_ (.A(_04602_),
    .B(_04607_),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_1 _11434_ (.A(_04029_),
    .B(_04608_),
    .Y(_04626_));
 sky130_fd_sc_hd__and2_1 _11435_ (.A(_04608_),
    .B(_04611_),
    .X(_04627_));
 sky130_fd_sc_hd__or2_1 _11436_ (.A(_04612_),
    .B(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__o221a_1 _11437_ (.A1(_04625_),
    .A2(_04626_),
    .B1(_04628_),
    .B2(_04030_),
    .C1(_04508_),
    .X(_04629_));
 sky130_fd_sc_hd__nor2_1 _11438_ (.A(_04530_),
    .B(_04601_),
    .Y(_04630_));
 sky130_fd_sc_hd__or3_1 _11439_ (.A(_04029_),
    .B(_04602_),
    .C(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__and2_1 _11440_ (.A(_04597_),
    .B(_04600_),
    .X(_04632_));
 sky130_fd_sc_hd__clkinv_4 _11441_ (.A(\gpout0.hpos[1] ),
    .Y(_04633_));
 sky130_fd_sc_hd__o31a_1 _11442_ (.A1(_04111_),
    .A2(_04601_),
    .A3(_04632_),
    .B1(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__or2_1 _11443_ (.A(_04593_),
    .B(_04596_),
    .X(_04635_));
 sky130_fd_sc_hd__nor2_1 _11444_ (.A(_04111_),
    .B(_04593_),
    .Y(_04636_));
 sky130_fd_sc_hd__or2_1 _11445_ (.A(_04589_),
    .B(_04592_),
    .X(_04637_));
 sky130_fd_sc_hd__a32oi_1 _11446_ (.A1(_04111_),
    .A2(_04597_),
    .A3(_04635_),
    .B1(_04636_),
    .B2(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__inv_2 _11447_ (.A(\gpout0.hpos[2] ),
    .Y(_04639_));
 sky130_fd_sc_hd__a221o_1 _11448_ (.A1(_04631_),
    .A2(_04634_),
    .B1(_04638_),
    .B2(_04508_),
    .C1(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__o31a_1 _11449_ (.A1(_04506_),
    .A2(_04624_),
    .A3(_04629_),
    .B1(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__buf_4 _11450_ (.A(\gpout0.hpos[4] ),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_4 _11451_ (.A(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__nor2_1 _11452_ (.A(_04513_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__o32a_1 _11453_ (.A1(_04513_),
    .A2(_04514_),
    .A3(_04641_),
    .B1(_04644_),
    .B2(_04478_),
    .X(_04645_));
 sky130_fd_sc_hd__nor2_1 _11454_ (.A(net72),
    .B(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__xnor2_1 _11455_ (.A(_04550_),
    .B(_04573_),
    .Y(_04647_));
 sky130_fd_sc_hd__or2_1 _11456_ (.A(_04029_),
    .B(_04576_),
    .X(_04648_));
 sky130_fd_sc_hd__a21oi_1 _11457_ (.A1(_04546_),
    .A2(_04575_),
    .B1(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__a211o_1 _11458_ (.A1(_04030_),
    .A2(_04647_),
    .B1(_04649_),
    .C1(_04508_),
    .X(_04650_));
 sky130_fd_sc_hd__and3_1 _11459_ (.A(_04557_),
    .B(_04570_),
    .C(_04571_),
    .X(_04651_));
 sky130_fd_sc_hd__or2_1 _11460_ (.A(_04029_),
    .B(_04572_),
    .X(_04652_));
 sky130_fd_sc_hd__xnor2_1 _11461_ (.A(_04559_),
    .B(_04569_),
    .Y(_04653_));
 sky130_fd_sc_hd__o221ai_1 _11462_ (.A1(_04651_),
    .A2(_04652_),
    .B1(_04653_),
    .B2(_04111_),
    .C1(_04508_),
    .Y(_04654_));
 sky130_fd_sc_hd__nor2_1 _11463_ (.A(_04508_),
    .B(_04589_),
    .Y(_04655_));
 sky130_fd_sc_hd__o31a_1 _11464_ (.A1(_04532_),
    .A2(_04585_),
    .A3(_04588_),
    .B1(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__nor2_1 _11465_ (.A(_04633_),
    .B(_04581_),
    .Y(_04657_));
 sky130_fd_sc_hd__o31a_1 _11466_ (.A1(_04540_),
    .A2(_04578_),
    .A3(_04580_),
    .B1(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__xnor2_1 _11467_ (.A(_04542_),
    .B(_04577_),
    .Y(_04659_));
 sky130_fd_sc_hd__a211o_1 _11468_ (.A1(_04582_),
    .A2(_04584_),
    .B1(_04534_),
    .C1(_04581_),
    .X(_04660_));
 sky130_fd_sc_hd__or3b_1 _11469_ (.A(_04507_),
    .B(_04585_),
    .C_N(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__o211ai_1 _11470_ (.A1(_04633_),
    .A2(_04659_),
    .B1(_04661_),
    .C1(_04030_),
    .Y(_04662_));
 sky130_fd_sc_hd__o311a_1 _11471_ (.A1(_04030_),
    .A2(_04656_),
    .A3(_04658_),
    .B1(_04662_),
    .C1(_04639_),
    .X(_04663_));
 sky130_fd_sc_hd__a311o_1 _11472_ (.A1(_04506_),
    .A2(_04650_),
    .A3(_04654_),
    .B1(_04643_),
    .C1(_04663_),
    .X(_04664_));
 sky130_fd_sc_hd__a22o_1 _11473_ (.A1(\rbzero.spi_registers.texadd2[0] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[0] ),
    .X(_04665_));
 sky130_fd_sc_hd__o21a_1 _11474_ (.A1(\rbzero.spi_registers.texadd3[0] ),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04666_));
 sky130_fd_sc_hd__o22a_1 _11475_ (.A1(\rbzero.spi_registers.texadd0[0] ),
    .A2(_04518_),
    .B1(_04665_),
    .B2(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__a22o_1 _11476_ (.A1(\rbzero.spi_registers.texadd2[1] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[1] ),
    .X(_04668_));
 sky130_fd_sc_hd__o21a_1 _11477_ (.A1(\rbzero.spi_registers.texadd3[1] ),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04669_));
 sky130_fd_sc_hd__o221a_1 _11478_ (.A1(\rbzero.spi_registers.texadd0[1] ),
    .A2(_04518_),
    .B1(_04668_),
    .B2(_04669_),
    .C1(_04111_),
    .X(_04670_));
 sky130_fd_sc_hd__a211o_1 _11479_ (.A1(_04030_),
    .A2(_04667_),
    .B1(_04670_),
    .C1(_04633_),
    .X(_04671_));
 sky130_fd_sc_hd__a22o_1 _11480_ (.A1(\rbzero.spi_registers.texadd2[2] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[2] ),
    .X(_04672_));
 sky130_fd_sc_hd__o21a_1 _11481_ (.A1(\rbzero.spi_registers.texadd3[2] ),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04673_));
 sky130_fd_sc_hd__o22a_1 _11482_ (.A1(\rbzero.spi_registers.texadd0[2] ),
    .A2(_04518_),
    .B1(_04672_),
    .B2(_04673_),
    .X(_04674_));
 sky130_fd_sc_hd__a22o_1 _11483_ (.A1(\rbzero.spi_registers.texadd2[3] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[3] ),
    .X(_04675_));
 sky130_fd_sc_hd__o21a_1 _11484_ (.A1(\rbzero.spi_registers.texadd3[3] ),
    .A2(_04603_),
    .B1(_04604_),
    .X(_04676_));
 sky130_fd_sc_hd__o221a_1 _11485_ (.A1(\rbzero.spi_registers.texadd0[3] ),
    .A2(_04518_),
    .B1(_04675_),
    .B2(_04676_),
    .C1(_04111_),
    .X(_04677_));
 sky130_fd_sc_hd__a211o_1 _11486_ (.A1(_04030_),
    .A2(_04674_),
    .B1(_04677_),
    .C1(_04508_),
    .X(_04678_));
 sky130_fd_sc_hd__and2_1 _11487_ (.A(_04566_),
    .B(_04567_),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _11488_ (.A(_04029_),
    .B(_04566_),
    .Y(_04680_));
 sky130_fd_sc_hd__a21oi_1 _11489_ (.A1(_04564_),
    .A2(_04565_),
    .B1(\rbzero.texu_hot[0] ),
    .Y(_04681_));
 sky130_fd_sc_hd__o32a_1 _11490_ (.A1(_04030_),
    .A2(_04568_),
    .A3(_04679_),
    .B1(_04680_),
    .B2(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__a22o_1 _11491_ (.A1(\rbzero.spi_registers.texadd2[4] ),
    .A2(_04522_),
    .B1(_04618_),
    .B2(\rbzero.spi_registers.texadd0[4] ),
    .X(_04683_));
 sky130_fd_sc_hd__a21oi_1 _11492_ (.A1(\rbzero.spi_registers.texadd1[4] ),
    .A2(_04525_),
    .B1(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__or3b_1 _11493_ (.A(\rbzero.wall_hot[1] ),
    .B(_04603_),
    .C_N(\rbzero.spi_registers.texadd3[4] ),
    .X(_04685_));
 sky130_fd_sc_hd__a31o_1 _11494_ (.A1(\rbzero.spi_registers.texadd3[5] ),
    .A2(_04604_),
    .A3(_04519_),
    .B1(_04029_),
    .X(_04686_));
 sky130_fd_sc_hd__a22o_1 _11495_ (.A1(\rbzero.spi_registers.texadd2[5] ),
    .A2(_04522_),
    .B1(_04525_),
    .B2(\rbzero.spi_registers.texadd1[5] ),
    .X(_04687_));
 sky130_fd_sc_hd__a211oi_1 _11496_ (.A1(\rbzero.spi_registers.texadd0[5] ),
    .A2(_04618_),
    .B1(_04686_),
    .C1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__a31o_1 _11497_ (.A1(_04029_),
    .A2(_04684_),
    .A3(_04685_),
    .B1(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__a21o_1 _11498_ (.A1(_04508_),
    .A2(_04689_),
    .B1(_04506_),
    .X(_04690_));
 sky130_fd_sc_hd__a21oi_1 _11499_ (.A1(_04633_),
    .A2(_04682_),
    .B1(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__a311o_1 _11500_ (.A1(_04506_),
    .A2(_04671_),
    .A3(_04678_),
    .B1(_04691_),
    .C1(_04513_),
    .X(_04692_));
 sky130_fd_sc_hd__or2_1 _11501_ (.A(_04481_),
    .B(_04472_),
    .X(_04693_));
 sky130_fd_sc_hd__a31o_1 _11502_ (.A1(_04664_),
    .A2(_04692_),
    .A3(_04693_),
    .B1(_04644_),
    .X(_04694_));
 sky130_fd_sc_hd__a32o_2 _11503_ (.A1(_04478_),
    .A2(_04505_),
    .A3(_04512_),
    .B1(_04646_),
    .B2(_04694_),
    .X(net73));
 sky130_fd_sc_hd__inv_2 _20688__4 (.A(clknet_1_0__leaf__03503_),
    .Y(net129));
 sky130_fd_sc_hd__clkinv_2 _11505_ (.A(net2),
    .Y(_04695_));
 sky130_fd_sc_hd__and3_2 _11506_ (.A(\gpout0.hpos[2] ),
    .B(\gpout0.hpos[1] ),
    .C(\gpout0.hpos[0] ),
    .X(_04696_));
 sky130_fd_sc_hd__or3_4 _11507_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(\gpout0.vpos[0] ),
    .X(_04697_));
 sky130_fd_sc_hd__inv_2 _11508_ (.A(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__clkbuf_4 _11509_ (.A(\gpout0.vpos[5] ),
    .X(_04699_));
 sky130_fd_sc_hd__nor2_2 _11510_ (.A(_04699_),
    .B(\gpout0.vpos[4] ),
    .Y(_04700_));
 sky130_fd_sc_hd__clkbuf_4 _11511_ (.A(\gpout0.vpos[4] ),
    .X(_04701_));
 sky130_fd_sc_hd__or2_2 _11512_ (.A(_04701_),
    .B(\gpout0.vpos[3] ),
    .X(_04702_));
 sky130_fd_sc_hd__nand2_1 _11513_ (.A(_04701_),
    .B(\gpout0.vpos[3] ),
    .Y(_04703_));
 sky130_fd_sc_hd__clkbuf_4 _11514_ (.A(_04699_),
    .X(_04704_));
 sky130_fd_sc_hd__nand2_2 _11515_ (.A(_04704_),
    .B(_04701_),
    .Y(_04705_));
 sky130_fd_sc_hd__and4b_1 _11516_ (.A_N(_04700_),
    .B(_04702_),
    .C(_04703_),
    .D(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__nor2_1 _11517_ (.A(_04633_),
    .B(_04110_),
    .Y(_04707_));
 sky130_fd_sc_hd__nand2_1 _11518_ (.A(\gpout0.hpos[2] ),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__nor2_1 _11519_ (.A(_04475_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__or2_1 _11520_ (.A(\gpout0.hpos[4] ),
    .B(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__o21ai_1 _11521_ (.A1(\gpout0.hpos[5] ),
    .A2(_04710_),
    .B1(_04479_),
    .Y(_04711_));
 sky130_fd_sc_hd__nor2_1 _11522_ (.A(_04501_),
    .B(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__a21oi_2 _11523_ (.A1(\gpout0.hpos[8] ),
    .A2(_04712_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04713_));
 sky130_fd_sc_hd__clkbuf_4 _11524_ (.A(\gpout0.vpos[7] ),
    .X(_04714_));
 sky130_fd_sc_hd__or4b_1 _11525_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.vpos[8] ),
    .C(_04714_),
    .D_N(net3),
    .X(_04715_));
 sky130_fd_sc_hd__inv_2 _11526_ (.A(\gpout0.vpos[3] ),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_2 _11527_ (.A(_04716_),
    .B(_04700_),
    .Y(_04717_));
 sky130_fd_sc_hd__clkbuf_4 _11528_ (.A(\gpout0.vpos[6] ),
    .X(_04718_));
 sky130_fd_sc_hd__o21a_1 _11529_ (.A1(_04717_),
    .A2(_04697_),
    .B1(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__nor3_4 _11530_ (.A(_04713_),
    .B(_04715_),
    .C(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__o31a_1 _11531_ (.A1(_04696_),
    .A2(_04698_),
    .A3(_04706_),
    .B1(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__xor2_1 _11532_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .B(_04474_),
    .X(_04722_));
 sky130_fd_sc_hd__buf_6 _11533_ (.A(\gpout0.vpos[3] ),
    .X(_04723_));
 sky130_fd_sc_hd__xor2_1 _11534_ (.A(_04723_),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .X(_04724_));
 sky130_fd_sc_hd__clkinv_2 _11535_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .Y(_04725_));
 sky130_fd_sc_hd__xnor2_1 _11536_ (.A(_04718_),
    .B(\rbzero.debug_overlay.playerY[3] ),
    .Y(_04726_));
 sky130_fd_sc_hd__o221a_1 _11537_ (.A1(_04714_),
    .A2(_04725_),
    .B1(\rbzero.debug_overlay.playerX[0] ),
    .B2(_04476_),
    .C1(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__or3b_1 _11538_ (.A(_04722_),
    .B(_04724_),
    .C_N(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__clkinv_2 _11539_ (.A(_04699_),
    .Y(_04729_));
 sky130_fd_sc_hd__inv_2 _11540_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .Y(_04730_));
 sky130_fd_sc_hd__a22o_1 _11541_ (.A1(_04729_),
    .A2(\rbzero.debug_overlay.playerY[2] ),
    .B1(_04730_),
    .B2(_04480_),
    .X(_04731_));
 sky130_fd_sc_hd__a221o_1 _11542_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_04476_),
    .B1(_04477_),
    .B2(\rbzero.debug_overlay.playerX[1] ),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__inv_2 _11543_ (.A(\gpout0.vpos[4] ),
    .Y(_04733_));
 sky130_fd_sc_hd__buf_2 _11544_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .X(_04734_));
 sky130_fd_sc_hd__inv_2 _11545_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .Y(_04735_));
 sky130_fd_sc_hd__inv_2 _11546_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .Y(_04736_));
 sky130_fd_sc_hd__a2bb2o_1 _11547_ (.A1_N(\rbzero.debug_overlay.playerY[1] ),
    .A2_N(_04733_),
    .B1(_04699_),
    .B2(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__a221o_1 _11548_ (.A1(_04733_),
    .A2(_04734_),
    .B1(_04735_),
    .B2(_04642_),
    .C1(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__inv_2 _11549_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .Y(_04739_));
 sky130_fd_sc_hd__a22o_1 _11550_ (.A1(_04714_),
    .A2(_04725_),
    .B1(_04739_),
    .B2(_04031_),
    .X(_04740_));
 sky130_fd_sc_hd__a221o_1 _11551_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_04501_),
    .B1(_04514_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .C1(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__or3_1 _11552_ (.A(_04732_),
    .B(_04738_),
    .C(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__nor2_2 _11553_ (.A(_04728_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__buf_2 _11554_ (.A(\gpout0.vpos[1] ),
    .X(_04744_));
 sky130_fd_sc_hd__inv_2 _11555_ (.A(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__inv_2 _11556_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .Y(_04746_));
 sky130_fd_sc_hd__nor2_1 _11557_ (.A(_04745_),
    .B(_04746_),
    .Y(_04747_));
 sky130_fd_sc_hd__nor2_1 _11558_ (.A(_04744_),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .Y(_04748_));
 sky130_fd_sc_hd__inv_2 _11559_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .Y(_04749_));
 sky130_fd_sc_hd__nor2_1 _11560_ (.A(_04749_),
    .B(_04111_),
    .Y(_04750_));
 sky130_fd_sc_hd__nor2_1 _11561_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(\gpout0.hpos[0] ),
    .Y(_04751_));
 sky130_fd_sc_hd__clkinv_2 _11562_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .Y(_04752_));
 sky130_fd_sc_hd__xnor2_1 _11563_ (.A(\gpout0.vpos[2] ),
    .B(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_04753_));
 sky130_fd_sc_hd__o221a_1 _11564_ (.A1(\gpout0.vpos[0] ),
    .A2(_04752_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .B2(_04639_),
    .C1(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__o221a_1 _11565_ (.A1(_04747_),
    .A2(_04748_),
    .B1(_04750_),
    .B2(_04751_),
    .C1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__xor2_1 _11566_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_04507_),
    .X(_04756_));
 sky130_fd_sc_hd__a221oi_1 _11567_ (.A1(\gpout0.vpos[0] ),
    .A2(_04752_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .B2(_04639_),
    .C1(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__or2_1 _11568_ (.A(_04714_),
    .B(_04718_),
    .X(_04758_));
 sky130_fd_sc_hd__o31a_1 _11569_ (.A1(_04717_),
    .A2(_04697_),
    .A3(_04758_),
    .B1(\gpout0.vpos[8] ),
    .X(_04759_));
 sky130_fd_sc_hd__or3b_1 _11570_ (.A(\gpout0.vpos[9] ),
    .B(_04034_),
    .C_N(net1),
    .X(_04760_));
 sky130_fd_sc_hd__or2_2 _11571_ (.A(_04031_),
    .B(_04480_),
    .X(_04761_));
 sky130_fd_sc_hd__or3_1 _11572_ (.A(_04471_),
    .B(_04642_),
    .C(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__o31a_1 _11573_ (.A1(_04474_),
    .A2(_04510_),
    .A3(_04762_),
    .B1(_04033_),
    .X(_04763_));
 sky130_fd_sc_hd__or3_4 _11574_ (.A(_04759_),
    .B(_04760_),
    .C(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__a31o_1 _11575_ (.A1(_04743_),
    .A2(_04755_),
    .A3(_04757_),
    .B1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__nand2_1 _11576_ (.A(_04510_),
    .B(_04697_),
    .Y(_04766_));
 sky130_fd_sc_hd__or2_1 _11577_ (.A(_04743_),
    .B(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__inv_2 _11578_ (.A(\gpout0.vpos[7] ),
    .Y(_04768_));
 sky130_fd_sc_hd__a22o_1 _11579_ (.A1(_04768_),
    .A2(\rbzero.map_overlay.i_mapdy[4] ),
    .B1(\rbzero.map_overlay.i_mapdy[2] ),
    .B2(_04729_),
    .X(_04769_));
 sky130_fd_sc_hd__inv_2 _11580_ (.A(\gpout0.vpos[6] ),
    .Y(_04770_));
 sky130_fd_sc_hd__inv_2 _11581_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .Y(_04771_));
 sky130_fd_sc_hd__xor2_1 _11582_ (.A(_04701_),
    .B(\rbzero.map_overlay.i_mapdy[1] ),
    .X(_04772_));
 sky130_fd_sc_hd__a221o_1 _11583_ (.A1(_04770_),
    .A2(\rbzero.map_overlay.i_mapdy[3] ),
    .B1(_04771_),
    .B2(_04699_),
    .C1(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__or4_1 _11584_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_overlay.i_mapdy[2] ),
    .C(\rbzero.map_overlay.i_mapdy[1] ),
    .D(\rbzero.map_overlay.i_mapdy[0] ),
    .X(_04774_));
 sky130_fd_sc_hd__o21a_1 _11585_ (.A1(\rbzero.map_overlay.i_mapdy[5] ),
    .A2(_04774_),
    .B1(_04768_),
    .X(_04775_));
 sky130_fd_sc_hd__inv_2 _11586_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .Y(_04776_));
 sky130_fd_sc_hd__o22a_1 _11587_ (.A1(_04770_),
    .A2(\rbzero.map_overlay.i_mapdy[3] ),
    .B1(_04776_),
    .B2(\gpout0.vpos[3] ),
    .X(_04777_));
 sky130_fd_sc_hd__o221a_1 _11588_ (.A1(_04716_),
    .A2(\rbzero.map_overlay.i_mapdy[0] ),
    .B1(_04775_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__or3b_1 _11589_ (.A(_04769_),
    .B(_04773_),
    .C_N(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__a22o_1 _11590_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04476_),
    .B1(_04477_),
    .B2(\rbzero.map_overlay.i_mapdx[1] ),
    .X(_04780_));
 sky130_fd_sc_hd__o22a_1 _11591_ (.A1(\rbzero.map_overlay.i_mapdx[4] ),
    .A2(_04501_),
    .B1(_04477_),
    .B2(\rbzero.map_overlay.i_mapdx[1] ),
    .X(_04781_));
 sky130_fd_sc_hd__or4_1 _11592_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(\rbzero.map_overlay.i_mapdx[2] ),
    .C(\rbzero.map_overlay.i_mapdx[1] ),
    .D(\rbzero.map_overlay.i_mapdx[0] ),
    .X(_04782_));
 sky130_fd_sc_hd__inv_2 _11593_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .Y(_04783_));
 sky130_fd_sc_hd__o21a_1 _11594_ (.A1(\rbzero.map_overlay.i_mapdx[5] ),
    .A2(_04782_),
    .B1(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__xnor2_1 _11595_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_04480_),
    .Y(_04785_));
 sky130_fd_sc_hd__o221a_1 _11596_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04476_),
    .B1(_04031_),
    .B2(_04784_),
    .C1(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__xnor2_1 _11597_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_04474_),
    .Y(_04787_));
 sky130_fd_sc_hd__and4b_1 _11598_ (.A_N(_04780_),
    .B(_04781_),
    .C(_04786_),
    .D(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__xor2_1 _11599_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_04031_),
    .X(_04789_));
 sky130_fd_sc_hd__a221o_1 _11600_ (.A1(\rbzero.map_overlay.i_otherx[0] ),
    .A2(_04476_),
    .B1(_04514_),
    .B2(\rbzero.map_overlay.i_otherx[3] ),
    .C1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__inv_2 _11601_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .Y(_04791_));
 sky130_fd_sc_hd__inv_2 _11602_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .Y(_04792_));
 sky130_fd_sc_hd__inv_2 _11603_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .Y(_04793_));
 sky130_fd_sc_hd__a22o_1 _11604_ (.A1(_04793_),
    .A2(_04480_),
    .B1(_04477_),
    .B2(\rbzero.map_overlay.i_otherx[1] ),
    .X(_04794_));
 sky130_fd_sc_hd__a221o_1 _11605_ (.A1(_04714_),
    .A2(_04791_),
    .B1(_04792_),
    .B2(_04642_),
    .C1(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__xnor2_1 _11606_ (.A(\gpout0.vpos[3] ),
    .B(\rbzero.map_overlay.i_othery[0] ),
    .Y(_04796_));
 sky130_fd_sc_hd__inv_2 _11607_ (.A(\rbzero.map_overlay.i_othery[3] ),
    .Y(_04797_));
 sky130_fd_sc_hd__xnor2_1 _11608_ (.A(\gpout0.vpos[4] ),
    .B(\rbzero.map_overlay.i_othery[1] ),
    .Y(_04798_));
 sky130_fd_sc_hd__o221a_1 _11609_ (.A1(_04718_),
    .A2(_04797_),
    .B1(\rbzero.map_overlay.i_otherx[0] ),
    .B2(_04476_),
    .C1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__xnor2_1 _11610_ (.A(\gpout0.vpos[5] ),
    .B(\rbzero.map_overlay.i_othery[2] ),
    .Y(_04800_));
 sky130_fd_sc_hd__clkinv_2 _11611_ (.A(_04473_),
    .Y(_04801_));
 sky130_fd_sc_hd__o2bb2a_1 _11612_ (.A1_N(\rbzero.map_overlay.i_otherx[2] ),
    .A2_N(_04801_),
    .B1(\gpout0.vpos[7] ),
    .B2(_04791_),
    .X(_04802_));
 sky130_fd_sc_hd__o221a_1 _11613_ (.A1(_04770_),
    .A2(\rbzero.map_overlay.i_othery[3] ),
    .B1(\rbzero.map_overlay.i_otherx[2] ),
    .B2(_04801_),
    .C1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__and4_1 _11614_ (.A(_04796_),
    .B(_04799_),
    .C(_04800_),
    .D(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__or3b_1 _11615_ (.A(_04790_),
    .B(_04795_),
    .C_N(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__o21a_1 _11616_ (.A1(_04779_),
    .A2(_04788_),
    .B1(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__nor2_1 _11617_ (.A(_04767_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__a21oi_4 _11618_ (.A1(\gpout0.hpos[8] ),
    .A2(_04761_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04808_));
 sky130_fd_sc_hd__mux2_1 _11619_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__nand2_1 _11620_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .Y(_04810_));
 sky130_fd_sc_hd__or2_1 _11621_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .X(_04811_));
 sky130_fd_sc_hd__nand3_1 _11622_ (.A(\rbzero.texV[4] ),
    .B(_04810_),
    .C(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__a21o_1 _11623_ (.A1(_04810_),
    .A2(_04811_),
    .B1(\rbzero.texV[4] ),
    .X(_04813_));
 sky130_fd_sc_hd__nand2_1 _11624_ (.A(_04812_),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__or2_1 _11625_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .X(_04815_));
 sky130_fd_sc_hd__nand2_1 _11626_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .Y(_04816_));
 sky130_fd_sc_hd__a21boi_1 _11627_ (.A1(\rbzero.texV[3] ),
    .A2(_04815_),
    .B1_N(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__xnor2_1 _11628_ (.A(_04814_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__nand2_1 _11629_ (.A(_04816_),
    .B(_04815_),
    .Y(_04819_));
 sky130_fd_sc_hd__xor2_1 _11630_ (.A(\rbzero.texV[3] ),
    .B(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__o211a_1 _11631_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(\rbzero.texV[1] ),
    .B1(\rbzero.texV[0] ),
    .C1(\rbzero.traced_texVinit[0] ),
    .X(_04821_));
 sky130_fd_sc_hd__a221o_1 _11632_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(\rbzero.texV[1] ),
    .B2(\rbzero.traced_texVinit[1] ),
    .C1(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__o21ai_1 _11633_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__or2_1 _11634_ (.A(_04820_),
    .B(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__nor2_1 _11635_ (.A(_04818_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__nand2_1 _11636_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_04826_));
 sky130_fd_sc_hd__or2_1 _11637_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .X(_04827_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(_04826_),
    .B(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__or2_1 _11639_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .X(_04829_));
 sky130_fd_sc_hd__nand2_1 _11640_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .Y(_04830_));
 sky130_fd_sc_hd__a21boi_1 _11641_ (.A1(\rbzero.texV[8] ),
    .A2(_04829_),
    .B1_N(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__nand2_1 _11642_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .Y(_04832_));
 sky130_fd_sc_hd__or2_1 _11643_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .X(_04833_));
 sky130_fd_sc_hd__nand3_1 _11644_ (.A(\rbzero.texV[7] ),
    .B(_04832_),
    .C(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__a21o_1 _11645_ (.A1(_04832_),
    .A2(_04833_),
    .B1(\rbzero.texV[7] ),
    .X(_04835_));
 sky130_fd_sc_hd__nand2_1 _11646_ (.A(_04834_),
    .B(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__nand2_1 _11647_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .Y(_04837_));
 sky130_fd_sc_hd__or2_1 _11648_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .X(_04838_));
 sky130_fd_sc_hd__nand3_1 _11649_ (.A(\rbzero.texV[6] ),
    .B(_04837_),
    .C(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand3_1 _11650_ (.A(_04836_),
    .B(_04837_),
    .C(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__a21o_1 _11651_ (.A1(_04837_),
    .A2(_04838_),
    .B1(\rbzero.texV[6] ),
    .X(_04841_));
 sky130_fd_sc_hd__nand2_1 _11652_ (.A(_04839_),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__and2_1 _11653_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .X(_04843_));
 sky130_fd_sc_hd__nor2_1 _11654_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .Y(_04844_));
 sky130_fd_sc_hd__nor2_1 _11655_ (.A(_04843_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__a21oi_2 _11656_ (.A1(\rbzero.texV[5] ),
    .A2(_04845_),
    .B1(_04843_),
    .Y(_04846_));
 sky130_fd_sc_hd__xnor2_1 _11657_ (.A(_04842_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__xnor2_1 _11658_ (.A(\rbzero.texV[5] ),
    .B(_04845_),
    .Y(_04848_));
 sky130_fd_sc_hd__a21oi_1 _11659_ (.A1(_04810_),
    .A2(_04812_),
    .B1(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__nor2_1 _11660_ (.A(_04814_),
    .B(_04817_),
    .Y(_04850_));
 sky130_fd_sc_hd__and3_1 _11661_ (.A(_04848_),
    .B(_04810_),
    .C(_04812_),
    .X(_04851_));
 sky130_fd_sc_hd__or2_1 _11662_ (.A(_04849_),
    .B(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__inv_2 _11663_ (.A(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__o21a_1 _11664_ (.A1(_04850_),
    .A2(_04825_),
    .B1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__nor2_1 _11665_ (.A(_04849_),
    .B(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__nor2_1 _11666_ (.A(_04847_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__o21bai_4 _11667_ (.A1(_04842_),
    .A2(_04846_),
    .B1_N(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__a21oi_1 _11668_ (.A1(_04837_),
    .A2(_04839_),
    .B1(_04836_),
    .Y(_04858_));
 sky130_fd_sc_hd__a21o_1 _11669_ (.A1(_04840_),
    .A2(_04857_),
    .B1(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__nand2_1 _11670_ (.A(_04830_),
    .B(_04829_),
    .Y(_04860_));
 sky130_fd_sc_hd__xor2_1 _11671_ (.A(\rbzero.texV[8] ),
    .B(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__nand3_1 _11672_ (.A(_04832_),
    .B(_04834_),
    .C(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__nand2_1 _11673_ (.A(_04859_),
    .B(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__a21o_1 _11674_ (.A1(_04832_),
    .A2(_04834_),
    .B1(_04861_),
    .X(_04864_));
 sky130_fd_sc_hd__o21a_1 _11675_ (.A1(_04828_),
    .A2(_04831_),
    .B1(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__a22oi_2 _11676_ (.A1(_04828_),
    .A2(_04831_),
    .B1(_04863_),
    .B2(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__xor2_1 _11677_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .X(_04867_));
 sky130_fd_sc_hd__xnor2_1 _11678_ (.A(_04826_),
    .B(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__a21oi_1 _11679_ (.A1(_04866_),
    .A2(_04868_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04869_));
 sky130_fd_sc_hd__o21a_4 _11680_ (.A1(_04866_),
    .A2(_04868_),
    .B1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__nand2_1 _11681_ (.A(_04818_),
    .B(_04824_),
    .Y(_04871_));
 sky130_fd_sc_hd__nor3b_1 _11682_ (.A(_04825_),
    .B(_04870_),
    .C_N(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__clkbuf_8 _11683_ (.A(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__nor3_1 _11684_ (.A(_04853_),
    .B(_04850_),
    .C(_04825_),
    .Y(_04874_));
 sky130_fd_sc_hd__nor3_4 _11685_ (.A(_04854_),
    .B(_04870_),
    .C(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__nor2_2 _11686_ (.A(_04873_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21oi_1 _11687_ (.A1(_04820_),
    .A2(_04823_),
    .B1(_04870_),
    .Y(_04877_));
 sky130_fd_sc_hd__and2_2 _11688_ (.A(_04824_),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__clkbuf_4 _11689_ (.A(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__nor2_1 _11690_ (.A(\rbzero.row_render.texu[0] ),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__inv_2 _11691_ (.A(\rbzero.row_render.texu[4] ),
    .Y(_04881_));
 sky130_fd_sc_hd__inv_2 _11692_ (.A(\rbzero.row_render.texu[3] ),
    .Y(_04882_));
 sky130_fd_sc_hd__and2_1 _11693_ (.A(_04847_),
    .B(_04855_),
    .X(_04883_));
 sky130_fd_sc_hd__nor3_4 _11694_ (.A(_04856_),
    .B(_04870_),
    .C(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__a41o_1 _11695_ (.A1(_04881_),
    .A2(_04882_),
    .A3(\rbzero.row_render.texu[2] ),
    .A4(\rbzero.row_render.texu[1] ),
    .B1(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__nor2_1 _11696_ (.A(\rbzero.row_render.texu[2] ),
    .B(\rbzero.row_render.texu[1] ),
    .Y(_04886_));
 sky130_fd_sc_hd__or3_2 _11697_ (.A(_04856_),
    .B(_04870_),
    .C(_04883_),
    .X(_04887_));
 sky130_fd_sc_hd__a31o_1 _11698_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(\rbzero.row_render.texu[3] ),
    .A3(_04886_),
    .B1(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__and3b_1 _11699_ (.A_N(\rbzero.row_render.texu[0] ),
    .B(_04885_),
    .C(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__a21o_1 _11700_ (.A1(_04876_),
    .A2(_04880_),
    .B1(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__or2_1 _11701_ (.A(\rbzero.row_render.side ),
    .B(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__buf_6 _11702_ (.A(_04824_),
    .X(_04892_));
 sky130_fd_sc_hd__buf_6 _11703_ (.A(_04877_),
    .X(_04893_));
 sky130_fd_sc_hd__nand2_4 _11704_ (.A(_04892_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__buf_4 _11705_ (.A(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__clkbuf_8 _11706_ (.A(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__buf_4 _11707_ (.A(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__clkbuf_4 _11708_ (.A(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__clkbuf_4 _11709_ (.A(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__inv_2 _11710_ (.A(\rbzero.row_render.side ),
    .Y(_04900_));
 sky130_fd_sc_hd__a31o_1 _11711_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04876_),
    .A3(_04899_),
    .B1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__and2b_1 _11712_ (.A_N(\rbzero.row_render.wall[0] ),
    .B(\rbzero.row_render.wall[1] ),
    .X(_04902_));
 sky130_fd_sc_hd__inv_2 _11713_ (.A(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__a21o_1 _11714_ (.A1(_04891_),
    .A2(_04901_),
    .B1(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__nor2b_2 _11715_ (.A(\rbzero.row_render.wall[1] ),
    .B_N(\rbzero.row_render.wall[0] ),
    .Y(_04905_));
 sky130_fd_sc_hd__inv_2 _11716_ (.A(net42),
    .Y(_04906_));
 sky130_fd_sc_hd__a21oi_1 _11717_ (.A1(_04900_),
    .A2(_04905_),
    .B1(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__buf_6 _11718_ (.A(_04887_),
    .X(_04908_));
 sky130_fd_sc_hd__a32o_1 _11719_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(\rbzero.row_render.texu[2] ),
    .A3(\rbzero.row_render.texu[1] ),
    .B1(_04908_),
    .B2(_04876_),
    .X(_04909_));
 sky130_fd_sc_hd__buf_4 _11720_ (.A(_04872_),
    .X(_04910_));
 sky130_fd_sc_hd__buf_4 _11721_ (.A(_04875_),
    .X(_04911_));
 sky130_fd_sc_hd__a32o_1 _11722_ (.A1(_04884_),
    .A2(_04910_),
    .A3(_04911_),
    .B1(_04886_),
    .B2(_04882_),
    .X(_04912_));
 sky130_fd_sc_hd__nor2_1 _11723_ (.A(\rbzero.row_render.side ),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__a31o_1 _11724_ (.A1(\rbzero.row_render.wall[0] ),
    .A2(_04909_),
    .A3(_04913_),
    .B1(_04905_),
    .X(_04914_));
 sky130_fd_sc_hd__inv_2 _11725_ (.A(_04912_),
    .Y(_04915_));
 sky130_fd_sc_hd__a41o_1 _11726_ (.A1(\rbzero.row_render.wall[0] ),
    .A2(\rbzero.row_render.wall[1] ),
    .A3(_04909_),
    .A4(_04915_),
    .B1(_04900_),
    .X(_04916_));
 sky130_fd_sc_hd__or3b_1 _11727_ (.A(_04902_),
    .B(_04914_),
    .C_N(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__buf_6 _11728_ (.A(_04884_),
    .X(_04918_));
 sky130_fd_sc_hd__buf_4 _11729_ (.A(_04894_),
    .X(_04919_));
 sky130_fd_sc_hd__buf_4 _11730_ (.A(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__and2_1 _11731_ (.A(\rbzero.tex_r0[52] ),
    .B(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__buf_4 _11732_ (.A(_04873_),
    .X(_04922_));
 sky130_fd_sc_hd__a31o_1 _11733_ (.A1(\rbzero.tex_r0[53] ),
    .A2(_04892_),
    .A3(_04893_),
    .B1(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__buf_4 _11734_ (.A(_04894_),
    .X(_04924_));
 sky130_fd_sc_hd__buf_4 _11735_ (.A(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__or3b_2 _11737_ (.A(_04825_),
    .B(_04870_),
    .C_N(_04871_),
    .X(_04927_));
 sky130_fd_sc_hd__buf_6 _11738_ (.A(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__buf_4 _11739_ (.A(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__buf_6 _11740_ (.A(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__buf_4 _11741_ (.A(_04875_),
    .X(_04931_));
 sky130_fd_sc_hd__buf_6 _11742_ (.A(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__o221a_1 _11743_ (.A1(_04921_),
    .A2(_04923_),
    .B1(_04926_),
    .B2(_04930_),
    .C1(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__buf_4 _11744_ (.A(_04922_),
    .X(_04934_));
 sky130_fd_sc_hd__mux2_1 _11745_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04925_),
    .X(_04935_));
 sky130_fd_sc_hd__clkbuf_4 _11746_ (.A(_04892_),
    .X(_04936_));
 sky130_fd_sc_hd__clkbuf_4 _11747_ (.A(_04893_),
    .X(_04937_));
 sky130_fd_sc_hd__and3_1 _11748_ (.A(\rbzero.tex_r0[51] ),
    .B(_04936_),
    .C(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__buf_6 _11749_ (.A(_04895_),
    .X(_04939_));
 sky130_fd_sc_hd__buf_4 _11750_ (.A(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__buf_6 _11751_ (.A(_04927_),
    .X(_04941_));
 sky130_fd_sc_hd__clkbuf_8 _11752_ (.A(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__a21o_1 _11753_ (.A1(\rbzero.tex_r0[50] ),
    .A2(_04940_),
    .B1(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__or3_2 _11754_ (.A(_04854_),
    .B(_04870_),
    .C(_04874_),
    .X(_04944_));
 sky130_fd_sc_hd__buf_6 _11755_ (.A(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__buf_6 _11756_ (.A(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__o221a_1 _11757_ (.A1(_04934_),
    .A2(_04935_),
    .B1(_04938_),
    .B2(_04943_),
    .C1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__inv_2 _11758_ (.A(_04840_),
    .Y(_04948_));
 sky130_fd_sc_hd__nor2_2 _11759_ (.A(_04948_),
    .B(_04858_),
    .Y(_04949_));
 sky130_fd_sc_hd__xnor2_4 _11760_ (.A(_04857_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nor2_8 _11761_ (.A(_04870_),
    .B(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__buf_6 _11762_ (.A(_04945_),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_1 _11763_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04919_),
    .X(_04953_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04919_),
    .X(_04954_));
 sky130_fd_sc_hd__mux2_1 _11765_ (.A0(_04953_),
    .A1(_04954_),
    .S(_04922_),
    .X(_04955_));
 sky130_fd_sc_hd__buf_4 _11766_ (.A(_04873_),
    .X(_04956_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04919_),
    .X(_04957_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04894_),
    .X(_04958_));
 sky130_fd_sc_hd__or2_1 _11769_ (.A(_04941_),
    .B(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__buf_6 _11770_ (.A(_04911_),
    .X(_04960_));
 sky130_fd_sc_hd__o211a_1 _11771_ (.A1(_04956_),
    .A2(_04957_),
    .B1(_04959_),
    .C1(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__a211o_1 _11772_ (.A1(_04952_),
    .A2(_04955_),
    .B1(_04961_),
    .C1(_04908_),
    .X(_04962_));
 sky130_fd_sc_hd__o311a_1 _11773_ (.A1(_04918_),
    .A2(_04933_),
    .A3(_04947_),
    .B1(_04951_),
    .C1(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__or2_4 _11774_ (.A(_04870_),
    .B(_04950_),
    .X(_04964_));
 sky130_fd_sc_hd__buf_6 _11775_ (.A(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__mux2_1 _11776_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04924_),
    .X(_04966_));
 sky130_fd_sc_hd__mux2_1 _11777_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04924_),
    .X(_04967_));
 sky130_fd_sc_hd__mux2_1 _11778_ (.A0(_04966_),
    .A1(_04967_),
    .S(_04910_),
    .X(_04968_));
 sky130_fd_sc_hd__mux2_1 _11779_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04919_),
    .X(_04969_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04894_),
    .X(_04970_));
 sky130_fd_sc_hd__or2_1 _11781_ (.A(_04928_),
    .B(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__o211a_1 _11782_ (.A1(_04922_),
    .A2(_04969_),
    .B1(_04971_),
    .C1(_04931_),
    .X(_04972_));
 sky130_fd_sc_hd__a211o_1 _11783_ (.A1(_04946_),
    .A2(_04968_),
    .B1(_04972_),
    .C1(_04884_),
    .X(_04973_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04924_),
    .X(_04974_));
 sky130_fd_sc_hd__mux2_1 _11785_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04924_),
    .X(_04975_));
 sky130_fd_sc_hd__mux2_1 _11786_ (.A0(_04974_),
    .A1(_04975_),
    .S(_04910_),
    .X(_04976_));
 sky130_fd_sc_hd__mux2_1 _11787_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04924_),
    .X(_04977_));
 sky130_fd_sc_hd__and3_1 _11788_ (.A(\rbzero.tex_r0[43] ),
    .B(_04892_),
    .C(_04893_),
    .X(_04978_));
 sky130_fd_sc_hd__a21o_1 _11789_ (.A1(\rbzero.tex_r0[42] ),
    .A2(_04939_),
    .B1(_04941_),
    .X(_04979_));
 sky130_fd_sc_hd__o221a_1 _11790_ (.A1(_04922_),
    .A2(_04977_),
    .B1(_04978_),
    .B2(_04979_),
    .C1(_04945_),
    .X(_04980_));
 sky130_fd_sc_hd__a211o_1 _11791_ (.A1(_04932_),
    .A2(_04976_),
    .B1(_04980_),
    .C1(_04908_),
    .X(_04981_));
 sky130_fd_sc_hd__and3_1 _11792_ (.A(_04859_),
    .B(_04864_),
    .C(_04862_),
    .X(_04982_));
 sky130_fd_sc_hd__a21o_1 _11793_ (.A1(_04864_),
    .A2(_04862_),
    .B1(_04859_),
    .X(_04983_));
 sky130_fd_sc_hd__or3b_1 _11794_ (.A(_04870_),
    .B(_04982_),
    .C_N(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__clkbuf_16 _11795_ (.A(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__a31o_1 _11796_ (.A1(_04965_),
    .A2(_04973_),
    .A3(_04981_),
    .B1(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__buf_6 _11797_ (.A(_04908_),
    .X(_04987_));
 sky130_fd_sc_hd__and2_1 _11798_ (.A(\rbzero.tex_r0[12] ),
    .B(_04920_),
    .X(_04988_));
 sky130_fd_sc_hd__a31o_1 _11799_ (.A1(\rbzero.tex_r0[13] ),
    .A2(_04892_),
    .A3(_04893_),
    .B1(_04922_),
    .X(_04989_));
 sky130_fd_sc_hd__mux2_1 _11800_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04925_),
    .X(_04990_));
 sky130_fd_sc_hd__buf_4 _11801_ (.A(_04942_),
    .X(_04991_));
 sky130_fd_sc_hd__o221a_1 _11802_ (.A1(_04988_),
    .A2(_04989_),
    .B1(_04990_),
    .B2(_04991_),
    .C1(_04932_),
    .X(_04992_));
 sky130_fd_sc_hd__mux2_1 _11803_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04925_),
    .X(_04993_));
 sky130_fd_sc_hd__and3_1 _11804_ (.A(\rbzero.tex_r0[11] ),
    .B(_04936_),
    .C(_04937_),
    .X(_04994_));
 sky130_fd_sc_hd__clkbuf_8 _11805_ (.A(_04941_),
    .X(_04995_));
 sky130_fd_sc_hd__a21o_1 _11806_ (.A1(\rbzero.tex_r0[10] ),
    .A2(_04940_),
    .B1(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__o221a_1 _11807_ (.A1(_04934_),
    .A2(_04993_),
    .B1(_04994_),
    .B2(_04996_),
    .C1(_04952_),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04919_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_04919_),
    .X(_04999_));
 sky130_fd_sc_hd__mux2_1 _11810_ (.A0(_04998_),
    .A1(_04999_),
    .S(_04922_),
    .X(_05000_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04939_),
    .X(_05001_));
 sky130_fd_sc_hd__mux2_1 _11812_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04895_),
    .X(_05002_));
 sky130_fd_sc_hd__or2_1 _11813_ (.A(_04941_),
    .B(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__o211a_1 _11814_ (.A1(_04956_),
    .A2(_05001_),
    .B1(_05003_),
    .C1(_04960_),
    .X(_05004_));
 sky130_fd_sc_hd__a211o_1 _11815_ (.A1(_04952_),
    .A2(_05000_),
    .B1(_05004_),
    .C1(_04918_),
    .X(_05005_));
 sky130_fd_sc_hd__o311a_1 _11816_ (.A1(_04987_),
    .A2(_04992_),
    .A3(_04997_),
    .B1(_04965_),
    .C1(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04919_),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_1 _11818_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04924_),
    .X(_05008_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(_05007_),
    .A1(_05008_),
    .S(_04910_),
    .X(_05009_));
 sky130_fd_sc_hd__and2_1 _11820_ (.A(\rbzero.tex_r0[20] ),
    .B(_04939_),
    .X(_05010_));
 sky130_fd_sc_hd__a31o_1 _11821_ (.A1(\rbzero.tex_r0[21] ),
    .A2(_04892_),
    .A3(_04893_),
    .B1(_04873_),
    .X(_05011_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04919_),
    .X(_05012_));
 sky130_fd_sc_hd__o221a_1 _11823_ (.A1(_05010_),
    .A2(_05011_),
    .B1(_05012_),
    .B2(_04942_),
    .C1(_04931_),
    .X(_05013_));
 sky130_fd_sc_hd__a211o_1 _11824_ (.A1(_04952_),
    .A2(_05009_),
    .B1(_05013_),
    .C1(_04884_),
    .X(_05014_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04924_),
    .X(_05015_));
 sky130_fd_sc_hd__mux2_1 _11826_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04924_),
    .X(_05016_));
 sky130_fd_sc_hd__mux2_1 _11827_ (.A0(_05015_),
    .A1(_05016_),
    .S(_04910_),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04919_),
    .X(_05018_));
 sky130_fd_sc_hd__mux2_1 _11829_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04894_),
    .X(_05019_));
 sky130_fd_sc_hd__or2_1 _11830_ (.A(_04928_),
    .B(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__o211a_1 _11831_ (.A1(_04956_),
    .A2(_05018_),
    .B1(_05020_),
    .C1(_04931_),
    .X(_05021_));
 sky130_fd_sc_hd__a211o_1 _11832_ (.A1(_04952_),
    .A2(_05017_),
    .B1(_05021_),
    .C1(_04908_),
    .X(_05022_));
 sky130_fd_sc_hd__inv_4 _11833_ (.A(_04985_),
    .Y(_05023_));
 sky130_fd_sc_hd__a31o_1 _11834_ (.A1(_04951_),
    .A2(_05014_),
    .A3(_05022_),
    .B1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__o221a_1 _11835_ (.A1(_04963_),
    .A2(_04986_),
    .B1(_05006_),
    .B2(_05024_),
    .C1(_04906_),
    .X(_05025_));
 sky130_fd_sc_hd__a31o_1 _11836_ (.A1(_04904_),
    .A2(_04907_),
    .A3(_04917_),
    .B1(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__buf_4 _11837_ (.A(_04928_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_8 _11838_ (.A(_04944_),
    .X(_05028_));
 sky130_fd_sc_hd__o211a_1 _11839_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_04928_),
    .B1(_04939_),
    .C1(\rbzero.floor_leak[0] ),
    .X(_05029_));
 sky130_fd_sc_hd__a221o_1 _11840_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_05027_),
    .B1(_05028_),
    .B2(\rbzero.floor_leak[2] ),
    .C1(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__o221a_1 _11841_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04908_),
    .B1(_04945_),
    .B2(\rbzero.floor_leak[2] ),
    .C1(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__a221o_1 _11842_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04987_),
    .B1(_04964_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__o221a_2 _11843_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_04985_),
    .B1(_04965_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__nand2_1 _11844_ (.A(_04908_),
    .B(_04876_),
    .Y(_05034_));
 sky130_fd_sc_hd__buf_4 _11845_ (.A(_04878_),
    .X(_05035_));
 sky130_fd_sc_hd__clkbuf_4 _11846_ (.A(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__or3_1 _11847_ (.A(_04922_),
    .B(_05036_),
    .C(_05023_),
    .X(_05037_));
 sky130_fd_sc_hd__or4_1 _11848_ (.A(_05034_),
    .B(_04951_),
    .C(_04808_),
    .D(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__inv_2 _11849_ (.A(\rbzero.row_render.size[2] ),
    .Y(_05039_));
 sky130_fd_sc_hd__nor2_1 _11850_ (.A(\rbzero.row_render.size[1] ),
    .B(\rbzero.row_render.size[0] ),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_1 _11851_ (.A(_05039_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__or2_1 _11852_ (.A(\rbzero.row_render.size[3] ),
    .B(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__or3_1 _11853_ (.A(\rbzero.row_render.size[5] ),
    .B(\rbzero.row_render.size[4] ),
    .C(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__and2_1 _11854_ (.A(\rbzero.row_render.size[6] ),
    .B(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__o21a_1 _11855_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_05044_),
    .B1(\rbzero.row_render.size[8] ),
    .X(_05045_));
 sky130_fd_sc_hd__a21oi_1 _11856_ (.A1(\rbzero.row_render.size[7] ),
    .A2(\rbzero.row_render.size[6] ),
    .B1(\rbzero.row_render.size[8] ),
    .Y(_05046_));
 sky130_fd_sc_hd__xnor2_1 _11857_ (.A(\rbzero.row_render.size[7] ),
    .B(\rbzero.row_render.size[6] ),
    .Y(_05047_));
 sky130_fd_sc_hd__and3_1 _11858_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(\rbzero.row_render.size[6] ),
    .X(_05048_));
 sky130_fd_sc_hd__nor2_1 _11859_ (.A(_05046_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__and2_1 _11860_ (.A(\rbzero.row_render.size[1] ),
    .B(_04633_),
    .X(_05050_));
 sky130_fd_sc_hd__o22a_1 _11861_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_04639_),
    .B1(_04633_),
    .B2(\rbzero.row_render.size[1] ),
    .X(_05051_));
 sky130_fd_sc_hd__o31a_1 _11862_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_04111_),
    .A3(_05050_),
    .B1(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__a221o_1 _11863_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_04475_),
    .B1(_04639_),
    .B2(\rbzero.row_render.size[2] ),
    .C1(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__o221a_1 _11864_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_04476_),
    .B1(_04477_),
    .B2(\rbzero.row_render.size[4] ),
    .C1(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__a221o_1 _11865_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_04801_),
    .B1(_04477_),
    .B2(\rbzero.row_render.size[4] ),
    .C1(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__o2bb2a_1 _11866_ (.A1_N(\rbzero.row_render.size[6] ),
    .A2_N(_04479_),
    .B1(_04801_),
    .B2(\rbzero.row_render.size[5] ),
    .X(_05056_));
 sky130_fd_sc_hd__nand2_1 _11867_ (.A(_05055_),
    .B(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__o221a_1 _11868_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_04479_),
    .B1(_05047_),
    .B2(_04031_),
    .C1(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__a221o_1 _11869_ (.A1(_04031_),
    .A2(_05047_),
    .B1(_05049_),
    .B2(\gpout0.hpos[8] ),
    .C1(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__and2b_1 _11870_ (.A_N(\rbzero.row_render.size[9] ),
    .B(\gpout0.hpos[9] ),
    .X(_05060_));
 sky130_fd_sc_hd__or2b_1 _11871_ (.A(\gpout0.hpos[9] ),
    .B_N(\rbzero.row_render.size[9] ),
    .X(_05061_));
 sky130_fd_sc_hd__o221a_1 _11872_ (.A1(\gpout0.hpos[8] ),
    .A2(_05049_),
    .B1(_05060_),
    .B2(_05046_),
    .C1(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__xnor2_1 _11873_ (.A(\rbzero.row_render.size[7] ),
    .B(_05044_),
    .Y(_05063_));
 sky130_fd_sc_hd__nor3_1 _11874_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(_05044_),
    .Y(_05064_));
 sky130_fd_sc_hd__nor2_1 _11875_ (.A(_05045_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__nor2_1 _11876_ (.A(\rbzero.row_render.size[6] ),
    .B(_05043_),
    .Y(_05066_));
 sky130_fd_sc_hd__nor2_1 _11877_ (.A(_05044_),
    .B(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__o21ai_1 _11878_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_05042_),
    .B1(\rbzero.row_render.size[5] ),
    .Y(_05068_));
 sky130_fd_sc_hd__nand2_1 _11879_ (.A(_05043_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__xnor2_1 _11880_ (.A(\rbzero.row_render.size[4] ),
    .B(_05042_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2_1 _11881_ (.A(\rbzero.row_render.size[3] ),
    .B(_05041_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _11882_ (.A(_05042_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__or2_1 _11883_ (.A(_05039_),
    .B(_05040_),
    .X(_05073_));
 sky130_fd_sc_hd__nand2_1 _11884_ (.A(_05041_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__or2_1 _11885_ (.A(\rbzero.row_render.size[0] ),
    .B(_04507_),
    .X(_05075_));
 sky130_fd_sc_hd__a31o_1 _11886_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_04509_),
    .A3(_05075_),
    .B1(_05040_),
    .X(_05076_));
 sky130_fd_sc_hd__a211o_1 _11887_ (.A1(\rbzero.row_render.size[2] ),
    .A2(\gpout0.hpos[2] ),
    .B1(_04707_),
    .C1(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__o221a_1 _11888_ (.A1(_04471_),
    .A2(_05072_),
    .B1(_05074_),
    .B2(\gpout0.hpos[2] ),
    .C1(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__a221o_1 _11889_ (.A1(_04471_),
    .A2(_05072_),
    .B1(_05070_),
    .B2(\gpout0.hpos[4] ),
    .C1(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__o221a_1 _11890_ (.A1(_04642_),
    .A2(_05070_),
    .B1(_05069_),
    .B2(\gpout0.hpos[5] ),
    .C1(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__a221o_1 _11891_ (.A1(_04473_),
    .A2(_05069_),
    .B1(_05067_),
    .B2(_04479_),
    .C1(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__o221a_1 _11892_ (.A1(_04479_),
    .A2(_05067_),
    .B1(_05063_),
    .B2(\gpout0.hpos[7] ),
    .C1(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__a221o_1 _11893_ (.A1(_04031_),
    .A2(_05063_),
    .B1(_05065_),
    .B2(\gpout0.hpos[8] ),
    .C1(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__or2_1 _11894_ (.A(\gpout0.hpos[8] ),
    .B(_05065_),
    .X(_05084_));
 sky130_fd_sc_hd__a21oi_1 _11895_ (.A1(_05083_),
    .A2(_05084_),
    .B1(\gpout0.hpos[9] ),
    .Y(_05085_));
 sky130_fd_sc_hd__a221o_1 _11896_ (.A1(\gpout0.hpos[9] ),
    .A2(_05046_),
    .B1(_05059_),
    .B2(_05062_),
    .C1(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__or4b_2 _11897_ (.A(\rbzero.row_render.size[10] ),
    .B(\rbzero.row_render.size[9] ),
    .C(_05045_),
    .D_N(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__a21oi_1 _11898_ (.A1(_05038_),
    .A2(_05087_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_05088_));
 sky130_fd_sc_hd__a21o_2 _11899_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_04985_),
    .B1(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__nor2_2 _11900_ (.A(_05033_),
    .B(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__mux2_1 _11901_ (.A0(_04809_),
    .A1(_05026_),
    .S(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__nor3_2 _11902_ (.A(_04759_),
    .B(_04760_),
    .C(_04763_),
    .Y(_05092_));
 sky130_fd_sc_hd__o22a_1 _11903_ (.A1(_04765_),
    .A2(_04807_),
    .B1(_05091_),
    .B2(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__nor2_1 _11904_ (.A(_04720_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__and3_2 _11905_ (.A(\rbzero.trace_state[3] ),
    .B(_04486_),
    .C(_04493_),
    .X(_05095_));
 sky130_fd_sc_hd__a21o_1 _11906_ (.A1(_04494_),
    .A2(_05095_),
    .B1(_04695_),
    .X(_05096_));
 sky130_fd_sc_hd__o21ai_1 _11907_ (.A1(_04721_),
    .A2(_05094_),
    .B1(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__o21a_4 _11908_ (.A1(\gpout0.hpos[7] ),
    .A2(\gpout0.hpos[8] ),
    .B1(\gpout0.hpos[9] ),
    .X(_05098_));
 sky130_fd_sc_hd__and3_1 _11909_ (.A(_04714_),
    .B(_04718_),
    .C(_04699_),
    .X(_05099_));
 sky130_fd_sc_hd__a21o_4 _11910_ (.A1(\gpout0.vpos[8] ),
    .A2(_05099_),
    .B1(\gpout0.vpos[9] ),
    .X(_05100_));
 sky130_fd_sc_hd__nor2_2 _11911_ (.A(_05098_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__o211a_2 _11912_ (.A1(_04494_),
    .A2(_04695_),
    .B1(_05097_),
    .C1(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__buf_4 _11913_ (.A(net45),
    .X(_05103_));
 sky130_fd_sc_hd__mux2_4 _11914_ (.A0(\reg_rgb[6] ),
    .A1(_05102_),
    .S(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__clkbuf_1 _11915_ (.A(_05104_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 _11916_ (.A(_04474_),
    .X(_05105_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_05105_),
    .B(_04035_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand2_2 _11918_ (.A(_04472_),
    .B(_04696_),
    .Y(_05107_));
 sky130_fd_sc_hd__xnor2_4 _11919_ (.A(_04514_),
    .B(_05107_),
    .Y(_05108_));
 sky130_fd_sc_hd__or2_1 _11920_ (.A(_04471_),
    .B(_04696_),
    .X(_05109_));
 sky130_fd_sc_hd__or2b_1 _11921_ (.A(_04709_),
    .B_N(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__and2_1 _11922_ (.A(_04501_),
    .B(_04711_),
    .X(_05111_));
 sky130_fd_sc_hd__or2_1 _11923_ (.A(_04712_),
    .B(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__inv_2 _11924_ (.A(_05108_),
    .Y(_05113_));
 sky130_fd_sc_hd__or3_1 _11925_ (.A(_04479_),
    .B(\gpout0.hpos[5] ),
    .C(_04710_),
    .X(_05114_));
 sky130_fd_sc_hd__o2bb2a_1 _11926_ (.A1_N(_04711_),
    .A2_N(_05114_),
    .B1(_05110_),
    .B2(\gpout0.hpos[4] ),
    .X(_05115_));
 sky130_fd_sc_hd__or3b_1 _11927_ (.A(_05112_),
    .B(_05113_),
    .C_N(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__or3b_1 _11928_ (.A(_04713_),
    .B(_05098_),
    .C_N(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__nor2_1 _11929_ (.A(_05110_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__and2_1 _11930_ (.A(_04477_),
    .B(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__o41a_2 _11931_ (.A1(_04479_),
    .A2(\gpout0.hpos[5] ),
    .A3(_04710_),
    .A4(_05109_),
    .B1(\gpout0.hpos[7] ),
    .X(_05120_));
 sky130_fd_sc_hd__xor2_4 _11932_ (.A(\gpout0.hpos[8] ),
    .B(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__xor2_2 _11933_ (.A(_05116_),
    .B(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__and4b_1 _11934_ (.A_N(_04473_),
    .B(_05108_),
    .C(_05119_),
    .D(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__nand2_2 _11935_ (.A(_05108_),
    .B(_05122_),
    .Y(_05124_));
 sky130_fd_sc_hd__a21bo_1 _11936_ (.A1(_04478_),
    .A2(_04696_),
    .B1_N(_04710_),
    .X(_05125_));
 sky130_fd_sc_hd__or2b_1 _11937_ (.A(_05117_),
    .B_N(_05110_),
    .X(_05126_));
 sky130_fd_sc_hd__or3_1 _11938_ (.A(_04473_),
    .B(_05125_),
    .C(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__nor2_1 _11939_ (.A(_05124_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__a31o_1 _11940_ (.A1(_04471_),
    .A2(_04642_),
    .A3(_04696_),
    .B1(\gpout0.hpos[5] ),
    .X(_05129_));
 sky130_fd_sc_hd__nand2_1 _11941_ (.A(_05107_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__and3_1 _11942_ (.A(_04642_),
    .B(_05118_),
    .C(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__and3_1 _11943_ (.A(_05108_),
    .B(_05131_),
    .C(_05122_),
    .X(_05132_));
 sky130_fd_sc_hd__or3_1 _11944_ (.A(_05123_),
    .B(_05128_),
    .C(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__and2b_1 _11945_ (.A_N(_05126_),
    .B(_05125_),
    .X(_05134_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(_05130_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__nor2_1 _11947_ (.A(_05124_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__or4_2 _11948_ (.A(_04477_),
    .B(_05110_),
    .C(_05117_),
    .D(_05130_),
    .X(_05137_));
 sky130_fd_sc_hd__nor2_1 _11949_ (.A(_05125_),
    .B(_05126_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_1 _11950_ (.A(_04473_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__o21ai_1 _11951_ (.A1(_05138_),
    .A2(_05131_),
    .B1(_05113_),
    .Y(_05140_));
 sky130_fd_sc_hd__and3_1 _11952_ (.A(_05107_),
    .B(_05129_),
    .C(_05134_),
    .X(_05141_));
 sky130_fd_sc_hd__and3_1 _11953_ (.A(_04479_),
    .B(_04473_),
    .C(_05119_),
    .X(_05142_));
 sky130_fd_sc_hd__a21oi_1 _11954_ (.A1(_04480_),
    .A2(_05141_),
    .B1(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__nand2_1 _11955_ (.A(_04479_),
    .B(\gpout0.hpos[5] ),
    .Y(_05144_));
 sky130_fd_sc_hd__mux2_1 _11956_ (.A0(_05144_),
    .A1(_05108_),
    .S(_05115_),
    .X(_05145_));
 sky130_fd_sc_hd__or2_1 _11957_ (.A(_05112_),
    .B(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__nand2_1 _11958_ (.A(_05112_),
    .B(_05145_),
    .Y(_05147_));
 sky130_fd_sc_hd__nand2_1 _11959_ (.A(_05146_),
    .B(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__a41o_1 _11960_ (.A1(_05137_),
    .A2(_05139_),
    .A3(_05140_),
    .A4(_05143_),
    .B1(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__or3b_4 _11961_ (.A(_05133_),
    .B(_05136_),
    .C_N(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__and3_2 _11962_ (.A(_05108_),
    .B(_05141_),
    .C(_05122_),
    .X(_05151_));
 sky130_fd_sc_hd__nor2_4 _11963_ (.A(_05137_),
    .B(_05124_),
    .Y(_05152_));
 sky130_fd_sc_hd__clkbuf_4 _11964_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_05153_));
 sky130_fd_sc_hd__and4bb_2 _11965_ (.A_N(_04473_),
    .B_N(_05121_),
    .C(_05119_),
    .D(_05113_),
    .X(_05154_));
 sky130_fd_sc_hd__nor3_4 _11966_ (.A(_05108_),
    .B(_05121_),
    .C(_05135_),
    .Y(_05155_));
 sky130_fd_sc_hd__a21o_1 _11967_ (.A1(_05146_),
    .A2(_05147_),
    .B1(_05121_),
    .X(_05156_));
 sky130_fd_sc_hd__inv_2 _11968_ (.A(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__and2_2 _11969_ (.A(_05142_),
    .B(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__a22o_1 _11970_ (.A1(\rbzero.debug_overlay.vplaneX[-4] ),
    .A2(_05155_),
    .B1(_05158_),
    .B2(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_05159_));
 sky130_fd_sc_hd__a211o_1 _11971_ (.A1(_05153_),
    .A2(_05154_),
    .B1(_05159_),
    .C1(_04723_),
    .X(_05160_));
 sky130_fd_sc_hd__a221o_1 _11972_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_05151_),
    .B1(_05152_),
    .B2(\rbzero.debug_overlay.vplaneX[-3] ),
    .C1(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__nor2_1 _11973_ (.A(_05108_),
    .B(_05156_),
    .Y(_05162_));
 sky130_fd_sc_hd__and2b_2 _11974_ (.A_N(_05127_),
    .B(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__and2_2 _11975_ (.A(_05131_),
    .B(_05162_),
    .X(_05164_));
 sky130_fd_sc_hd__and3_2 _11976_ (.A(_04480_),
    .B(_05141_),
    .C(_05157_),
    .X(_05165_));
 sky130_fd_sc_hd__a22o_1 _11977_ (.A1(\rbzero.debug_overlay.vplaneX[-7] ),
    .A2(_05164_),
    .B1(_05165_),
    .B2(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_05166_));
 sky130_fd_sc_hd__and4_2 _11978_ (.A(_04473_),
    .B(_05108_),
    .C(_05119_),
    .D(_05122_),
    .X(_05167_));
 sky130_fd_sc_hd__nor2_4 _11979_ (.A(_05139_),
    .B(_05124_),
    .Y(_05168_));
 sky130_fd_sc_hd__a22o_1 _11980_ (.A1(\rbzero.debug_overlay.vplaneX[-1] ),
    .A2(_05167_),
    .B1(_05168_),
    .B2(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_05169_));
 sky130_fd_sc_hd__a211o_1 _11981_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(_05163_),
    .B1(_05166_),
    .C1(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__a211oi_1 _11982_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_05150_),
    .B1(_05161_),
    .C1(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__buf_4 _11983_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_4 _11984_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_05173_));
 sky130_fd_sc_hd__a21bo_1 _11985_ (.A1(_05173_),
    .A2(_05154_),
    .B1_N(\gpout0.vpos[3] ),
    .X(_05174_));
 sky130_fd_sc_hd__a221o_1 _11986_ (.A1(\rbzero.debug_overlay.vplaneY[-4] ),
    .A2(_05155_),
    .B1(_05158_),
    .B2(_05172_),
    .C1(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__a221o_1 _11987_ (.A1(\rbzero.debug_overlay.vplaneY[0] ),
    .A2(_05151_),
    .B1(_05152_),
    .B2(\rbzero.debug_overlay.vplaneY[-3] ),
    .C1(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_4 _11988_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_05177_));
 sky130_fd_sc_hd__a22o_1 _11989_ (.A1(\rbzero.debug_overlay.vplaneY[-7] ),
    .A2(_05164_),
    .B1(_05163_),
    .B2(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_05178_));
 sky130_fd_sc_hd__a21o_1 _11990_ (.A1(\rbzero.debug_overlay.vplaneY[-8] ),
    .A2(_05165_),
    .B1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__a221o_1 _11991_ (.A1(\rbzero.debug_overlay.vplaneY[-1] ),
    .A2(_05167_),
    .B1(_05168_),
    .B2(_05177_),
    .C1(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__a211o_1 _11992_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(_05150_),
    .B1(_05176_),
    .C1(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__or3b_1 _11993_ (.A(_04705_),
    .B(_05171_),
    .C_N(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__or2_2 _11994_ (.A(_04699_),
    .B(_04703_),
    .X(_05183_));
 sky130_fd_sc_hd__a22o_1 _11995_ (.A1(\rbzero.debug_overlay.facingY[-1] ),
    .A2(_05167_),
    .B1(_05165_),
    .B2(\rbzero.debug_overlay.facingY[-8] ),
    .X(_05184_));
 sky130_fd_sc_hd__a22o_1 _11996_ (.A1(\rbzero.debug_overlay.facingY[-4] ),
    .A2(_05155_),
    .B1(_05158_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .X(_05185_));
 sky130_fd_sc_hd__a22o_1 _11997_ (.A1(\rbzero.debug_overlay.facingY[-7] ),
    .A2(_05164_),
    .B1(_05152_),
    .B2(\rbzero.debug_overlay.facingY[-3] ),
    .X(_05186_));
 sky130_fd_sc_hd__a221o_1 _11998_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_05163_),
    .B1(_05168_),
    .B2(\rbzero.debug_overlay.facingY[-2] ),
    .C1(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__a211o_1 _11999_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_05154_),
    .B1(_05185_),
    .C1(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__a211o_1 _12000_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_05151_),
    .B1(_05184_),
    .C1(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__a21oi_1 _12001_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_05150_),
    .B1(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__or3_1 _12002_ (.A(_04729_),
    .B(_04702_),
    .C(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__a22o_1 _12003_ (.A1(\rbzero.debug_overlay.facingX[-7] ),
    .A2(_05164_),
    .B1(_05152_),
    .B2(\rbzero.debug_overlay.facingX[-3] ),
    .X(_05192_));
 sky130_fd_sc_hd__a22o_1 _12004_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_05155_),
    .B1(_05154_),
    .B2(\rbzero.debug_overlay.facingX[-5] ),
    .X(_05193_));
 sky130_fd_sc_hd__a22o_1 _12005_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(_05167_),
    .B1(_05168_),
    .B2(\rbzero.debug_overlay.facingX[-2] ),
    .X(_05194_));
 sky130_fd_sc_hd__a221o_1 _12006_ (.A1(\rbzero.debug_overlay.facingX[0] ),
    .A2(_05151_),
    .B1(_05163_),
    .B2(\rbzero.debug_overlay.facingX[-6] ),
    .C1(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__a2111o_1 _12007_ (.A1(\rbzero.debug_overlay.facingX[-9] ),
    .A2(_05158_),
    .B1(_05183_),
    .C1(_05193_),
    .D1(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__a211o_1 _12008_ (.A1(\rbzero.debug_overlay.facingX[-8] ),
    .A2(_05165_),
    .B1(_05192_),
    .C1(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__a21oi_1 _12009_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_05150_),
    .B1(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__a31oi_2 _12010_ (.A1(_05182_),
    .A2(_05183_),
    .A3(_05191_),
    .B1(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__a22o_1 _12011_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_05151_),
    .B1(_05152_),
    .B2(\rbzero.debug_overlay.playerX[-3] ),
    .X(_05200_));
 sky130_fd_sc_hd__a221o_1 _12012_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_05164_),
    .B1(_05168_),
    .B2(\rbzero.debug_overlay.playerX[-2] ),
    .C1(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__a22o_1 _12013_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_05167_),
    .B1(_05163_),
    .B2(\rbzero.debug_overlay.playerX[-6] ),
    .X(_05202_));
 sky130_fd_sc_hd__a22o_1 _12014_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_05128_),
    .B1(_05132_),
    .B2(\rbzero.debug_overlay.playerX[1] ),
    .X(_05203_));
 sky130_fd_sc_hd__a221o_1 _12015_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_05154_),
    .B1(_05158_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__nor2_1 _12016_ (.A(_05148_),
    .B(_05137_),
    .Y(_05205_));
 sky130_fd_sc_hd__a221o_1 _12017_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_05136_),
    .B1(_05205_),
    .B2(\rbzero.debug_overlay.playerX[5] ),
    .C1(_04717_),
    .X(_05206_));
 sky130_fd_sc_hd__a221o_1 _12018_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_05155_),
    .B1(_05165_),
    .B2(\rbzero.debug_overlay.playerX[-8] ),
    .C1(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__a2111o_1 _12019_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_05123_),
    .B1(_05202_),
    .C1(_05204_),
    .D1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__or2_1 _12020_ (.A(_05201_),
    .B(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__nand2_1 _12021_ (.A(\gpout0.vpos[3] ),
    .B(_04700_),
    .Y(_05210_));
 sky130_fd_sc_hd__a221o_1 _12022_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_05155_),
    .B1(_05205_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .C1(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__a221o_1 _12023_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_05154_),
    .B1(_05158_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .C1(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__a22o_1 _12024_ (.A1(_04734_),
    .A2(_05132_),
    .B1(_05152_),
    .B2(\rbzero.debug_overlay.playerY[-3] ),
    .X(_05213_));
 sky130_fd_sc_hd__a221o_1 _12025_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_05128_),
    .B1(_05136_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .C1(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__a22o_1 _12026_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_05151_),
    .B1(_05165_),
    .B2(\rbzero.debug_overlay.playerY[-8] ),
    .X(_05215_));
 sky130_fd_sc_hd__a22o_1 _12027_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_05164_),
    .B1(_05167_),
    .B2(\rbzero.debug_overlay.playerY[-1] ),
    .X(_05216_));
 sky130_fd_sc_hd__a221o_1 _12028_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_05123_),
    .B1(_05168_),
    .B2(\rbzero.debug_overlay.playerY[-2] ),
    .C1(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__a211o_1 _12029_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_05163_),
    .B1(_05215_),
    .C1(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__or3_1 _12030_ (.A(_05212_),
    .B(_05214_),
    .C(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__and4_1 _12031_ (.A(_04708_),
    .B(_04697_),
    .C(_05209_),
    .D(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__o21ai_1 _12032_ (.A1(_04700_),
    .A2(_05199_),
    .B1(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__o311a_1 _12033_ (.A1(_04708_),
    .A2(_04762_),
    .A3(_05106_),
    .B1(_05221_),
    .C1(_04720_),
    .X(_05222_));
 sky130_fd_sc_hd__buf_6 _12034_ (.A(_04918_),
    .X(_05223_));
 sky130_fd_sc_hd__clkbuf_4 _12035_ (.A(_04991_),
    .X(_05224_));
 sky130_fd_sc_hd__buf_4 _12036_ (.A(_04896_),
    .X(_05225_));
 sky130_fd_sc_hd__buf_4 _12037_ (.A(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__buf_4 _12038_ (.A(_04879_),
    .X(_05227_));
 sky130_fd_sc_hd__or2_1 _12039_ (.A(\rbzero.tex_r1[14] ),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__buf_4 _12040_ (.A(_04934_),
    .X(_05229_));
 sky130_fd_sc_hd__o211a_1 _12041_ (.A1(\rbzero.tex_r1[15] ),
    .A2(_05226_),
    .B1(_05228_),
    .C1(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__clkbuf_4 _12042_ (.A(_05027_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_4 _12043_ (.A(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__clkbuf_4 _12044_ (.A(_05227_),
    .X(_05233_));
 sky130_fd_sc_hd__a31o_1 _12045_ (.A1(\rbzero.tex_r1[13] ),
    .A2(_05232_),
    .A3(_05233_),
    .B1(_04952_),
    .X(_05234_));
 sky130_fd_sc_hd__a311o_1 _12046_ (.A1(\rbzero.tex_r1[12] ),
    .A2(_05224_),
    .A3(_04899_),
    .B1(_05230_),
    .C1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__or2_1 _12047_ (.A(\rbzero.tex_r1[10] ),
    .B(_05227_),
    .X(_05236_));
 sky130_fd_sc_hd__o211a_1 _12048_ (.A1(\rbzero.tex_r1[11] ),
    .A2(_05226_),
    .B1(_05236_),
    .C1(_05229_),
    .X(_05237_));
 sky130_fd_sc_hd__buf_6 _12049_ (.A(_04960_),
    .X(_05238_));
 sky130_fd_sc_hd__a31o_1 _12050_ (.A1(\rbzero.tex_r1[9] ),
    .A2(_05232_),
    .A3(_05233_),
    .B1(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__a311o_1 _12051_ (.A1(\rbzero.tex_r1[8] ),
    .A2(_05224_),
    .A3(_04899_),
    .B1(_05237_),
    .C1(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__buf_6 _12052_ (.A(_04951_),
    .X(_05241_));
 sky130_fd_sc_hd__buf_4 _12053_ (.A(_04940_),
    .X(_05242_));
 sky130_fd_sc_hd__clkbuf_4 _12054_ (.A(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_4 _12055_ (.A(_05035_),
    .X(_05244_));
 sky130_fd_sc_hd__clkbuf_4 _12056_ (.A(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__or2_1 _12057_ (.A(\rbzero.tex_r1[6] ),
    .B(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__o211a_1 _12058_ (.A1(\rbzero.tex_r1[7] ),
    .A2(_05243_),
    .B1(_05246_),
    .C1(_05229_),
    .X(_05247_));
 sky130_fd_sc_hd__a31o_1 _12059_ (.A1(\rbzero.tex_r1[5] ),
    .A2(_04930_),
    .A3(_05245_),
    .B1(_04946_),
    .X(_05248_));
 sky130_fd_sc_hd__a31o_1 _12060_ (.A1(\rbzero.tex_r1[4] ),
    .A2(_05224_),
    .A3(_04899_),
    .B1(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__or2_1 _12061_ (.A(\rbzero.tex_r1[2] ),
    .B(_05245_),
    .X(_05250_));
 sky130_fd_sc_hd__o211a_1 _12062_ (.A1(\rbzero.tex_r1[3] ),
    .A2(_04899_),
    .B1(_05250_),
    .C1(_05229_),
    .X(_05251_));
 sky130_fd_sc_hd__a31o_1 _12063_ (.A1(\rbzero.tex_r1[1] ),
    .A2(_04991_),
    .A3(_05233_),
    .B1(_04932_),
    .X(_05252_));
 sky130_fd_sc_hd__a31o_1 _12064_ (.A1(\rbzero.tex_r1[0] ),
    .A2(_05224_),
    .A3(_04899_),
    .B1(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__buf_4 _12065_ (.A(_04908_),
    .X(_05254_));
 sky130_fd_sc_hd__o221a_1 _12066_ (.A1(_05247_),
    .A2(_05249_),
    .B1(_05251_),
    .B2(_05253_),
    .C1(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__a311o_1 _12067_ (.A1(_05223_),
    .A2(_05235_),
    .A3(_05240_),
    .B1(_05241_),
    .C1(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__or2_1 _12068_ (.A(\rbzero.tex_r1[30] ),
    .B(_05227_),
    .X(_05257_));
 sky130_fd_sc_hd__o211a_1 _12069_ (.A1(\rbzero.tex_r1[31] ),
    .A2(_05226_),
    .B1(_05257_),
    .C1(_05229_),
    .X(_05258_));
 sky130_fd_sc_hd__a31o_1 _12070_ (.A1(\rbzero.tex_r1[29] ),
    .A2(_05232_),
    .A3(_05233_),
    .B1(_04952_),
    .X(_05259_));
 sky130_fd_sc_hd__a311o_1 _12071_ (.A1(\rbzero.tex_r1[28] ),
    .A2(_05224_),
    .A3(_04899_),
    .B1(_05258_),
    .C1(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__or2_1 _12072_ (.A(\rbzero.tex_r1[26] ),
    .B(_05227_),
    .X(_05261_));
 sky130_fd_sc_hd__o211a_1 _12073_ (.A1(\rbzero.tex_r1[27] ),
    .A2(_05226_),
    .B1(_05261_),
    .C1(_05229_),
    .X(_05262_));
 sky130_fd_sc_hd__buf_4 _12074_ (.A(_04995_),
    .X(_05263_));
 sky130_fd_sc_hd__a31o_1 _12075_ (.A1(\rbzero.tex_r1[25] ),
    .A2(_05263_),
    .A3(_05233_),
    .B1(_05238_),
    .X(_05264_));
 sky130_fd_sc_hd__a311o_1 _12076_ (.A1(\rbzero.tex_r1[24] ),
    .A2(_05224_),
    .A3(_04899_),
    .B1(_05262_),
    .C1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__or2_1 _12077_ (.A(\rbzero.tex_r1[22] ),
    .B(_05227_),
    .X(_05266_));
 sky130_fd_sc_hd__o211a_1 _12078_ (.A1(\rbzero.tex_r1[23] ),
    .A2(_05243_),
    .B1(_05266_),
    .C1(_05229_),
    .X(_05267_));
 sky130_fd_sc_hd__a31o_1 _12079_ (.A1(\rbzero.tex_r1[21] ),
    .A2(_04930_),
    .A3(_05245_),
    .B1(_04946_),
    .X(_05268_));
 sky130_fd_sc_hd__a31o_1 _12080_ (.A1(\rbzero.tex_r1[20] ),
    .A2(_05224_),
    .A3(_05243_),
    .B1(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__or2_1 _12081_ (.A(\rbzero.tex_r1[18] ),
    .B(_05245_),
    .X(_05270_));
 sky130_fd_sc_hd__o211a_1 _12082_ (.A1(\rbzero.tex_r1[19] ),
    .A2(_05243_),
    .B1(_05270_),
    .C1(_05229_),
    .X(_05271_));
 sky130_fd_sc_hd__a31o_1 _12083_ (.A1(\rbzero.tex_r1[17] ),
    .A2(_04991_),
    .A3(_05233_),
    .B1(_04932_),
    .X(_05272_));
 sky130_fd_sc_hd__a31o_1 _12084_ (.A1(\rbzero.tex_r1[16] ),
    .A2(_05224_),
    .A3(_04899_),
    .B1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__o221a_1 _12085_ (.A1(_05267_),
    .A2(_05269_),
    .B1(_05271_),
    .B2(_05273_),
    .C1(_05254_),
    .X(_05274_));
 sky130_fd_sc_hd__a311o_1 _12086_ (.A1(_05223_),
    .A2(_05260_),
    .A3(_05265_),
    .B1(_04965_),
    .C1(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__buf_4 _12087_ (.A(_04939_),
    .X(_05276_));
 sky130_fd_sc_hd__clkbuf_8 _12088_ (.A(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__or2_1 _12089_ (.A(\rbzero.tex_r1[62] ),
    .B(_05036_),
    .X(_05278_));
 sky130_fd_sc_hd__o211a_1 _12090_ (.A1(\rbzero.tex_r1[63] ),
    .A2(_05277_),
    .B1(_05278_),
    .C1(_04934_),
    .X(_05279_));
 sky130_fd_sc_hd__a31o_1 _12091_ (.A1(\rbzero.tex_r1[61] ),
    .A2(_05231_),
    .A3(_05233_),
    .B1(_04946_),
    .X(_05280_));
 sky130_fd_sc_hd__a311o_1 _12092_ (.A1(\rbzero.tex_r1[60] ),
    .A2(_05232_),
    .A3(_05243_),
    .B1(_05279_),
    .C1(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__or2_1 _12093_ (.A(\rbzero.tex_r1[58] ),
    .B(_05244_),
    .X(_05282_));
 sky130_fd_sc_hd__o211a_1 _12094_ (.A1(\rbzero.tex_r1[59] ),
    .A2(_05277_),
    .B1(_05282_),
    .C1(_04934_),
    .X(_05283_));
 sky130_fd_sc_hd__a31o_1 _12095_ (.A1(\rbzero.tex_r1[57] ),
    .A2(_05231_),
    .A3(_05245_),
    .B1(_04932_),
    .X(_05284_));
 sky130_fd_sc_hd__a311o_1 _12096_ (.A1(\rbzero.tex_r1[56] ),
    .A2(_05232_),
    .A3(_05243_),
    .B1(_05283_),
    .C1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__or2_1 _12097_ (.A(\rbzero.tex_r1[54] ),
    .B(_05036_),
    .X(_05286_));
 sky130_fd_sc_hd__buf_4 _12098_ (.A(_04956_),
    .X(_05287_));
 sky130_fd_sc_hd__o211a_1 _12099_ (.A1(\rbzero.tex_r1[55] ),
    .A2(_05242_),
    .B1(_05286_),
    .C1(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__clkbuf_4 _12100_ (.A(_04879_),
    .X(_05289_));
 sky130_fd_sc_hd__a31o_1 _12101_ (.A1(\rbzero.tex_r1[53] ),
    .A2(_05027_),
    .A3(_05289_),
    .B1(_04945_),
    .X(_05290_));
 sky130_fd_sc_hd__a31o_1 _12102_ (.A1(\rbzero.tex_r1[52] ),
    .A2(_04991_),
    .A3(_04898_),
    .B1(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__or2_1 _12103_ (.A(\rbzero.tex_r1[50] ),
    .B(_05289_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_8 _12104_ (.A(_04873_),
    .X(_05293_));
 sky130_fd_sc_hd__buf_6 _12105_ (.A(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__o211a_1 _12106_ (.A1(\rbzero.tex_r1[51] ),
    .A2(_04898_),
    .B1(_05292_),
    .C1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__a31o_1 _12107_ (.A1(\rbzero.tex_r1[49] ),
    .A2(_04942_),
    .A3(_05227_),
    .B1(_04931_),
    .X(_05296_));
 sky130_fd_sc_hd__a31o_1 _12108_ (.A1(\rbzero.tex_r1[48] ),
    .A2(_05263_),
    .A3(_04898_),
    .B1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__o221a_1 _12109_ (.A1(_05288_),
    .A2(_05291_),
    .B1(_05295_),
    .B2(_05297_),
    .C1(_05254_),
    .X(_05298_));
 sky130_fd_sc_hd__a311o_1 _12110_ (.A1(_05223_),
    .A2(_05281_),
    .A3(_05285_),
    .B1(_04965_),
    .C1(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__or2_1 _12111_ (.A(\rbzero.tex_r1[46] ),
    .B(_05244_),
    .X(_05300_));
 sky130_fd_sc_hd__o211a_1 _12112_ (.A1(\rbzero.tex_r1[47] ),
    .A2(_05277_),
    .B1(_05300_),
    .C1(_04934_),
    .X(_05301_));
 sky130_fd_sc_hd__a31o_1 _12113_ (.A1(\rbzero.tex_r1[45] ),
    .A2(_05231_),
    .A3(_05245_),
    .B1(_04946_),
    .X(_05302_));
 sky130_fd_sc_hd__a311o_1 _12114_ (.A1(\rbzero.tex_r1[44] ),
    .A2(_05232_),
    .A3(_05243_),
    .B1(_05301_),
    .C1(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__buf_4 _12115_ (.A(_04925_),
    .X(_05304_));
 sky130_fd_sc_hd__or2_1 _12116_ (.A(\rbzero.tex_r1[42] ),
    .B(_05244_),
    .X(_05305_));
 sky130_fd_sc_hd__o211a_1 _12117_ (.A1(\rbzero.tex_r1[43] ),
    .A2(_05304_),
    .B1(_05305_),
    .C1(_04934_),
    .X(_05306_));
 sky130_fd_sc_hd__a31o_1 _12118_ (.A1(\rbzero.tex_r1[41] ),
    .A2(_05231_),
    .A3(_05245_),
    .B1(_04960_),
    .X(_05307_));
 sky130_fd_sc_hd__a311o_1 _12119_ (.A1(\rbzero.tex_r1[40] ),
    .A2(_05232_),
    .A3(_05226_),
    .B1(_05306_),
    .C1(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__or2_1 _12120_ (.A(\rbzero.tex_r1[38] ),
    .B(_05036_),
    .X(_05309_));
 sky130_fd_sc_hd__o211a_1 _12121_ (.A1(\rbzero.tex_r1[39] ),
    .A2(_05242_),
    .B1(_05309_),
    .C1(_05287_),
    .X(_05310_));
 sky130_fd_sc_hd__a31o_1 _12122_ (.A1(\rbzero.tex_r1[37] ),
    .A2(_05027_),
    .A3(_05289_),
    .B1(_04945_),
    .X(_05311_));
 sky130_fd_sc_hd__a31o_1 _12123_ (.A1(\rbzero.tex_r1[36] ),
    .A2(_04991_),
    .A3(_04898_),
    .B1(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__or2_1 _12124_ (.A(\rbzero.tex_r1[34] ),
    .B(_05036_),
    .X(_05313_));
 sky130_fd_sc_hd__o211a_1 _12125_ (.A1(\rbzero.tex_r1[35] ),
    .A2(_04898_),
    .B1(_05313_),
    .C1(_05287_),
    .X(_05314_));
 sky130_fd_sc_hd__a31o_1 _12126_ (.A1(\rbzero.tex_r1[33] ),
    .A2(_04942_),
    .A3(_05227_),
    .B1(_04931_),
    .X(_05315_));
 sky130_fd_sc_hd__a31o_1 _12127_ (.A1(\rbzero.tex_r1[32] ),
    .A2(_05263_),
    .A3(_04898_),
    .B1(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__o221a_1 _12128_ (.A1(_05310_),
    .A2(_05312_),
    .B1(_05314_),
    .B2(_05316_),
    .C1(_05254_),
    .X(_05317_));
 sky130_fd_sc_hd__a311o_1 _12129_ (.A1(_05223_),
    .A2(_05303_),
    .A3(_05308_),
    .B1(_05241_),
    .C1(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__buf_4 _12130_ (.A(net42),
    .X(_05319_));
 sky130_fd_sc_hd__a31o_1 _12131_ (.A1(_05023_),
    .A2(_05299_),
    .A3(_05318_),
    .B1(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__a31oi_4 _12132_ (.A1(_04985_),
    .A2(_05256_),
    .A3(_05275_),
    .B1(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__nand2_1 _12133_ (.A(\rbzero.row_render.side ),
    .B(_04890_),
    .Y(_05322_));
 sky130_fd_sc_hd__and2_1 _12134_ (.A(_04902_),
    .B(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__o21ai_1 _12135_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_05241_),
    .B1(_04905_),
    .Y(_05324_));
 sky130_fd_sc_hd__a21o_1 _12136_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_05241_),
    .B1(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__o211a_1 _12137_ (.A1(_04914_),
    .A2(_05323_),
    .B1(_05325_),
    .C1(_05319_),
    .X(_05326_));
 sky130_fd_sc_hd__or3b_1 _12138_ (.A(_05321_),
    .B(_05326_),
    .C_N(_05090_),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(\rbzero.color_sky[1] ),
    .A1(\rbzero.color_floor[1] ),
    .S(_04808_),
    .X(_05328_));
 sky130_fd_sc_hd__o21ai_1 _12140_ (.A1(_05033_),
    .A2(_05089_),
    .B1(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__nor2_1 _12141_ (.A(_04743_),
    .B(_04766_),
    .Y(_05330_));
 sky130_fd_sc_hd__a2bb2o_1 _12142_ (.A1_N(\gpout0.vpos[4] ),
    .A2_N(_04642_),
    .B1(_04471_),
    .B2(\gpout0.vpos[3] ),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_1 _12143_ (.A1(_04701_),
    .A2(_04642_),
    .B1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__nand2_1 _12144_ (.A(_04699_),
    .B(_04474_),
    .Y(_05333_));
 sky130_fd_sc_hd__or2_1 _12145_ (.A(_04699_),
    .B(_04473_),
    .X(_05334_));
 sky130_fd_sc_hd__o2111a_1 _12146_ (.A1(\gpout0.vpos[3] ),
    .A2(_04471_),
    .B1(_04514_),
    .C1(_05333_),
    .D1(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__o2bb2a_1 _12147_ (.A1_N(_05332_),
    .A2_N(_05335_),
    .B1(_04714_),
    .B2(_04717_),
    .X(_05336_));
 sky130_fd_sc_hd__and4_1 _12148_ (.A(_04031_),
    .B(_04480_),
    .C(_04474_),
    .D(_04478_),
    .X(_05337_));
 sky130_fd_sc_hd__a211oi_1 _12149_ (.A1(_05333_),
    .A2(_05334_),
    .B1(_04723_),
    .C1(_04471_),
    .Y(_05338_));
 sky130_fd_sc_hd__a311oi_1 _12150_ (.A1(_04701_),
    .A2(_04723_),
    .A3(_05099_),
    .B1(_05337_),
    .C1(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__a211o_1 _12151_ (.A1(_04702_),
    .A2(_04703_),
    .B1(_05333_),
    .C1(_04477_),
    .X(_05340_));
 sky130_fd_sc_hd__o211a_1 _12152_ (.A1(_04718_),
    .A2(_05336_),
    .B1(_05339_),
    .C1(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__o21ai_1 _12153_ (.A1(_04474_),
    .A2(_04762_),
    .B1(_05341_),
    .Y(_05342_));
 sky130_fd_sc_hd__and2_1 _12154_ (.A(_05330_),
    .B(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__or3b_1 _12155_ (.A(_04770_),
    .B(_04031_),
    .C_N(_04644_),
    .X(_05344_));
 sky130_fd_sc_hd__nand2_1 _12156_ (.A(_04701_),
    .B(_04480_),
    .Y(_05345_));
 sky130_fd_sc_hd__or4_1 _12157_ (.A(_04714_),
    .B(_04723_),
    .C(_05334_),
    .D(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__xnor2_1 _12158_ (.A(_04723_),
    .B(_04642_),
    .Y(_05347_));
 sky130_fd_sc_hd__nor2_1 _12159_ (.A(_04699_),
    .B(_04513_),
    .Y(_05348_));
 sky130_fd_sc_hd__nor2_1 _12160_ (.A(_04729_),
    .B(_04476_),
    .Y(_05349_));
 sky130_fd_sc_hd__or2_1 _12161_ (.A(\gpout0.vpos[4] ),
    .B(_04480_),
    .X(_05350_));
 sky130_fd_sc_hd__nand2_1 _12162_ (.A(_04718_),
    .B(_04474_),
    .Y(_05351_));
 sky130_fd_sc_hd__or2_1 _12163_ (.A(_04718_),
    .B(_04474_),
    .X(_05352_));
 sky130_fd_sc_hd__and4_1 _12164_ (.A(_05345_),
    .B(_05350_),
    .C(_05351_),
    .D(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__or4b_1 _12165_ (.A(_05347_),
    .B(_05348_),
    .C(_05349_),
    .D_N(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__o21ai_2 _12166_ (.A1(_05344_),
    .A2(_05346_),
    .B1(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__inv_2 _12167_ (.A(_04805_),
    .Y(_05356_));
 sky130_fd_sc_hd__nor2_1 _12168_ (.A(_05356_),
    .B(_04788_),
    .Y(_05357_));
 sky130_fd_sc_hd__nor2_1 _12169_ (.A(_04767_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__a311oi_2 _12170_ (.A1(_04779_),
    .A2(_05343_),
    .A3(_05355_),
    .B1(_05358_),
    .C1(_04765_),
    .Y(_05359_));
 sky130_fd_sc_hd__a31oi_1 _12171_ (.A1(_04764_),
    .A2(_05327_),
    .A3(_05329_),
    .B1(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__nor2_1 _12172_ (.A(_04720_),
    .B(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__o21ai_1 _12173_ (.A1(_05222_),
    .A2(_05361_),
    .B1(_05096_),
    .Y(_05362_));
 sky130_fd_sc_hd__o211ai_4 _12174_ (.A1(_04493_),
    .A2(_04695_),
    .B1(_05101_),
    .C1(_05362_),
    .Y(_05363_));
 sky130_fd_sc_hd__clkinv_2 _12175_ (.A(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__mux2_2 _12176_ (.A0(\reg_rgb[7] ),
    .A1(_05364_),
    .S(_05103_),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_1 _12177_ (.A(_05365_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _12178_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04920_),
    .X(_05366_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04920_),
    .X(_05367_));
 sky130_fd_sc_hd__mux2_1 _12180_ (.A0(_05366_),
    .A1(_05367_),
    .S(_04930_),
    .X(_05368_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_04920_),
    .X(_05369_));
 sky130_fd_sc_hd__mux2_1 _12182_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_04920_),
    .X(_05370_));
 sky130_fd_sc_hd__buf_4 _12183_ (.A(_04910_),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _12184_ (.A0(_05369_),
    .A1(_05370_),
    .S(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__buf_6 _12185_ (.A(_04946_),
    .X(_05373_));
 sky130_fd_sc_hd__mux2_1 _12186_ (.A0(_05368_),
    .A1(_05372_),
    .S(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__mux2_1 _12187_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_05277_),
    .X(_05375_));
 sky130_fd_sc_hd__and3_1 _12188_ (.A(\rbzero.tex_g0[11] ),
    .B(_04936_),
    .C(_04937_),
    .X(_05376_));
 sky130_fd_sc_hd__a21o_1 _12189_ (.A1(\rbzero.tex_g0[10] ),
    .A2(_05226_),
    .B1(_05263_),
    .X(_05377_));
 sky130_fd_sc_hd__o221a_1 _12190_ (.A1(_05229_),
    .A2(_05375_),
    .B1(_05376_),
    .B2(_05377_),
    .C1(_05373_),
    .X(_05378_));
 sky130_fd_sc_hd__mux2_1 _12191_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04940_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _12192_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_04940_),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _12193_ (.A0(_05379_),
    .A1(_05380_),
    .S(_05294_),
    .X(_05381_));
 sky130_fd_sc_hd__a21o_1 _12194_ (.A1(_05238_),
    .A2(_05381_),
    .B1(_05254_),
    .X(_05382_));
 sky130_fd_sc_hd__o221a_1 _12195_ (.A1(_05223_),
    .A2(_05374_),
    .B1(_05378_),
    .B2(_05382_),
    .C1(_04965_),
    .X(_05383_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_05276_),
    .X(_05384_));
 sky130_fd_sc_hd__mux2_1 _12197_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_05276_),
    .X(_05385_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(_05384_),
    .A1(_05385_),
    .S(_05263_),
    .X(_05386_));
 sky130_fd_sc_hd__mux2_1 _12199_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_05276_),
    .X(_05387_));
 sky130_fd_sc_hd__and3_1 _12200_ (.A(\rbzero.tex_g0[27] ),
    .B(_04936_),
    .C(_04937_),
    .X(_05388_));
 sky130_fd_sc_hd__buf_4 _12201_ (.A(_04929_),
    .X(_05389_));
 sky130_fd_sc_hd__a21o_1 _12202_ (.A1(\rbzero.tex_g0[26] ),
    .A2(_05304_),
    .B1(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__o221a_1 _12203_ (.A1(_05294_),
    .A2(_05387_),
    .B1(_05388_),
    .B2(_05390_),
    .C1(_04952_),
    .X(_05391_));
 sky130_fd_sc_hd__a211o_1 _12204_ (.A1(_05238_),
    .A2(_05386_),
    .B1(_05391_),
    .C1(_05254_),
    .X(_05392_));
 sky130_fd_sc_hd__mux2_1 _12205_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_05276_),
    .X(_05393_));
 sky130_fd_sc_hd__mux2_1 _12206_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_05276_),
    .X(_05394_));
 sky130_fd_sc_hd__mux2_1 _12207_ (.A0(_05393_),
    .A1(_05394_),
    .S(_05287_),
    .X(_05395_));
 sky130_fd_sc_hd__and2_1 _12208_ (.A(\rbzero.tex_g0[20] ),
    .B(_05225_),
    .X(_05396_));
 sky130_fd_sc_hd__a31o_1 _12209_ (.A1(\rbzero.tex_g0[21] ),
    .A2(_04936_),
    .A3(_04937_),
    .B1(_05293_),
    .X(_05397_));
 sky130_fd_sc_hd__mux2_1 _12210_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_05276_),
    .X(_05398_));
 sky130_fd_sc_hd__o221a_1 _12211_ (.A1(_05396_),
    .A2(_05397_),
    .B1(_05398_),
    .B2(_05263_),
    .C1(_04932_),
    .X(_05399_));
 sky130_fd_sc_hd__a211o_1 _12212_ (.A1(_05373_),
    .A2(_05395_),
    .B1(_05399_),
    .C1(_04918_),
    .X(_05400_));
 sky130_fd_sc_hd__a31o_1 _12213_ (.A1(_05241_),
    .A2(_05392_),
    .A3(_05400_),
    .B1(_05023_),
    .X(_05401_));
 sky130_fd_sc_hd__and2_1 _12214_ (.A(\rbzero.tex_g0[52] ),
    .B(_05226_),
    .X(_05402_));
 sky130_fd_sc_hd__a31o_1 _12215_ (.A1(\rbzero.tex_g0[53] ),
    .A2(_04936_),
    .A3(_04937_),
    .B1(_05294_),
    .X(_05403_));
 sky130_fd_sc_hd__mux2_1 _12216_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_05277_),
    .X(_05404_));
 sky130_fd_sc_hd__o221a_1 _12217_ (.A1(_05402_),
    .A2(_05403_),
    .B1(_05404_),
    .B2(_05224_),
    .C1(_05238_),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_1 _12218_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_05277_),
    .X(_05406_));
 sky130_fd_sc_hd__and3_1 _12219_ (.A(\rbzero.tex_g0[51] ),
    .B(_04936_),
    .C(_04937_),
    .X(_05407_));
 sky130_fd_sc_hd__a21o_1 _12220_ (.A1(\rbzero.tex_g0[50] ),
    .A2(_05226_),
    .B1(_05263_),
    .X(_05408_));
 sky130_fd_sc_hd__o221a_1 _12221_ (.A1(_05229_),
    .A2(_05406_),
    .B1(_05407_),
    .B2(_05408_),
    .C1(_05373_),
    .X(_05409_));
 sky130_fd_sc_hd__mux2_1 _12222_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_04897_),
    .X(_05410_));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04897_),
    .X(_05411_));
 sky130_fd_sc_hd__mux2_1 _12224_ (.A0(_05410_),
    .A1(_05411_),
    .S(_05294_),
    .X(_05412_));
 sky130_fd_sc_hd__mux2_1 _12225_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_05225_),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_04896_),
    .X(_05414_));
 sky130_fd_sc_hd__or2_1 _12227_ (.A(_04930_),
    .B(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__o211a_1 _12228_ (.A1(_05294_),
    .A2(_05413_),
    .B1(_05415_),
    .C1(_05238_),
    .X(_05416_));
 sky130_fd_sc_hd__a211o_1 _12229_ (.A1(_05373_),
    .A2(_05412_),
    .B1(_05416_),
    .C1(_05254_),
    .X(_05417_));
 sky130_fd_sc_hd__o311a_1 _12230_ (.A1(_05223_),
    .A2(_05405_),
    .A3(_05409_),
    .B1(_05241_),
    .C1(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__mux2_1 _12231_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04940_),
    .X(_05419_));
 sky130_fd_sc_hd__mux2_1 _12232_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04940_),
    .X(_05420_));
 sky130_fd_sc_hd__mux2_1 _12233_ (.A0(_05419_),
    .A1(_05420_),
    .S(_05287_),
    .X(_05421_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04897_),
    .X(_05422_));
 sky130_fd_sc_hd__mux2_1 _12235_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04939_),
    .X(_05423_));
 sky130_fd_sc_hd__or2_1 _12236_ (.A(_05389_),
    .B(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__o211a_1 _12237_ (.A1(_05294_),
    .A2(_05422_),
    .B1(_05424_),
    .C1(_05238_),
    .X(_05425_));
 sky130_fd_sc_hd__a211o_1 _12238_ (.A1(_05373_),
    .A2(_05421_),
    .B1(_05425_),
    .C1(_05223_),
    .X(_05426_));
 sky130_fd_sc_hd__mux2_1 _12239_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04940_),
    .X(_05427_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_05276_),
    .X(_05428_));
 sky130_fd_sc_hd__mux2_1 _12241_ (.A0(_05427_),
    .A1(_05428_),
    .S(_05287_),
    .X(_05429_));
 sky130_fd_sc_hd__buf_4 _12242_ (.A(_04924_),
    .X(_05430_));
 sky130_fd_sc_hd__buf_4 _12243_ (.A(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__and2_1 _12244_ (.A(\rbzero.tex_g0[44] ),
    .B(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__a31o_1 _12245_ (.A1(\rbzero.tex_g0[45] ),
    .A2(_04936_),
    .A3(_04937_),
    .B1(_05293_),
    .X(_05433_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04940_),
    .X(_05434_));
 sky130_fd_sc_hd__o221a_1 _12247_ (.A1(_05432_),
    .A2(_05433_),
    .B1(_05434_),
    .B2(_05263_),
    .C1(_05238_),
    .X(_05435_));
 sky130_fd_sc_hd__a211o_1 _12248_ (.A1(_05373_),
    .A2(_05429_),
    .B1(_05435_),
    .C1(_05254_),
    .X(_05436_));
 sky130_fd_sc_hd__a31o_1 _12249_ (.A1(_04965_),
    .A2(_05426_),
    .A3(_05436_),
    .B1(_04985_),
    .X(_05437_));
 sky130_fd_sc_hd__o221a_2 _12250_ (.A1(_05383_),
    .A2(_05401_),
    .B1(_05418_),
    .B2(_05437_),
    .C1(_04906_),
    .X(_05438_));
 sky130_fd_sc_hd__and3_1 _12251_ (.A(_05294_),
    .B(_04932_),
    .C(_05233_),
    .X(_05439_));
 sky130_fd_sc_hd__a31oi_1 _12252_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04876_),
    .A3(_04899_),
    .B1(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__o21ai_1 _12253_ (.A1(_04889_),
    .A2(_05440_),
    .B1(\rbzero.row_render.side ),
    .Y(_05441_));
 sky130_fd_sc_hd__a31o_1 _12254_ (.A1(\rbzero.row_render.side ),
    .A2(\rbzero.row_render.wall[0] ),
    .A3(_04912_),
    .B1(_04905_),
    .X(_05442_));
 sky130_fd_sc_hd__a31o_1 _12255_ (.A1(_04891_),
    .A2(_04902_),
    .A3(_05441_),
    .B1(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__a211o_1 _12256_ (.A1(_04907_),
    .A2(_05443_),
    .B1(_05033_),
    .C1(_05089_),
    .X(_05444_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_04808_),
    .X(_05445_));
 sky130_fd_sc_hd__o221ai_4 _12258_ (.A1(_05438_),
    .A2(_05444_),
    .B1(_05445_),
    .B2(_05090_),
    .C1(_04764_),
    .Y(_05446_));
 sky130_fd_sc_hd__nand2_1 _12259_ (.A(_05092_),
    .B(_04743_),
    .Y(_05447_));
 sky130_fd_sc_hd__and3b_1 _12260_ (.A_N(_04720_),
    .B(_05446_),
    .C(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__o21ai_1 _12261_ (.A1(_04721_),
    .A2(_05448_),
    .B1(_05096_),
    .Y(_05449_));
 sky130_fd_sc_hd__o211a_2 _12262_ (.A1(_04486_),
    .A2(_04695_),
    .B1(_05101_),
    .C1(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__mux2_2 _12263_ (.A0(\reg_rgb[14] ),
    .A1(_05450_),
    .S(_05103_),
    .X(_05451_));
 sky130_fd_sc_hd__clkbuf_1 _12264_ (.A(_05451_),
    .X(net65));
 sky130_fd_sc_hd__or2_1 _12265_ (.A(\rbzero.tex_g1[14] ),
    .B(_05036_),
    .X(_05452_));
 sky130_fd_sc_hd__o211a_1 _12266_ (.A1(\rbzero.tex_g1[15] ),
    .A2(_05277_),
    .B1(_05452_),
    .C1(_05287_),
    .X(_05453_));
 sky130_fd_sc_hd__a31o_1 _12267_ (.A1(\rbzero.tex_g1[13] ),
    .A2(_05231_),
    .A3(_05233_),
    .B1(_04946_),
    .X(_05454_));
 sky130_fd_sc_hd__a311o_1 _12268_ (.A1(\rbzero.tex_g1[12] ),
    .A2(_05224_),
    .A3(_05243_),
    .B1(_05453_),
    .C1(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__or2_1 _12269_ (.A(\rbzero.tex_g1[10] ),
    .B(_05036_),
    .X(_05456_));
 sky130_fd_sc_hd__o211a_1 _12270_ (.A1(\rbzero.tex_g1[11] ),
    .A2(_05277_),
    .B1(_05456_),
    .C1(_04934_),
    .X(_05457_));
 sky130_fd_sc_hd__a31o_1 _12271_ (.A1(\rbzero.tex_g1[9] ),
    .A2(_05231_),
    .A3(_05233_),
    .B1(_04932_),
    .X(_05458_));
 sky130_fd_sc_hd__a311o_1 _12272_ (.A1(\rbzero.tex_g1[8] ),
    .A2(_05232_),
    .A3(_05243_),
    .B1(_05457_),
    .C1(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__or2_1 _12273_ (.A(\rbzero.tex_g1[6] ),
    .B(_05036_),
    .X(_05460_));
 sky130_fd_sc_hd__o211a_1 _12274_ (.A1(\rbzero.tex_g1[7] ),
    .A2(_05242_),
    .B1(_05460_),
    .C1(_05287_),
    .X(_05461_));
 sky130_fd_sc_hd__a31o_1 _12275_ (.A1(\rbzero.tex_g1[5] ),
    .A2(_05027_),
    .A3(_05289_),
    .B1(_04945_),
    .X(_05462_));
 sky130_fd_sc_hd__a31o_1 _12276_ (.A1(\rbzero.tex_g1[4] ),
    .A2(_04991_),
    .A3(_04898_),
    .B1(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__or2_1 _12277_ (.A(\rbzero.tex_g1[2] ),
    .B(_05289_),
    .X(_05464_));
 sky130_fd_sc_hd__o211a_1 _12278_ (.A1(\rbzero.tex_g1[3] ),
    .A2(_04898_),
    .B1(_05464_),
    .C1(_05294_),
    .X(_05465_));
 sky130_fd_sc_hd__a31o_1 _12279_ (.A1(\rbzero.tex_g1[1] ),
    .A2(_04942_),
    .A3(_05227_),
    .B1(_04931_),
    .X(_05466_));
 sky130_fd_sc_hd__a31o_1 _12280_ (.A1(\rbzero.tex_g1[0] ),
    .A2(_05263_),
    .A3(_05226_),
    .B1(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__o221a_1 _12281_ (.A1(_05461_),
    .A2(_05463_),
    .B1(_05465_),
    .B2(_05467_),
    .C1(_05254_),
    .X(_05468_));
 sky130_fd_sc_hd__a311o_1 _12282_ (.A1(_05223_),
    .A2(_05455_),
    .A3(_05459_),
    .B1(_05241_),
    .C1(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__or2_1 _12283_ (.A(\rbzero.tex_g1[30] ),
    .B(_05244_),
    .X(_05470_));
 sky130_fd_sc_hd__o211a_1 _12284_ (.A1(\rbzero.tex_g1[31] ),
    .A2(_05277_),
    .B1(_05470_),
    .C1(_04934_),
    .X(_05471_));
 sky130_fd_sc_hd__a31o_1 _12285_ (.A1(\rbzero.tex_g1[29] ),
    .A2(_05231_),
    .A3(_05245_),
    .B1(_04946_),
    .X(_05472_));
 sky130_fd_sc_hd__a311o_1 _12286_ (.A1(\rbzero.tex_g1[28] ),
    .A2(_05232_),
    .A3(_05243_),
    .B1(_05471_),
    .C1(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__or2_1 _12287_ (.A(\rbzero.tex_g1[26] ),
    .B(_05244_),
    .X(_05474_));
 sky130_fd_sc_hd__o211a_1 _12288_ (.A1(\rbzero.tex_g1[27] ),
    .A2(_05304_),
    .B1(_05474_),
    .C1(_04934_),
    .X(_05475_));
 sky130_fd_sc_hd__a31o_1 _12289_ (.A1(\rbzero.tex_g1[25] ),
    .A2(_04930_),
    .A3(_05245_),
    .B1(_04960_),
    .X(_05476_));
 sky130_fd_sc_hd__a311o_1 _12290_ (.A1(\rbzero.tex_g1[24] ),
    .A2(_05232_),
    .A3(_05226_),
    .B1(_05475_),
    .C1(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__or2_1 _12291_ (.A(\rbzero.tex_g1[22] ),
    .B(_05036_),
    .X(_05478_));
 sky130_fd_sc_hd__o211a_1 _12292_ (.A1(\rbzero.tex_g1[23] ),
    .A2(_05242_),
    .B1(_05478_),
    .C1(_05287_),
    .X(_05479_));
 sky130_fd_sc_hd__a31o_1 _12293_ (.A1(\rbzero.tex_g1[21] ),
    .A2(_05027_),
    .A3(_05289_),
    .B1(_05028_),
    .X(_05480_));
 sky130_fd_sc_hd__a31o_1 _12294_ (.A1(\rbzero.tex_g1[20] ),
    .A2(_04991_),
    .A3(_05242_),
    .B1(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__or2_1 _12295_ (.A(\rbzero.tex_g1[18] ),
    .B(_05036_),
    .X(_05482_));
 sky130_fd_sc_hd__o211a_1 _12296_ (.A1(\rbzero.tex_g1[19] ),
    .A2(_05242_),
    .B1(_05482_),
    .C1(_05287_),
    .X(_05483_));
 sky130_fd_sc_hd__a31o_1 _12297_ (.A1(\rbzero.tex_g1[17] ),
    .A2(_04942_),
    .A3(_05227_),
    .B1(_04931_),
    .X(_05484_));
 sky130_fd_sc_hd__a31o_1 _12298_ (.A1(\rbzero.tex_g1[16] ),
    .A2(_05263_),
    .A3(_04898_),
    .B1(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__o221a_1 _12299_ (.A1(_05479_),
    .A2(_05481_),
    .B1(_05483_),
    .B2(_05485_),
    .C1(_05254_),
    .X(_05486_));
 sky130_fd_sc_hd__a311o_1 _12300_ (.A1(_05223_),
    .A2(_05473_),
    .A3(_05477_),
    .B1(_04965_),
    .C1(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__or2_1 _12301_ (.A(\rbzero.tex_g1[46] ),
    .B(_04879_),
    .X(_05488_));
 sky130_fd_sc_hd__o211a_1 _12302_ (.A1(\rbzero.tex_g1[47] ),
    .A2(_05276_),
    .B1(_05488_),
    .C1(_04956_),
    .X(_05489_));
 sky130_fd_sc_hd__a31o_1 _12303_ (.A1(\rbzero.tex_g1[45] ),
    .A2(_04942_),
    .A3(_05289_),
    .B1(_04945_),
    .X(_05490_));
 sky130_fd_sc_hd__a311o_1 _12304_ (.A1(\rbzero.tex_g1[44] ),
    .A2(_04991_),
    .A3(_05242_),
    .B1(_05489_),
    .C1(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__or2_1 _12305_ (.A(\rbzero.tex_g1[42] ),
    .B(_04879_),
    .X(_05492_));
 sky130_fd_sc_hd__o211a_1 _12306_ (.A1(\rbzero.tex_g1[43] ),
    .A2(_04920_),
    .B1(_05492_),
    .C1(_04922_),
    .X(_05493_));
 sky130_fd_sc_hd__a31o_1 _12307_ (.A1(\rbzero.tex_g1[41] ),
    .A2(_05027_),
    .A3(_05289_),
    .B1(_04931_),
    .X(_05494_));
 sky130_fd_sc_hd__a311o_1 _12308_ (.A1(\rbzero.tex_g1[40] ),
    .A2(_05231_),
    .A3(_05242_),
    .B1(_05493_),
    .C1(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__or2_1 _12309_ (.A(\rbzero.tex_g1[38] ),
    .B(_04879_),
    .X(_05496_));
 sky130_fd_sc_hd__o211a_1 _12310_ (.A1(\rbzero.tex_g1[39] ),
    .A2(_04897_),
    .B1(_05496_),
    .C1(_04956_),
    .X(_05497_));
 sky130_fd_sc_hd__clkbuf_4 _12311_ (.A(_04878_),
    .X(_05498_));
 sky130_fd_sc_hd__a31o_1 _12312_ (.A1(\rbzero.tex_g1[37] ),
    .A2(_04928_),
    .A3(_05498_),
    .B1(_05028_),
    .X(_05499_));
 sky130_fd_sc_hd__a31o_1 _12313_ (.A1(\rbzero.tex_g1[36] ),
    .A2(_04942_),
    .A3(_04897_),
    .B1(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__or2_1 _12314_ (.A(\rbzero.tex_g1[34] ),
    .B(_04879_),
    .X(_05501_));
 sky130_fd_sc_hd__o211a_1 _12315_ (.A1(\rbzero.tex_g1[35] ),
    .A2(_04897_),
    .B1(_05501_),
    .C1(_05293_),
    .X(_05502_));
 sky130_fd_sc_hd__a31o_1 _12316_ (.A1(\rbzero.tex_g1[33] ),
    .A2(_04941_),
    .A3(_05498_),
    .B1(_04911_),
    .X(_05503_));
 sky130_fd_sc_hd__a31o_1 _12317_ (.A1(\rbzero.tex_g1[32] ),
    .A2(_04995_),
    .A3(_05225_),
    .B1(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__o221a_1 _12318_ (.A1(_05497_),
    .A2(_05500_),
    .B1(_05502_),
    .B2(_05504_),
    .C1(_04908_),
    .X(_05505_));
 sky130_fd_sc_hd__a311o_1 _12319_ (.A1(_04918_),
    .A2(_05491_),
    .A3(_05495_),
    .B1(_04951_),
    .C1(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__or2_1 _12320_ (.A(\rbzero.tex_g1[54] ),
    .B(_04879_),
    .X(_05507_));
 sky130_fd_sc_hd__o211a_1 _12321_ (.A1(\rbzero.tex_g1[55] ),
    .A2(_05276_),
    .B1(_05507_),
    .C1(_04956_),
    .X(_05508_));
 sky130_fd_sc_hd__a31o_1 _12322_ (.A1(\rbzero.tex_g1[53] ),
    .A2(_05027_),
    .A3(_05289_),
    .B1(_04945_),
    .X(_05509_));
 sky130_fd_sc_hd__a311o_1 _12323_ (.A1(\rbzero.tex_g1[52] ),
    .A2(_04991_),
    .A3(_05242_),
    .B1(_05508_),
    .C1(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__or2_1 _12324_ (.A(\rbzero.tex_g1[50] ),
    .B(_05035_),
    .X(_05511_));
 sky130_fd_sc_hd__o211a_1 _12325_ (.A1(\rbzero.tex_g1[51] ),
    .A2(_04920_),
    .B1(_05511_),
    .C1(_04922_),
    .X(_05512_));
 sky130_fd_sc_hd__a31o_1 _12326_ (.A1(\rbzero.tex_g1[49] ),
    .A2(_05027_),
    .A3(_05289_),
    .B1(_04931_),
    .X(_05513_));
 sky130_fd_sc_hd__a311o_1 _12327_ (.A1(\rbzero.tex_g1[48] ),
    .A2(_05231_),
    .A3(_05277_),
    .B1(_05512_),
    .C1(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__or2_1 _12328_ (.A(\rbzero.tex_g1[62] ),
    .B(_04879_),
    .X(_05515_));
 sky130_fd_sc_hd__o211a_1 _12329_ (.A1(\rbzero.tex_g1[63] ),
    .A2(_04940_),
    .B1(_05515_),
    .C1(_04956_),
    .X(_05516_));
 sky130_fd_sc_hd__a31o_1 _12330_ (.A1(\rbzero.tex_g1[61] ),
    .A2(_04928_),
    .A3(_05498_),
    .B1(_05028_),
    .X(_05517_));
 sky130_fd_sc_hd__a31o_1 _12331_ (.A1(\rbzero.tex_g1[60] ),
    .A2(_04942_),
    .A3(_04897_),
    .B1(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__or2_1 _12332_ (.A(\rbzero.tex_g1[58] ),
    .B(_04879_),
    .X(_05519_));
 sky130_fd_sc_hd__o211a_1 _12333_ (.A1(\rbzero.tex_g1[59] ),
    .A2(_04897_),
    .B1(_05519_),
    .C1(_04956_),
    .X(_05520_));
 sky130_fd_sc_hd__a31o_1 _12334_ (.A1(\rbzero.tex_g1[57] ),
    .A2(_04941_),
    .A3(_05498_),
    .B1(_04911_),
    .X(_05521_));
 sky130_fd_sc_hd__a31o_1 _12335_ (.A1(\rbzero.tex_g1[56] ),
    .A2(_04995_),
    .A3(_04897_),
    .B1(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__o221a_1 _12336_ (.A1(_05516_),
    .A2(_05518_),
    .B1(_05520_),
    .B2(_05522_),
    .C1(_04884_),
    .X(_05523_));
 sky130_fd_sc_hd__a311o_1 _12337_ (.A1(_04987_),
    .A2(_05510_),
    .A3(_05514_),
    .B1(_04964_),
    .C1(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__a31o_1 _12338_ (.A1(_05023_),
    .A2(_05506_),
    .A3(_05524_),
    .B1(net42),
    .X(_05525_));
 sky130_fd_sc_hd__a31oi_4 _12339_ (.A1(_04985_),
    .A2(_05469_),
    .A3(_05487_),
    .B1(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__xnor2_1 _12340_ (.A(\rbzero.row_render.texu[2] ),
    .B(_05373_),
    .Y(_05527_));
 sky130_fd_sc_hd__nor2_1 _12341_ (.A(_04903_),
    .B(_05322_),
    .Y(_05528_));
 sky130_fd_sc_hd__a211oi_1 _12342_ (.A1(_04905_),
    .A2(_05527_),
    .B1(_05528_),
    .C1(_04906_),
    .Y(_05529_));
 sky130_fd_sc_hd__or3b_1 _12343_ (.A(_05526_),
    .B(_05529_),
    .C_N(_05090_),
    .X(_05530_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_04808_),
    .X(_05531_));
 sky130_fd_sc_hd__o21ai_1 _12345_ (.A1(_05033_),
    .A2(_05089_),
    .B1(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__inv_2 _12346_ (.A(_05355_),
    .Y(_05533_));
 sky130_fd_sc_hd__and2_1 _12347_ (.A(_04779_),
    .B(_05357_),
    .X(_05534_));
 sky130_fd_sc_hd__a31oi_1 _12348_ (.A1(_05343_),
    .A2(_05533_),
    .A3(_05534_),
    .B1(_04765_),
    .Y(_05535_));
 sky130_fd_sc_hd__a31oi_1 _12349_ (.A1(_04764_),
    .A2(_05530_),
    .A3(_05532_),
    .B1(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__nor2_1 _12350_ (.A(_04720_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_1 _12351_ (.A1(_05222_),
    .A2(_05537_),
    .B1(_05096_),
    .Y(_05538_));
 sky130_fd_sc_hd__o211a_2 _12352_ (.A1(\rbzero.trace_state[3] ),
    .A2(_04695_),
    .B1(_05101_),
    .C1(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__mux2_2 _12353_ (.A0(\reg_rgb[15] ),
    .A1(_05539_),
    .S(_05103_),
    .X(_05540_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_05540_),
    .X(net66));
 sky130_fd_sc_hd__o21a_1 _12355_ (.A1(_04891_),
    .A2(_05439_),
    .B1(_05323_),
    .X(_05541_));
 sky130_fd_sc_hd__a211o_1 _12356_ (.A1(\rbzero.row_render.wall[0] ),
    .A2(_04913_),
    .B1(_05442_),
    .C1(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__or2_1 _12357_ (.A(\rbzero.tex_b0[26] ),
    .B(_05498_),
    .X(_05543_));
 sky130_fd_sc_hd__o211a_1 _12358_ (.A1(\rbzero.tex_b0[27] ),
    .A2(_05225_),
    .B1(_05543_),
    .C1(_05293_),
    .X(_05544_));
 sky130_fd_sc_hd__a31o_1 _12359_ (.A1(\rbzero.tex_b0[25] ),
    .A2(_04941_),
    .A3(_05498_),
    .B1(_04911_),
    .X(_05545_));
 sky130_fd_sc_hd__a31o_1 _12360_ (.A1(\rbzero.tex_b0[24] ),
    .A2(_04995_),
    .A3(_05225_),
    .B1(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__or2_1 _12361_ (.A(\rbzero.tex_b0[30] ),
    .B(_05498_),
    .X(_05547_));
 sky130_fd_sc_hd__o211a_1 _12362_ (.A1(\rbzero.tex_b0[31] ),
    .A2(_05225_),
    .B1(_05547_),
    .C1(_05293_),
    .X(_05548_));
 sky130_fd_sc_hd__clkbuf_4 _12363_ (.A(_04878_),
    .X(_05549_));
 sky130_fd_sc_hd__a31o_1 _12364_ (.A1(\rbzero.tex_b0[29] ),
    .A2(_04941_),
    .A3(_05549_),
    .B1(_05028_),
    .X(_05550_));
 sky130_fd_sc_hd__a31o_1 _12365_ (.A1(\rbzero.tex_b0[28] ),
    .A2(_04995_),
    .A3(_05431_),
    .B1(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__o221a_1 _12366_ (.A1(_05544_),
    .A2(_05546_),
    .B1(_05548_),
    .B2(_05551_),
    .C1(_04918_),
    .X(_05552_));
 sky130_fd_sc_hd__or2_1 _12367_ (.A(\rbzero.tex_b0[22] ),
    .B(_05498_),
    .X(_05553_));
 sky130_fd_sc_hd__o211a_1 _12368_ (.A1(\rbzero.tex_b0[23] ),
    .A2(_05225_),
    .B1(_05553_),
    .C1(_05293_),
    .X(_05554_));
 sky130_fd_sc_hd__a31o_1 _12369_ (.A1(\rbzero.tex_b0[21] ),
    .A2(_04941_),
    .A3(_05549_),
    .B1(_05028_),
    .X(_05555_));
 sky130_fd_sc_hd__a31o_1 _12370_ (.A1(\rbzero.tex_b0[20] ),
    .A2(_04995_),
    .A3(_05431_),
    .B1(_05555_),
    .X(_05556_));
 sky130_fd_sc_hd__or2_1 _12371_ (.A(\rbzero.tex_b0[18] ),
    .B(_05498_),
    .X(_05557_));
 sky130_fd_sc_hd__o211a_1 _12372_ (.A1(\rbzero.tex_b0[19] ),
    .A2(_05431_),
    .B1(_05557_),
    .C1(_05293_),
    .X(_05558_));
 sky130_fd_sc_hd__clkbuf_4 _12373_ (.A(_04927_),
    .X(_05559_));
 sky130_fd_sc_hd__a31o_1 _12374_ (.A1(\rbzero.tex_b0[17] ),
    .A2(_05559_),
    .A3(_05549_),
    .B1(_04911_),
    .X(_05560_));
 sky130_fd_sc_hd__a31o_1 _12375_ (.A1(\rbzero.tex_b0[16] ),
    .A2(_05389_),
    .A3(_05304_),
    .B1(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__o221a_1 _12376_ (.A1(_05554_),
    .A2(_05556_),
    .B1(_05558_),
    .B2(_05561_),
    .C1(_04987_),
    .X(_05562_));
 sky130_fd_sc_hd__or2_1 _12377_ (.A(\rbzero.tex_b0[6] ),
    .B(_04878_),
    .X(_05563_));
 sky130_fd_sc_hd__o211a_1 _12378_ (.A1(\rbzero.tex_b0[7] ),
    .A2(_04896_),
    .B1(_05563_),
    .C1(_04873_),
    .X(_05564_));
 sky130_fd_sc_hd__a31o_1 _12379_ (.A1(\rbzero.tex_b0[5] ),
    .A2(_05559_),
    .A3(_05549_),
    .B1(_05028_),
    .X(_05565_));
 sky130_fd_sc_hd__a311o_1 _12380_ (.A1(\rbzero.tex_b0[4] ),
    .A2(_04995_),
    .A3(_05225_),
    .B1(_05564_),
    .C1(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__or2_1 _12381_ (.A(\rbzero.tex_b0[2] ),
    .B(_04878_),
    .X(_05567_));
 sky130_fd_sc_hd__o211a_1 _12382_ (.A1(\rbzero.tex_b0[3] ),
    .A2(_04896_),
    .B1(_05567_),
    .C1(_04873_),
    .X(_05568_));
 sky130_fd_sc_hd__a31o_1 _12383_ (.A1(\rbzero.tex_b0[1] ),
    .A2(_05559_),
    .A3(_05549_),
    .B1(_04911_),
    .X(_05569_));
 sky130_fd_sc_hd__a311o_1 _12384_ (.A1(\rbzero.tex_b0[0] ),
    .A2(_04995_),
    .A3(_05225_),
    .B1(_05568_),
    .C1(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__or2_1 _12385_ (.A(\rbzero.tex_b0[10] ),
    .B(_04878_),
    .X(_05571_));
 sky130_fd_sc_hd__o211a_1 _12386_ (.A1(\rbzero.tex_b0[11] ),
    .A2(_05430_),
    .B1(_05571_),
    .C1(_04910_),
    .X(_05572_));
 sky130_fd_sc_hd__a31o_1 _12387_ (.A1(\rbzero.tex_b0[9] ),
    .A2(_04927_),
    .A3(_05035_),
    .B1(_04875_),
    .X(_05573_));
 sky130_fd_sc_hd__a31o_1 _12388_ (.A1(\rbzero.tex_b0[8] ),
    .A2(_05559_),
    .A3(_05430_),
    .B1(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__or2_1 _12389_ (.A(\rbzero.tex_b0[14] ),
    .B(_05035_),
    .X(_05575_));
 sky130_fd_sc_hd__o211a_1 _12390_ (.A1(\rbzero.tex_b0[15] ),
    .A2(_05430_),
    .B1(_05575_),
    .C1(_04910_),
    .X(_05576_));
 sky130_fd_sc_hd__a31o_1 _12391_ (.A1(\rbzero.tex_b0[13] ),
    .A2(_04928_),
    .A3(_05035_),
    .B1(_04944_),
    .X(_05577_));
 sky130_fd_sc_hd__a31o_1 _12392_ (.A1(\rbzero.tex_b0[12] ),
    .A2(_04929_),
    .A3(_05430_),
    .B1(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__o221a_1 _12393_ (.A1(_05572_),
    .A2(_05574_),
    .B1(_05576_),
    .B2(_05578_),
    .C1(_04884_),
    .X(_05579_));
 sky130_fd_sc_hd__a311o_1 _12394_ (.A1(_04987_),
    .A2(_05566_),
    .A3(_05570_),
    .B1(_04951_),
    .C1(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__o311a_1 _12395_ (.A1(_04965_),
    .A2(_05552_),
    .A3(_05562_),
    .B1(_05580_),
    .C1(_04985_),
    .X(_05581_));
 sky130_fd_sc_hd__or2_1 _12396_ (.A(\rbzero.tex_b0[42] ),
    .B(_05498_),
    .X(_05582_));
 sky130_fd_sc_hd__o211a_1 _12397_ (.A1(\rbzero.tex_b0[43] ),
    .A2(_05431_),
    .B1(_05582_),
    .C1(_05293_),
    .X(_05583_));
 sky130_fd_sc_hd__a31o_1 _12398_ (.A1(\rbzero.tex_b0[41] ),
    .A2(_05559_),
    .A3(_05549_),
    .B1(_04911_),
    .X(_05584_));
 sky130_fd_sc_hd__a31o_1 _12399_ (.A1(\rbzero.tex_b0[40] ),
    .A2(_05389_),
    .A3(_05431_),
    .B1(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__or2_1 _12400_ (.A(\rbzero.tex_b0[46] ),
    .B(_05549_),
    .X(_05586_));
 sky130_fd_sc_hd__o211a_1 _12401_ (.A1(\rbzero.tex_b0[47] ),
    .A2(_05431_),
    .B1(_05586_),
    .C1(_05371_),
    .X(_05587_));
 sky130_fd_sc_hd__a31o_1 _12402_ (.A1(\rbzero.tex_b0[45] ),
    .A2(_05559_),
    .A3(_05549_),
    .B1(_05028_),
    .X(_05588_));
 sky130_fd_sc_hd__a31o_1 _12403_ (.A1(\rbzero.tex_b0[44] ),
    .A2(_05389_),
    .A3(_05304_),
    .B1(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__o221a_1 _12404_ (.A1(_05583_),
    .A2(_05585_),
    .B1(_05587_),
    .B2(_05589_),
    .C1(_04918_),
    .X(_05590_));
 sky130_fd_sc_hd__or2_1 _12405_ (.A(\rbzero.tex_b0[38] ),
    .B(_05549_),
    .X(_05591_));
 sky130_fd_sc_hd__o211a_1 _12406_ (.A1(\rbzero.tex_b0[39] ),
    .A2(_05304_),
    .B1(_05591_),
    .C1(_05371_),
    .X(_05592_));
 sky130_fd_sc_hd__a31o_1 _12407_ (.A1(\rbzero.tex_b0[37] ),
    .A2(_05559_),
    .A3(_05244_),
    .B1(_05028_),
    .X(_05593_));
 sky130_fd_sc_hd__a31o_1 _12408_ (.A1(\rbzero.tex_b0[36] ),
    .A2(_05389_),
    .A3(_05304_),
    .B1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__or2_1 _12409_ (.A(\rbzero.tex_b0[34] ),
    .B(_05549_),
    .X(_05595_));
 sky130_fd_sc_hd__o211a_1 _12410_ (.A1(\rbzero.tex_b0[35] ),
    .A2(_05304_),
    .B1(_05595_),
    .C1(_05371_),
    .X(_05596_));
 sky130_fd_sc_hd__a31o_1 _12411_ (.A1(\rbzero.tex_b0[33] ),
    .A2(_04929_),
    .A3(_05244_),
    .B1(_04911_),
    .X(_05597_));
 sky130_fd_sc_hd__a31o_1 _12412_ (.A1(\rbzero.tex_b0[32] ),
    .A2(_05389_),
    .A3(_05304_),
    .B1(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__o221a_1 _12413_ (.A1(_05592_),
    .A2(_05594_),
    .B1(_05596_),
    .B2(_05598_),
    .C1(_04987_),
    .X(_05599_));
 sky130_fd_sc_hd__or2_1 _12414_ (.A(\rbzero.tex_b0[54] ),
    .B(_04878_),
    .X(_05600_));
 sky130_fd_sc_hd__o211a_1 _12415_ (.A1(\rbzero.tex_b0[55] ),
    .A2(_04896_),
    .B1(_05600_),
    .C1(_04873_),
    .X(_05601_));
 sky130_fd_sc_hd__a31o_1 _12416_ (.A1(\rbzero.tex_b0[53] ),
    .A2(_05559_),
    .A3(_05244_),
    .B1(_05028_),
    .X(_05602_));
 sky130_fd_sc_hd__a311o_1 _12417_ (.A1(\rbzero.tex_b0[52] ),
    .A2(_05389_),
    .A3(_05431_),
    .B1(_05601_),
    .C1(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__or2_1 _12418_ (.A(\rbzero.tex_b0[50] ),
    .B(_04878_),
    .X(_05604_));
 sky130_fd_sc_hd__o211a_1 _12419_ (.A1(\rbzero.tex_b0[51] ),
    .A2(_04896_),
    .B1(_05604_),
    .C1(_04873_),
    .X(_05605_));
 sky130_fd_sc_hd__a31o_1 _12420_ (.A1(\rbzero.tex_b0[49] ),
    .A2(_05559_),
    .A3(_05244_),
    .B1(_04911_),
    .X(_05606_));
 sky130_fd_sc_hd__a311o_1 _12421_ (.A1(\rbzero.tex_b0[48] ),
    .A2(_05389_),
    .A3(_05431_),
    .B1(_05605_),
    .C1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__or2_1 _12422_ (.A(\rbzero.tex_b0[58] ),
    .B(_05035_),
    .X(_05608_));
 sky130_fd_sc_hd__o211a_1 _12423_ (.A1(\rbzero.tex_b0[59] ),
    .A2(_05430_),
    .B1(_05608_),
    .C1(_04910_),
    .X(_05609_));
 sky130_fd_sc_hd__a31o_1 _12424_ (.A1(\rbzero.tex_b0[57] ),
    .A2(_04928_),
    .A3(_05035_),
    .B1(_04875_),
    .X(_05610_));
 sky130_fd_sc_hd__a31o_1 _12425_ (.A1(\rbzero.tex_b0[56] ),
    .A2(_04929_),
    .A3(_04925_),
    .B1(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__or2_1 _12426_ (.A(\rbzero.tex_b0[62] ),
    .B(_05035_),
    .X(_05612_));
 sky130_fd_sc_hd__o211a_1 _12427_ (.A1(\rbzero.tex_b0[63] ),
    .A2(_04925_),
    .B1(_05612_),
    .C1(_04910_),
    .X(_05613_));
 sky130_fd_sc_hd__a31o_1 _12428_ (.A1(\rbzero.tex_b0[61] ),
    .A2(_04928_),
    .A3(_05035_),
    .B1(_04944_),
    .X(_05614_));
 sky130_fd_sc_hd__a31o_1 _12429_ (.A1(\rbzero.tex_b0[60] ),
    .A2(_04929_),
    .A3(_04925_),
    .B1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__o221a_1 _12430_ (.A1(_05609_),
    .A2(_05611_),
    .B1(_05613_),
    .B2(_05615_),
    .C1(_04884_),
    .X(_05616_));
 sky130_fd_sc_hd__a311o_1 _12431_ (.A1(_04987_),
    .A2(_05603_),
    .A3(_05607_),
    .B1(_04964_),
    .C1(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__o311a_1 _12432_ (.A1(_05241_),
    .A2(_05590_),
    .A3(_05599_),
    .B1(_05617_),
    .C1(_05023_),
    .X(_05618_));
 sky130_fd_sc_hd__nor2_1 _12433_ (.A(_05581_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__o2bb2a_1 _12434_ (.A1_N(_04907_),
    .A2_N(_05542_),
    .B1(_05619_),
    .B2(_05319_),
    .X(_05620_));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_04808_),
    .X(_05621_));
 sky130_fd_sc_hd__o21ai_1 _12436_ (.A1(_05033_),
    .A2(_05089_),
    .B1(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__o31ai_2 _12437_ (.A1(_05033_),
    .A2(_05089_),
    .A3(_05620_),
    .B1(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__or2_1 _12438_ (.A(_05092_),
    .B(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__o21a_1 _12439_ (.A1(_05342_),
    .A2(_05355_),
    .B1(_05534_),
    .X(_05625_));
 sky130_fd_sc_hd__or3_1 _12440_ (.A(_04764_),
    .B(_04766_),
    .C(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a31o_1 _12441_ (.A1(_05447_),
    .A2(_05624_),
    .A3(_05626_),
    .B1(_04720_),
    .X(_05627_));
 sky130_fd_sc_hd__and2_1 _12442_ (.A(_05096_),
    .B(_05101_),
    .X(_05628_));
 sky130_fd_sc_hd__and3b_2 _12443_ (.A_N(_04721_),
    .B(_05627_),
    .C(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__mux2_2 _12444_ (.A0(\reg_rgb[22] ),
    .A1(_05629_),
    .S(_05103_),
    .X(_05630_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12445_ (.A(_05630_),
    .X(net67));
 sky130_fd_sc_hd__mux2_1 _12446_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_04808_),
    .X(_05631_));
 sky130_fd_sc_hd__o21ai_1 _12447_ (.A1(_04889_),
    .A2(_04880_),
    .B1(\rbzero.row_render.side ),
    .Y(_05632_));
 sky130_fd_sc_hd__o21ai_1 _12448_ (.A1(_04876_),
    .A2(_04889_),
    .B1(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__nand2_1 _12449_ (.A(\rbzero.row_render.wall[1] ),
    .B(_04913_),
    .Y(_05634_));
 sky130_fd_sc_hd__a22o_1 _12450_ (.A1(_04902_),
    .A2(_05633_),
    .B1(_05634_),
    .B2(\rbzero.row_render.wall[0] ),
    .X(_05635_));
 sky130_fd_sc_hd__and3_1 _12451_ (.A(\rbzero.row_render.texu[0] ),
    .B(_04936_),
    .C(_04937_),
    .X(_05636_));
 sky130_fd_sc_hd__o21ai_1 _12452_ (.A1(_04880_),
    .A2(_05636_),
    .B1(_04905_),
    .Y(_05637_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04896_),
    .X(_05638_));
 sky130_fd_sc_hd__mux2_1 _12454_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04939_),
    .X(_05639_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(_05638_),
    .A1(_05639_),
    .S(_04956_),
    .X(_05640_));
 sky130_fd_sc_hd__mux2_1 _12456_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04939_),
    .X(_05641_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04939_),
    .X(_05642_));
 sky130_fd_sc_hd__mux2_1 _12458_ (.A0(_05641_),
    .A1(_05642_),
    .S(_04995_),
    .X(_05643_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(_05640_),
    .A1(_05643_),
    .S(_04932_),
    .X(_05644_));
 sky130_fd_sc_hd__and2_1 _12460_ (.A(\rbzero.tex_b1[62] ),
    .B(_05304_),
    .X(_05645_));
 sky130_fd_sc_hd__a31o_1 _12461_ (.A1(\rbzero.tex_b1[63] ),
    .A2(_04936_),
    .A3(_04937_),
    .B1(_04930_),
    .X(_05646_));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_05431_),
    .X(_05647_));
 sky130_fd_sc_hd__o221a_1 _12463_ (.A1(_05645_),
    .A2(_05646_),
    .B1(_05647_),
    .B2(_05294_),
    .C1(_05238_),
    .X(_05648_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_05430_),
    .X(_05649_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_05430_),
    .X(_05650_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(_05649_),
    .A1(_05650_),
    .S(_05371_),
    .X(_05651_));
 sky130_fd_sc_hd__a21o_1 _12467_ (.A1(_05373_),
    .A2(_05651_),
    .B1(_04987_),
    .X(_05652_));
 sky130_fd_sc_hd__o221a_1 _12468_ (.A1(_05223_),
    .A2(_05644_),
    .B1(_05648_),
    .B2(_05652_),
    .C1(_05241_),
    .X(_05653_));
 sky130_fd_sc_hd__buf_4 _12469_ (.A(_04895_),
    .X(_05654_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_05654_),
    .X(_05656_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(_05655_),
    .A1(_05656_),
    .S(_04930_),
    .X(_05657_));
 sky130_fd_sc_hd__and3_1 _12473_ (.A(\rbzero.tex_b1[39] ),
    .B(_04892_),
    .C(_04893_),
    .X(_05658_));
 sky130_fd_sc_hd__a21o_1 _12474_ (.A1(\rbzero.tex_b1[38] ),
    .A2(_04920_),
    .B1(_04929_),
    .X(_05659_));
 sky130_fd_sc_hd__mux2_1 _12475_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_05654_),
    .X(_05660_));
 sky130_fd_sc_hd__o221a_1 _12476_ (.A1(_05658_),
    .A2(_05659_),
    .B1(_05660_),
    .B2(_05371_),
    .C1(_04960_),
    .X(_05661_));
 sky130_fd_sc_hd__a211o_1 _12477_ (.A1(_04952_),
    .A2(_05657_),
    .B1(_05661_),
    .C1(_04918_),
    .X(_05662_));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_05654_),
    .X(_05663_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_05654_),
    .X(_05664_));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(_05663_),
    .A1(_05664_),
    .S(_05389_),
    .X(_05665_));
 sky130_fd_sc_hd__and2_1 _12481_ (.A(\rbzero.tex_b1[46] ),
    .B(_04925_),
    .X(_05666_));
 sky130_fd_sc_hd__a31o_1 _12482_ (.A1(\rbzero.tex_b1[47] ),
    .A2(_04892_),
    .A3(_04893_),
    .B1(_04929_),
    .X(_05667_));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_05654_),
    .X(_05668_));
 sky130_fd_sc_hd__o221a_1 _12484_ (.A1(_05666_),
    .A2(_05667_),
    .B1(_05668_),
    .B2(_05371_),
    .C1(_04960_),
    .X(_05669_));
 sky130_fd_sc_hd__a211o_1 _12485_ (.A1(_04952_),
    .A2(_05665_),
    .B1(_05669_),
    .C1(_04987_),
    .X(_05670_));
 sky130_fd_sc_hd__a31o_1 _12486_ (.A1(_04965_),
    .A2(_05662_),
    .A3(_05670_),
    .B1(_04985_),
    .X(_05671_));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_05654_),
    .X(_05672_));
 sky130_fd_sc_hd__or2_1 _12488_ (.A(_04930_),
    .B(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__mux2_1 _12489_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_05430_),
    .X(_05674_));
 sky130_fd_sc_hd__o21a_1 _12490_ (.A1(_05371_),
    .A2(_05674_),
    .B1(_04945_),
    .X(_05675_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04896_),
    .X(_05676_));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04896_),
    .X(_05677_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(_05676_),
    .A1(_05677_),
    .S(_05293_),
    .X(_05678_));
 sky130_fd_sc_hd__a221o_1 _12494_ (.A1(_05673_),
    .A2(_05675_),
    .B1(_05678_),
    .B2(_05238_),
    .C1(_04918_),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_05430_),
    .X(_05680_));
 sky130_fd_sc_hd__mux2_1 _12496_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_05654_),
    .X(_05681_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(_05680_),
    .A1(_05681_),
    .S(_04930_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _12498_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_05654_),
    .X(_05683_));
 sky130_fd_sc_hd__and2_1 _12499_ (.A(\rbzero.tex_b1[30] ),
    .B(_04925_),
    .X(_05684_));
 sky130_fd_sc_hd__a31o_1 _12500_ (.A1(\rbzero.tex_b1[31] ),
    .A2(_04892_),
    .A3(_04893_),
    .B1(_04929_),
    .X(_05685_));
 sky130_fd_sc_hd__o221a_1 _12501_ (.A1(_05371_),
    .A2(_05683_),
    .B1(_05684_),
    .B2(_05685_),
    .C1(_04960_),
    .X(_05686_));
 sky130_fd_sc_hd__a211o_1 _12502_ (.A1(_05373_),
    .A2(_05682_),
    .B1(_05686_),
    .C1(_04987_),
    .X(_05687_));
 sky130_fd_sc_hd__mux2_1 _12503_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_04895_),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_1 _12504_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_04895_),
    .X(_05689_));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(_05688_),
    .A1(_05689_),
    .S(_04873_),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_1 _12506_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04895_),
    .X(_05691_));
 sky130_fd_sc_hd__mux2_1 _12507_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04895_),
    .X(_05692_));
 sky130_fd_sc_hd__mux2_1 _12508_ (.A0(_05691_),
    .A1(_05692_),
    .S(_05559_),
    .X(_05693_));
 sky130_fd_sc_hd__mux2_1 _12509_ (.A0(_05690_),
    .A1(_05693_),
    .S(_04960_),
    .X(_05694_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_05654_),
    .X(_05695_));
 sky130_fd_sc_hd__and2_1 _12511_ (.A(\rbzero.tex_b1[14] ),
    .B(_04920_),
    .X(_05696_));
 sky130_fd_sc_hd__a31o_1 _12512_ (.A1(\rbzero.tex_b1[15] ),
    .A2(_04892_),
    .A3(_04893_),
    .B1(_05027_),
    .X(_05697_));
 sky130_fd_sc_hd__o221a_1 _12513_ (.A1(_05371_),
    .A2(_05695_),
    .B1(_05696_),
    .B2(_05697_),
    .C1(_04960_),
    .X(_05698_));
 sky130_fd_sc_hd__mux2_1 _12514_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04895_),
    .X(_05699_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04895_),
    .X(_05700_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(_05699_),
    .A1(_05700_),
    .S(_04929_),
    .X(_05701_));
 sky130_fd_sc_hd__a21o_1 _12517_ (.A1(_04946_),
    .A2(_05701_),
    .B1(_04908_),
    .X(_05702_));
 sky130_fd_sc_hd__o221a_1 _12518_ (.A1(_04918_),
    .A2(_05694_),
    .B1(_05698_),
    .B2(_05702_),
    .C1(_04964_),
    .X(_05703_));
 sky130_fd_sc_hd__a31o_1 _12519_ (.A1(_05241_),
    .A2(_05679_),
    .A3(_05687_),
    .B1(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__o221a_2 _12520_ (.A1(_05653_),
    .A2(_05671_),
    .B1(_05704_),
    .B2(_05023_),
    .C1(_04906_),
    .X(_05705_));
 sky130_fd_sc_hd__a31o_1 _12521_ (.A1(_05319_),
    .A2(_05635_),
    .A3(_05637_),
    .B1(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__mux2_1 _12522_ (.A0(_05631_),
    .A1(_05706_),
    .S(_05090_),
    .X(_05707_));
 sky130_fd_sc_hd__a31o_1 _12523_ (.A1(_05092_),
    .A2(_05330_),
    .A3(_05625_),
    .B1(_04720_),
    .X(_05708_));
 sky130_fd_sc_hd__a21o_1 _12524_ (.A1(_04764_),
    .A2(_05707_),
    .B1(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__and3b_2 _12525_ (.A_N(_05222_),
    .B(_05628_),
    .C(_05709_),
    .X(_05710_));
 sky130_fd_sc_hd__mux2_2 _12526_ (.A0(\reg_rgb[23] ),
    .A1(_05710_),
    .S(_05103_),
    .X(_05711_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12527_ (.A(_05711_),
    .X(net68));
 sky130_fd_sc_hd__mux2_4 _12528_ (.A0(reg_vsync),
    .A1(_04488_),
    .S(_05103_),
    .X(_05712_));
 sky130_fd_sc_hd__clkbuf_1 _12529_ (.A(_05712_),
    .X(net75));
 sky130_fd_sc_hd__inv_2 _12530_ (.A(\rbzero.hsync ),
    .Y(_05713_));
 sky130_fd_sc_hd__mux2_2 _12531_ (.A0(reg_hsync),
    .A1(_05713_),
    .S(_05103_),
    .X(_05714_));
 sky130_fd_sc_hd__clkbuf_1 _12532_ (.A(_05714_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 _12533_ (.A(net4),
    .X(_05715_));
 sky130_fd_sc_hd__or2_1 _12534_ (.A(_05715_),
    .B(_05102_),
    .X(_05716_));
 sky130_fd_sc_hd__inv_2 _12535_ (.A(net7),
    .Y(_05717_));
 sky130_fd_sc_hd__nor2_1 _12536_ (.A(_05717_),
    .B(net8),
    .Y(_05718_));
 sky130_fd_sc_hd__nand2_1 _12537_ (.A(_05715_),
    .B(_05363_),
    .Y(_05719_));
 sky130_fd_sc_hd__mux4_1 _12538_ (.A0(_05450_),
    .A1(_05539_),
    .A2(_05629_),
    .A3(_05710_),
    .S0(_05715_),
    .S1(net7),
    .X(_05720_));
 sky130_fd_sc_hd__a32o_1 _12539_ (.A1(_05716_),
    .A2(_05718_),
    .A3(_05719_),
    .B1(_05720_),
    .B2(net8),
    .X(_05721_));
 sky130_fd_sc_hd__and4b_1 _12540_ (.A_N(net9),
    .B(_05721_),
    .C(net5),
    .D(net6),
    .X(_05722_));
 sky130_fd_sc_hd__and2b_1 _12541_ (.A_N(net8),
    .B(net9),
    .X(_05723_));
 sky130_fd_sc_hd__inv_2 _12542_ (.A(net6),
    .Y(_05724_));
 sky130_fd_sc_hd__nor2_1 _12543_ (.A(net7),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__and2b_1 _12544_ (.A_N(net5),
    .B(net4),
    .X(_05726_));
 sky130_fd_sc_hd__nor2_1 _12545_ (.A(net5),
    .B(net4),
    .Y(_05727_));
 sky130_fd_sc_hd__a22o_1 _12546_ (.A1(net72),
    .A2(_05726_),
    .B1(_05727_),
    .B2(_05100_),
    .X(_05728_));
 sky130_fd_sc_hd__and2_1 _12547_ (.A(net5),
    .B(net4),
    .X(_05729_));
 sky130_fd_sc_hd__and2b_1 _12548_ (.A_N(net4),
    .B(net5),
    .X(_05730_));
 sky130_fd_sc_hd__a22o_1 _12549_ (.A1(_05098_),
    .A2(_05729_),
    .B1(_05730_),
    .B2(net44),
    .X(_05731_));
 sky130_fd_sc_hd__nor2_1 _12550_ (.A(net7),
    .B(net6),
    .Y(_05732_));
 sky130_fd_sc_hd__a22o_1 _12551_ (.A1(_05725_),
    .A2(_05728_),
    .B1(_05731_),
    .B2(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__buf_4 _12552_ (.A(net55),
    .X(_05734_));
 sky130_fd_sc_hd__nor2_1 _12553_ (.A(net9),
    .B(net8),
    .Y(_05735_));
 sky130_fd_sc_hd__a41o_1 _12554_ (.A1(_05734_),
    .A2(_05729_),
    .A3(_05735_),
    .A4(_05725_),
    .B1(_05723_),
    .X(_05736_));
 sky130_fd_sc_hd__a22o_1 _12555_ (.A1(_05319_),
    .A2(_05729_),
    .B1(_05730_),
    .B2(net41),
    .X(_05737_));
 sky130_fd_sc_hd__a22o_1 _12556_ (.A1(net40),
    .A2(_05726_),
    .B1(_05727_),
    .B2(net52),
    .X(_05738_));
 sky130_fd_sc_hd__or3_1 _12557_ (.A(_05717_),
    .B(_05737_),
    .C(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__a221o_1 _12558_ (.A1(net46),
    .A2(_05726_),
    .B1(_05727_),
    .B2(net43),
    .C1(net7),
    .X(_05740_));
 sky130_fd_sc_hd__a21o_1 _12559_ (.A1(_05734_),
    .A2(_05735_),
    .B1(net51),
    .X(_05741_));
 sky130_fd_sc_hd__a22o_1 _12560_ (.A1(net50),
    .A2(_05730_),
    .B1(_05741_),
    .B2(_05729_),
    .X(_05742_));
 sky130_fd_sc_hd__a32o_1 _12561_ (.A1(_05724_),
    .A2(_05739_),
    .A3(_05740_),
    .B1(_05725_),
    .B2(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__a22o_1 _12562_ (.A1(net54),
    .A2(_05726_),
    .B1(_05727_),
    .B2(net53),
    .X(_05744_));
 sky130_fd_sc_hd__a21o_1 _12563_ (.A1(net56),
    .A2(_05730_),
    .B1(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__a21oi_2 _12564_ (.A1(net128),
    .A2(net5),
    .B1(_05715_),
    .Y(_05746_));
 sky130_fd_sc_hd__a221o_2 _12565_ (.A1(_04468_),
    .A2(_05726_),
    .B1(_05729_),
    .B2(\gpout0.clk_div[1] ),
    .C1(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__a22o_2 _12566_ (.A1(_05725_),
    .A2(_05745_),
    .B1(_05747_),
    .B2(_05732_),
    .X(_05748_));
 sky130_fd_sc_hd__a22o_2 _12567_ (.A1(_05736_),
    .A2(_05743_),
    .B1(_05748_),
    .B2(_05735_),
    .X(_05749_));
 sky130_fd_sc_hd__a21oi_1 _12568_ (.A1(net5),
    .A2(net6),
    .B1(net7),
    .Y(_05750_));
 sky130_fd_sc_hd__and3b_1 _12569_ (.A_N(_05750_),
    .B(net8),
    .C(net9),
    .X(_05751_));
 sky130_fd_sc_hd__buf_2 _12570_ (.A(\gpout0.vpos[2] ),
    .X(_05752_));
 sky130_fd_sc_hd__buf_2 _12571_ (.A(_04723_),
    .X(_05753_));
 sky130_fd_sc_hd__mux2_1 _12572_ (.A0(_05752_),
    .A1(_05753_),
    .S(_05715_),
    .X(_05754_));
 sky130_fd_sc_hd__buf_2 _12573_ (.A(_04718_),
    .X(_05755_));
 sky130_fd_sc_hd__buf_2 _12574_ (.A(_04714_),
    .X(_05756_));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(_05755_),
    .A1(_05756_),
    .S(_05715_),
    .X(_05757_));
 sky130_fd_sc_hd__clkbuf_4 _12576_ (.A(_04701_),
    .X(_05758_));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(_05758_),
    .A1(_04704_),
    .S(_05715_),
    .X(_05759_));
 sky130_fd_sc_hd__buf_2 _12578_ (.A(\gpout0.vpos[0] ),
    .X(_05760_));
 sky130_fd_sc_hd__buf_2 _12579_ (.A(\gpout0.vpos[8] ),
    .X(_05761_));
 sky130_fd_sc_hd__buf_2 _12580_ (.A(\gpout0.vpos[9] ),
    .X(_05762_));
 sky130_fd_sc_hd__mux4_1 _12581_ (.A0(_05760_),
    .A1(_04744_),
    .A2(_05761_),
    .A3(_05762_),
    .S0(_05715_),
    .S1(net7),
    .X(_05763_));
 sky130_fd_sc_hd__mux4_1 _12582_ (.A0(_05754_),
    .A1(_05757_),
    .A2(_05759_),
    .A3(_05763_),
    .S0(net6),
    .S1(net5),
    .X(_05764_));
 sky130_fd_sc_hd__mux4_1 _12583_ (.A0(_04643_),
    .A1(_05105_),
    .A2(_04481_),
    .A3(_04032_),
    .S0(_05715_),
    .S1(net5),
    .X(_05765_));
 sky130_fd_sc_hd__or2_1 _12584_ (.A(net6),
    .B(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(_04033_),
    .A1(_04034_),
    .S(_05715_),
    .X(_05767_));
 sky130_fd_sc_hd__mux4_1 _12586_ (.A0(\gpout0.hpos[0] ),
    .A1(_04507_),
    .A2(_04506_),
    .A3(_04513_),
    .S0(net4),
    .S1(net5),
    .X(_05768_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(_05767_),
    .A1(_05768_),
    .S(net7),
    .X(_05769_));
 sky130_fd_sc_hd__a22o_1 _12588_ (.A1(net6),
    .A2(_05718_),
    .B1(_05750_),
    .B2(net8),
    .X(_05770_));
 sky130_fd_sc_hd__o211a_1 _12589_ (.A1(_05724_),
    .A2(_05769_),
    .B1(_05770_),
    .C1(net9),
    .X(_05771_));
 sky130_fd_sc_hd__a22o_1 _12590_ (.A1(_05751_),
    .A2(_05764_),
    .B1(_05766_),
    .B2(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__a211o_2 _12591_ (.A1(_05723_),
    .A2(_05733_),
    .B1(_05749_),
    .C1(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__nand3_1 _12592_ (.A(_05727_),
    .B(_05735_),
    .C(_05732_),
    .Y(_05774_));
 sky130_fd_sc_hd__o22a_2 _12593_ (.A1(_05722_),
    .A2(_05773_),
    .B1(_05774_),
    .B2(_05450_),
    .X(_05775_));
 sky130_fd_sc_hd__mux2_2 _12594_ (.A0(\reg_gpout[0] ),
    .A1(clknet_1_1__leaf__05775_),
    .S(_05103_),
    .X(_05776_));
 sky130_fd_sc_hd__buf_1 _12595_ (.A(_05776_),
    .X(net57));
 sky130_fd_sc_hd__inv_2 _12596_ (.A(net14),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_1 _12597_ (.A(net13),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__inv_2 _12598_ (.A(_05102_),
    .Y(_05779_));
 sky130_fd_sc_hd__clkbuf_4 _12599_ (.A(net10),
    .X(_05780_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(_05779_),
    .A1(_05363_),
    .S(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__mux4_1 _12601_ (.A0(_05450_),
    .A1(_05539_),
    .A2(_05629_),
    .A3(_05710_),
    .S0(_05780_),
    .S1(net13),
    .X(_05782_));
 sky130_fd_sc_hd__a2bb2o_1 _12602_ (.A1_N(_05778_),
    .A2_N(_05781_),
    .B1(net14),
    .B2(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__and4b_1 _12603_ (.A_N(net15),
    .B(_05783_),
    .C(net11),
    .D(net12),
    .X(_05784_));
 sky130_fd_sc_hd__inv_2 _12604_ (.A(net12),
    .Y(_05785_));
 sky130_fd_sc_hd__nor2_1 _12605_ (.A(net13),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__and2b_1 _12606_ (.A_N(net11),
    .B(net10),
    .X(_05787_));
 sky130_fd_sc_hd__nor2_1 _12607_ (.A(net11),
    .B(_05780_),
    .Y(_05788_));
 sky130_fd_sc_hd__a22o_1 _12608_ (.A1(net72),
    .A2(_05787_),
    .B1(_05788_),
    .B2(_05100_),
    .X(_05789_));
 sky130_fd_sc_hd__and2_1 _12609_ (.A(net11),
    .B(_05780_),
    .X(_05790_));
 sky130_fd_sc_hd__nor2_1 _12610_ (.A(net13),
    .B(net12),
    .Y(_05791_));
 sky130_fd_sc_hd__and3_1 _12611_ (.A(_05098_),
    .B(_05790_),
    .C(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__and2b_1 _12612_ (.A_N(net10),
    .B(net11),
    .X(_05793_));
 sky130_fd_sc_hd__and3_1 _12613_ (.A(net44),
    .B(_05793_),
    .C(_05791_),
    .X(_05794_));
 sky130_fd_sc_hd__a211o_1 _12614_ (.A1(_05786_),
    .A2(_05789_),
    .B1(_05792_),
    .C1(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__and2_1 _12615_ (.A(_05777_),
    .B(net15),
    .X(_05796_));
 sky130_fd_sc_hd__nor2_1 _12616_ (.A(net14),
    .B(net15),
    .Y(_05797_));
 sky130_fd_sc_hd__a21o_1 _12617_ (.A1(_05734_),
    .A2(_05797_),
    .B1(net51),
    .X(_05798_));
 sky130_fd_sc_hd__a22o_1 _12618_ (.A1(_05790_),
    .A2(_05798_),
    .B1(_05793_),
    .B2(net50),
    .X(_05799_));
 sky130_fd_sc_hd__a22o_1 _12619_ (.A1(net46),
    .A2(_05787_),
    .B1(_05788_),
    .B2(net43),
    .X(_05800_));
 sky130_fd_sc_hd__a22o_1 _12620_ (.A1(net40),
    .A2(_05787_),
    .B1(_05788_),
    .B2(net52),
    .X(_05801_));
 sky130_fd_sc_hd__a221o_1 _12621_ (.A1(_05319_),
    .A2(_05790_),
    .B1(_05793_),
    .B2(net41),
    .C1(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__mux2_1 _12622_ (.A0(_05800_),
    .A1(_05802_),
    .S(net13),
    .X(_05803_));
 sky130_fd_sc_hd__a22o_1 _12623_ (.A1(_05799_),
    .A2(_05786_),
    .B1(_05803_),
    .B2(_05785_),
    .X(_05804_));
 sky130_fd_sc_hd__a41o_1 _12624_ (.A1(_05734_),
    .A2(_05790_),
    .A3(_05797_),
    .A4(_05786_),
    .B1(_05796_),
    .X(_05805_));
 sky130_fd_sc_hd__a21o_1 _12625_ (.A1(net11),
    .A2(net12),
    .B1(net13),
    .X(_05806_));
 sky130_fd_sc_hd__mux2_1 _12626_ (.A0(_05752_),
    .A1(_04723_),
    .S(_05780_),
    .X(_05807_));
 sky130_fd_sc_hd__mux2_1 _12627_ (.A0(_05755_),
    .A1(_05756_),
    .S(_05780_),
    .X(_05808_));
 sky130_fd_sc_hd__mux2_1 _12628_ (.A0(_04701_),
    .A1(_04704_),
    .S(_05780_),
    .X(_05809_));
 sky130_fd_sc_hd__mux4_1 _12629_ (.A0(_05760_),
    .A1(_04744_),
    .A2(_05761_),
    .A3(_05762_),
    .S0(_05780_),
    .S1(net13),
    .X(_05810_));
 sky130_fd_sc_hd__mux4_1 _12630_ (.A0(_05807_),
    .A1(_05808_),
    .A2(_05809_),
    .A3(_05810_),
    .S0(net12),
    .S1(net11),
    .X(_05811_));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(_04033_),
    .A1(_04034_),
    .S(_05780_),
    .X(_05812_));
 sky130_fd_sc_hd__mux4_1 _12632_ (.A0(\gpout0.hpos[0] ),
    .A1(_04507_),
    .A2(\gpout0.hpos[2] ),
    .A3(_04513_),
    .S0(net10),
    .S1(net11),
    .X(_05813_));
 sky130_fd_sc_hd__mux2_1 _12633_ (.A0(_05812_),
    .A1(_05813_),
    .S(net13),
    .X(_05814_));
 sky130_fd_sc_hd__mux4_1 _12634_ (.A0(_04643_),
    .A1(_05105_),
    .A2(_04481_),
    .A3(_04032_),
    .S0(_05780_),
    .S1(net11),
    .X(_05815_));
 sky130_fd_sc_hd__or2_1 _12635_ (.A(net12),
    .B(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__o22ai_1 _12636_ (.A1(_05785_),
    .A2(_05778_),
    .B1(_05806_),
    .B2(_05777_),
    .Y(_05817_));
 sky130_fd_sc_hd__o2111a_1 _12637_ (.A1(_05785_),
    .A2(_05814_),
    .B1(_05816_),
    .C1(_05817_),
    .D1(net15),
    .X(_05818_));
 sky130_fd_sc_hd__a41o_1 _12638_ (.A1(net14),
    .A2(net15),
    .A3(_05806_),
    .A4(_05811_),
    .B1(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__and2_1 _12639_ (.A(_05788_),
    .B(_05791_),
    .X(_05820_));
 sky130_fd_sc_hd__and3_1 _12640_ (.A(net49),
    .B(_05787_),
    .C(_05791_),
    .X(_05821_));
 sky130_fd_sc_hd__a22o_1 _12641_ (.A1(net56),
    .A2(_05793_),
    .B1(_05787_),
    .B2(net54),
    .X(_05822_));
 sky130_fd_sc_hd__a21o_1 _12642_ (.A1(net53),
    .A2(_05788_),
    .B1(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__and3_1 _12643_ (.A(\gpout1.clk_div[1] ),
    .B(_05790_),
    .C(_05791_),
    .X(_05824_));
 sky130_fd_sc_hd__buf_1 _12644_ (.A(clknet_leaf_44_i_clk),
    .X(_05825_));
 sky130_fd_sc_hd__and3_2 _12645_ (.A(clknet_1_0__leaf__05825_),
    .B(_05793_),
    .C(_05791_),
    .X(_05826_));
 sky130_fd_sc_hd__a211o_2 _12646_ (.A1(_05786_),
    .A2(_05823_),
    .B1(_05824_),
    .C1(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__o31a_2 _12647_ (.A1(_05820_),
    .A2(_05821_),
    .A3(_05827_),
    .B1(_05797_),
    .X(_05828_));
 sky130_fd_sc_hd__a211o_2 _12648_ (.A1(_05804_),
    .A2(_05805_),
    .B1(_05819_),
    .C1(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__a21o_2 _12649_ (.A1(_05795_),
    .A2(_05796_),
    .B1(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__nand2_1 _12650_ (.A(_05797_),
    .B(_05820_),
    .Y(_05831_));
 sky130_fd_sc_hd__o22a_2 _12651_ (.A1(_05784_),
    .A2(_05830_),
    .B1(_05831_),
    .B2(_05539_),
    .X(_05832_));
 sky130_fd_sc_hd__mux2_2 _12652_ (.A0(\reg_gpout[1] ),
    .A1(clknet_1_1__leaf__05832_),
    .S(_05103_),
    .X(_05833_));
 sky130_fd_sc_hd__buf_1 _12653_ (.A(_05833_),
    .X(net58));
 sky130_fd_sc_hd__nor2_1 _12654_ (.A(net21),
    .B(net20),
    .Y(_05834_));
 sky130_fd_sc_hd__buf_2 _12655_ (.A(net17),
    .X(_05835_));
 sky130_fd_sc_hd__clkbuf_4 _12656_ (.A(net16),
    .X(_05836_));
 sky130_fd_sc_hd__nor2_1 _12657_ (.A(_05835_),
    .B(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__nor2_1 _12658_ (.A(net19),
    .B(net18),
    .Y(_05838_));
 sky130_fd_sc_hd__and2_1 _12659_ (.A(_05837_),
    .B(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__inv_2 _12660_ (.A(net19),
    .Y(_05840_));
 sky130_fd_sc_hd__mux2_1 _12661_ (.A0(_05779_),
    .A1(_05363_),
    .S(_05836_),
    .X(_05841_));
 sky130_fd_sc_hd__mux4_1 _12662_ (.A0(_05450_),
    .A1(_05539_),
    .A2(_05629_),
    .A3(_05710_),
    .S0(_05836_),
    .S1(net19),
    .X(_05842_));
 sky130_fd_sc_hd__nand2_1 _12663_ (.A(net20),
    .B(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__o31a_1 _12664_ (.A1(_05840_),
    .A2(net20),
    .A3(_05841_),
    .B1(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__buf_2 _12665_ (.A(net18),
    .X(_05845_));
 sky130_fd_sc_hd__or4bb_1 _12666_ (.A(net21),
    .B(_05844_),
    .C_N(_05835_),
    .D_N(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__inv_2 _12667_ (.A(net20),
    .Y(_05847_));
 sky130_fd_sc_hd__and2b_1 _12668_ (.A_N(_05835_),
    .B(net16),
    .X(_05848_));
 sky130_fd_sc_hd__a22o_1 _12669_ (.A1(_05100_),
    .A2(_05837_),
    .B1(_05848_),
    .B2(net72),
    .X(_05849_));
 sky130_fd_sc_hd__and2b_1 _12670_ (.A_N(net16),
    .B(net17),
    .X(_05850_));
 sky130_fd_sc_hd__and3_1 _12671_ (.A(_05835_),
    .B(net16),
    .C(_05838_),
    .X(_05851_));
 sky130_fd_sc_hd__a32o_1 _12672_ (.A1(net44),
    .A2(_05838_),
    .A3(_05850_),
    .B1(_05851_),
    .B2(_05098_),
    .X(_05852_));
 sky130_fd_sc_hd__a31o_1 _12673_ (.A1(_05840_),
    .A2(_05845_),
    .A3(_05849_),
    .B1(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__nand2_1 _12674_ (.A(_05835_),
    .B(_05836_),
    .Y(_05854_));
 sky130_fd_sc_hd__nand2_1 _12675_ (.A(_05734_),
    .B(_05834_),
    .Y(_05855_));
 sky130_fd_sc_hd__nand2_1 _12676_ (.A(_05840_),
    .B(_05845_),
    .Y(_05856_));
 sky130_fd_sc_hd__inv_2 _12677_ (.A(net21),
    .Y(_05857_));
 sky130_fd_sc_hd__o32a_1 _12678_ (.A1(_05854_),
    .A2(_05855_),
    .A3(_05856_),
    .B1(net20),
    .B2(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__a21oi_1 _12679_ (.A1(_05734_),
    .A2(_05834_),
    .B1(net51),
    .Y(_05859_));
 sky130_fd_sc_hd__o2bb2a_1 _12680_ (.A1_N(net50),
    .A2_N(_05850_),
    .B1(_05854_),
    .B2(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__mux4_1 _12681_ (.A0(net52),
    .A1(net41),
    .A2(net40),
    .A3(_05319_),
    .S0(_05835_),
    .S1(_05836_),
    .X(_05861_));
 sky130_fd_sc_hd__a221o_1 _12682_ (.A1(net43),
    .A2(_05837_),
    .B1(_05848_),
    .B2(net46),
    .C1(net19),
    .X(_05862_));
 sky130_fd_sc_hd__o21ai_1 _12683_ (.A1(_05840_),
    .A2(_05861_),
    .B1(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__o22a_1 _12684_ (.A1(_05860_),
    .A2(_05856_),
    .B1(_05863_),
    .B2(_05845_),
    .X(_05864_));
 sky130_fd_sc_hd__a22o_1 _12685_ (.A1(net53),
    .A2(_05837_),
    .B1(_05850_),
    .B2(net56),
    .X(_05865_));
 sky130_fd_sc_hd__a21o_1 _12686_ (.A1(net54),
    .A2(_05848_),
    .B1(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__a32o_2 _12687_ (.A1(clknet_1_0__leaf__05825_),
    .A2(_05838_),
    .A3(_05850_),
    .B1(_05851_),
    .B2(\gpout2.clk_div[1] ),
    .X(_05867_));
 sky130_fd_sc_hd__a311o_2 _12688_ (.A1(net47),
    .A2(_05838_),
    .A3(_05848_),
    .B1(_05867_),
    .C1(_05839_),
    .X(_05868_));
 sky130_fd_sc_hd__a31o_2 _12689_ (.A1(_05840_),
    .A2(_05845_),
    .A3(_05866_),
    .B1(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__a2bb2o_2 _12690_ (.A1_N(_05858_),
    .A2_N(_05864_),
    .B1(_05869_),
    .B2(_05834_),
    .X(_05870_));
 sky130_fd_sc_hd__a21o_1 _12691_ (.A1(_05835_),
    .A2(_05845_),
    .B1(net19),
    .X(_05871_));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(_05752_),
    .A1(_05753_),
    .S(_05836_),
    .X(_05872_));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(_05755_),
    .A1(_05756_),
    .S(_05836_),
    .X(_05873_));
 sky130_fd_sc_hd__mux2_1 _12694_ (.A0(_05758_),
    .A1(_04704_),
    .S(_05836_),
    .X(_05874_));
 sky130_fd_sc_hd__mux4_1 _12695_ (.A0(_05760_),
    .A1(_04744_),
    .A2(_05761_),
    .A3(_05762_),
    .S0(_05836_),
    .S1(net19),
    .X(_05875_));
 sky130_fd_sc_hd__mux4_1 _12696_ (.A0(_05872_),
    .A1(_05873_),
    .A2(_05874_),
    .A3(_05875_),
    .S0(_05845_),
    .S1(_05835_),
    .X(_05876_));
 sky130_fd_sc_hd__mux4_1 _12697_ (.A0(_04643_),
    .A1(_05105_),
    .A2(_04481_),
    .A3(_04032_),
    .S0(_05836_),
    .S1(_05835_),
    .X(_05877_));
 sky130_fd_sc_hd__mux2_1 _12698_ (.A0(_04033_),
    .A1(_04034_),
    .S(net16),
    .X(_05878_));
 sky130_fd_sc_hd__mux4_1 _12699_ (.A0(\gpout0.hpos[0] ),
    .A1(_04507_),
    .A2(\gpout0.hpos[2] ),
    .A3(_04513_),
    .S0(net16),
    .S1(_05835_),
    .X(_05879_));
 sky130_fd_sc_hd__mux2_1 _12700_ (.A0(_05878_),
    .A1(_05879_),
    .S(net19),
    .X(_05880_));
 sky130_fd_sc_hd__or2b_1 _12701_ (.A(_05880_),
    .B_N(_05845_),
    .X(_05881_));
 sky130_fd_sc_hd__nor2_1 _12702_ (.A(_05847_),
    .B(_05871_),
    .Y(_05882_));
 sky130_fd_sc_hd__a31o_1 _12703_ (.A1(net19),
    .A2(_05845_),
    .A3(_05847_),
    .B1(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__o2111a_1 _12704_ (.A1(_05845_),
    .A2(_05877_),
    .B1(_05881_),
    .C1(net21),
    .D1(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__a41o_1 _12705_ (.A1(net21),
    .A2(net20),
    .A3(_05871_),
    .A4(_05876_),
    .B1(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__a311oi_2 _12706_ (.A1(net21),
    .A2(_05847_),
    .A3(_05853_),
    .B1(_05870_),
    .C1(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__a32oi_2 _12707_ (.A1(_05779_),
    .A2(_05834_),
    .A3(_05839_),
    .B1(_05846_),
    .B2(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__mux2_2 _12708_ (.A0(\reg_gpout[2] ),
    .A1(clknet_1_1__leaf__05887_),
    .S(net45),
    .X(_05888_));
 sky130_fd_sc_hd__buf_1 _12709_ (.A(_05888_),
    .X(net59));
 sky130_fd_sc_hd__nor2_1 _12710_ (.A(net27),
    .B(net26),
    .Y(_05889_));
 sky130_fd_sc_hd__nor2_1 _12711_ (.A(net23),
    .B(net22),
    .Y(_05890_));
 sky130_fd_sc_hd__nor2_1 _12712_ (.A(net25),
    .B(net24),
    .Y(_05891_));
 sky130_fd_sc_hd__and3_1 _12713_ (.A(_05889_),
    .B(_05890_),
    .C(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__inv_2 _12714_ (.A(net24),
    .Y(_05893_));
 sky130_fd_sc_hd__nor2_1 _12715_ (.A(net25),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__inv_2 _12716_ (.A(net22),
    .Y(_05895_));
 sky130_fd_sc_hd__nor2_1 _12717_ (.A(net23),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__a22o_1 _12718_ (.A1(net72),
    .A2(_05896_),
    .B1(_05890_),
    .B2(_05100_),
    .X(_05897_));
 sky130_fd_sc_hd__and3_1 _12719_ (.A(net23),
    .B(net22),
    .C(_05891_),
    .X(_05898_));
 sky130_fd_sc_hd__inv_2 _12720_ (.A(net23),
    .Y(_05899_));
 sky130_fd_sc_hd__nor2_1 _12721_ (.A(_05899_),
    .B(net22),
    .Y(_05900_));
 sky130_fd_sc_hd__and3_1 _12722_ (.A(net44),
    .B(_05900_),
    .C(_05891_),
    .X(_05901_));
 sky130_fd_sc_hd__a221o_1 _12723_ (.A1(_05894_),
    .A2(_05897_),
    .B1(_05898_),
    .B2(_05098_),
    .C1(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__and2b_1 _12724_ (.A_N(net26),
    .B(net27),
    .X(_05903_));
 sky130_fd_sc_hd__clkbuf_4 _12725_ (.A(net22),
    .X(_05904_));
 sky130_fd_sc_hd__or2_1 _12726_ (.A(_05904_),
    .B(_05102_),
    .X(_05905_));
 sky130_fd_sc_hd__and2b_1 _12727_ (.A_N(net26),
    .B(net25),
    .X(_05906_));
 sky130_fd_sc_hd__nand2_1 _12728_ (.A(_05904_),
    .B(_05363_),
    .Y(_05907_));
 sky130_fd_sc_hd__mux4_1 _12729_ (.A0(_05450_),
    .A1(_05539_),
    .A2(_05629_),
    .A3(_05710_),
    .S0(_05904_),
    .S1(net25),
    .X(_05908_));
 sky130_fd_sc_hd__a32o_1 _12730_ (.A1(_05905_),
    .A2(_05906_),
    .A3(_05907_),
    .B1(_05908_),
    .B2(net26),
    .X(_05909_));
 sky130_fd_sc_hd__and4b_1 _12731_ (.A_N(net27),
    .B(_05909_),
    .C(net23),
    .D(net24),
    .X(_05910_));
 sky130_fd_sc_hd__a21o_1 _12732_ (.A1(_05902_),
    .A2(_05903_),
    .B1(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__a21oi_1 _12733_ (.A1(net23),
    .A2(net24),
    .B1(net25),
    .Y(_05912_));
 sky130_fd_sc_hd__and3b_1 _12734_ (.A_N(_05912_),
    .B(net26),
    .C(net27),
    .X(_05913_));
 sky130_fd_sc_hd__mux2_1 _12735_ (.A0(_05758_),
    .A1(_04704_),
    .S(_05904_),
    .X(_05914_));
 sky130_fd_sc_hd__mux4_1 _12736_ (.A0(_05760_),
    .A1(_04744_),
    .A2(_05761_),
    .A3(_05762_),
    .S0(_05904_),
    .S1(net25),
    .X(_05915_));
 sky130_fd_sc_hd__mux2_1 _12737_ (.A0(_05752_),
    .A1(_05753_),
    .S(_05904_),
    .X(_05916_));
 sky130_fd_sc_hd__mux2_1 _12738_ (.A0(_05755_),
    .A1(_05756_),
    .S(_05904_),
    .X(_05917_));
 sky130_fd_sc_hd__mux4_1 _12739_ (.A0(_05914_),
    .A1(_05915_),
    .A2(_05916_),
    .A3(_05917_),
    .S0(net24),
    .S1(_05899_),
    .X(_05918_));
 sky130_fd_sc_hd__mux2_1 _12740_ (.A0(_04033_),
    .A1(_04034_),
    .S(_05904_),
    .X(_05919_));
 sky130_fd_sc_hd__mux4_1 _12741_ (.A0(_04029_),
    .A1(_04507_),
    .A2(_04506_),
    .A3(_04513_),
    .S0(_05904_),
    .S1(net23),
    .X(_05920_));
 sky130_fd_sc_hd__mux2_1 _12742_ (.A0(_05919_),
    .A1(_05920_),
    .S(net25),
    .X(_05921_));
 sky130_fd_sc_hd__mux4_1 _12743_ (.A0(_04643_),
    .A1(_05105_),
    .A2(_04481_),
    .A3(_04032_),
    .S0(_05904_),
    .S1(net23),
    .X(_05922_));
 sky130_fd_sc_hd__or2_1 _12744_ (.A(net24),
    .B(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__a22o_1 _12745_ (.A1(net24),
    .A2(_05906_),
    .B1(_05912_),
    .B2(net26),
    .X(_05924_));
 sky130_fd_sc_hd__o2111a_1 _12746_ (.A1(_05893_),
    .A2(_05921_),
    .B1(_05923_),
    .C1(_05924_),
    .D1(net27),
    .X(_05925_));
 sky130_fd_sc_hd__and2_1 _12747_ (.A(net53),
    .B(_05890_),
    .X(_05926_));
 sky130_fd_sc_hd__a221o_1 _12748_ (.A1(net56),
    .A2(_05900_),
    .B1(_05896_),
    .B2(net54),
    .C1(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__o211a_1 _12749_ (.A1(net48),
    .A2(_05895_),
    .B1(_05891_),
    .C1(_05899_),
    .X(_05928_));
 sky130_fd_sc_hd__a32o_2 _12750_ (.A1(clknet_1_0__leaf__05825_),
    .A2(_05900_),
    .A3(_05891_),
    .B1(_05898_),
    .B2(\gpout3.clk_div[1] ),
    .X(_05929_));
 sky130_fd_sc_hd__a211o_2 _12751_ (.A1(_05894_),
    .A2(_05927_),
    .B1(_05928_),
    .C1(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__nor2_1 _12752_ (.A(_05899_),
    .B(_05895_),
    .Y(_05931_));
 sky130_fd_sc_hd__a41o_1 _12753_ (.A1(_05734_),
    .A2(_05931_),
    .A3(_05889_),
    .A4(_05894_),
    .B1(_05903_),
    .X(_05932_));
 sky130_fd_sc_hd__a21o_1 _12754_ (.A1(net55),
    .A2(_05889_),
    .B1(net51),
    .X(_05933_));
 sky130_fd_sc_hd__a22o_1 _12755_ (.A1(_05931_),
    .A2(_05933_),
    .B1(_05900_),
    .B2(net50),
    .X(_05934_));
 sky130_fd_sc_hd__a22o_1 _12756_ (.A1(net46),
    .A2(_05896_),
    .B1(_05890_),
    .B2(net43),
    .X(_05935_));
 sky130_fd_sc_hd__a22o_1 _12757_ (.A1(net40),
    .A2(_05896_),
    .B1(_05890_),
    .B2(net52),
    .X(_05936_));
 sky130_fd_sc_hd__a221o_1 _12758_ (.A1(_05319_),
    .A2(_05931_),
    .B1(_05900_),
    .B2(net41),
    .C1(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__mux2_1 _12759_ (.A0(_05935_),
    .A1(_05937_),
    .S(net25),
    .X(_05938_));
 sky130_fd_sc_hd__a22o_1 _12760_ (.A1(_05934_),
    .A2(_05894_),
    .B1(_05938_),
    .B2(_05893_),
    .X(_05939_));
 sky130_fd_sc_hd__a22o_2 _12761_ (.A1(_05889_),
    .A2(_05930_),
    .B1(_05932_),
    .B2(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__a211o_2 _12762_ (.A1(_05913_),
    .A2(_05918_),
    .B1(_05925_),
    .C1(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__o2bb2a_2 _12763_ (.A1_N(_05363_),
    .A2_N(_05892_),
    .B1(_05911_),
    .B2(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__mux2_2 _12764_ (.A0(\reg_gpout[3] ),
    .A1(clknet_1_0__leaf__05942_),
    .S(net45),
    .X(_05943_));
 sky130_fd_sc_hd__buf_1 _12765_ (.A(_05943_),
    .X(net60));
 sky130_fd_sc_hd__buf_2 _12766_ (.A(net29),
    .X(_05944_));
 sky130_fd_sc_hd__inv_2 _12767_ (.A(net33),
    .Y(_05945_));
 sky130_fd_sc_hd__clkbuf_4 _12768_ (.A(net28),
    .X(_05946_));
 sky130_fd_sc_hd__or2_1 _12769_ (.A(_05946_),
    .B(_05102_),
    .X(_05947_));
 sky130_fd_sc_hd__inv_2 _12770_ (.A(net31),
    .Y(_05948_));
 sky130_fd_sc_hd__nor2_1 _12771_ (.A(_05948_),
    .B(net32),
    .Y(_05949_));
 sky130_fd_sc_hd__nand2_1 _12772_ (.A(_05946_),
    .B(_05363_),
    .Y(_05950_));
 sky130_fd_sc_hd__mux4_1 _12773_ (.A0(_05450_),
    .A1(_05539_),
    .A2(_05629_),
    .A3(_05710_),
    .S0(_05946_),
    .S1(net31),
    .X(_05951_));
 sky130_fd_sc_hd__a32o_1 _12774_ (.A1(_05947_),
    .A2(_05949_),
    .A3(_05950_),
    .B1(_05951_),
    .B2(net32),
    .X(_05952_));
 sky130_fd_sc_hd__and4_1 _12775_ (.A(_05944_),
    .B(net30),
    .C(_05945_),
    .D(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__inv_2 _12776_ (.A(net32),
    .Y(_05954_));
 sky130_fd_sc_hd__nor2_1 _12777_ (.A(_05944_),
    .B(_05946_),
    .Y(_05955_));
 sky130_fd_sc_hd__and2b_1 _12778_ (.A_N(_05944_),
    .B(net28),
    .X(_05956_));
 sky130_fd_sc_hd__a22o_1 _12779_ (.A1(_05100_),
    .A2(_05955_),
    .B1(_05956_),
    .B2(net72),
    .X(_05957_));
 sky130_fd_sc_hd__and2b_1 _12780_ (.A_N(net28),
    .B(net29),
    .X(_05958_));
 sky130_fd_sc_hd__nor2_2 _12781_ (.A(net31),
    .B(net30),
    .Y(_05959_));
 sky130_fd_sc_hd__and4_1 _12782_ (.A(_05944_),
    .B(_05946_),
    .C(_05098_),
    .D(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__a31o_1 _12783_ (.A1(net44),
    .A2(_05958_),
    .A3(_05959_),
    .B1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__a31o_1 _12784_ (.A1(_05948_),
    .A2(net30),
    .A3(_05957_),
    .B1(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__a21oi_1 _12785_ (.A1(_05944_),
    .A2(net30),
    .B1(net31),
    .Y(_05963_));
 sky130_fd_sc_hd__mux2_1 _12786_ (.A0(_05752_),
    .A1(_04723_),
    .S(_05946_),
    .X(_05964_));
 sky130_fd_sc_hd__mux2_1 _12787_ (.A0(_04718_),
    .A1(_04714_),
    .S(net28),
    .X(_05965_));
 sky130_fd_sc_hd__mux2_1 _12788_ (.A0(_04701_),
    .A1(_04704_),
    .S(net28),
    .X(_05966_));
 sky130_fd_sc_hd__mux4_1 _12789_ (.A0(_05760_),
    .A1(_04744_),
    .A2(_05761_),
    .A3(_05762_),
    .S0(net28),
    .S1(net31),
    .X(_05967_));
 sky130_fd_sc_hd__mux4_1 _12790_ (.A0(_05964_),
    .A1(_05965_),
    .A2(_05966_),
    .A3(_05967_),
    .S0(net30),
    .S1(_05944_),
    .X(_05968_));
 sky130_fd_sc_hd__and4b_1 _12791_ (.A_N(_05963_),
    .B(_05968_),
    .C(net32),
    .D(net33),
    .X(_05969_));
 sky130_fd_sc_hd__mux4_1 _12792_ (.A0(_04643_),
    .A1(_05105_),
    .A2(_04481_),
    .A3(_04032_),
    .S0(_05946_),
    .S1(_05944_),
    .X(_05970_));
 sky130_fd_sc_hd__mux2_1 _12793_ (.A0(_04033_),
    .A1(_04034_),
    .S(net28),
    .X(_05971_));
 sky130_fd_sc_hd__mux4_1 _12794_ (.A0(\gpout0.hpos[0] ),
    .A1(_04507_),
    .A2(\gpout0.hpos[2] ),
    .A3(_04513_),
    .S0(net28),
    .S1(net29),
    .X(_05972_));
 sky130_fd_sc_hd__mux2_1 _12795_ (.A0(_05971_),
    .A1(_05972_),
    .S(net31),
    .X(_05973_));
 sky130_fd_sc_hd__or2b_1 _12796_ (.A(_05973_),
    .B_N(net30),
    .X(_05974_));
 sky130_fd_sc_hd__a22o_1 _12797_ (.A1(net30),
    .A2(_05949_),
    .B1(_05963_),
    .B2(net32),
    .X(_05975_));
 sky130_fd_sc_hd__o2111a_1 _12798_ (.A1(net30),
    .A2(_05970_),
    .B1(_05974_),
    .C1(net33),
    .D1(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__nand2_1 _12799_ (.A(_05944_),
    .B(_05946_),
    .Y(_05977_));
 sky130_fd_sc_hd__nor2_1 _12800_ (.A(net32),
    .B(net33),
    .Y(_05978_));
 sky130_fd_sc_hd__nand2_1 _12801_ (.A(_05734_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(_05948_),
    .B(net30),
    .Y(_05980_));
 sky130_fd_sc_hd__o32a_1 _12803_ (.A1(_05977_),
    .A2(_05979_),
    .A3(_05980_),
    .B1(_05945_),
    .B2(net32),
    .X(_05981_));
 sky130_fd_sc_hd__a21oi_1 _12804_ (.A1(net55),
    .A2(_05978_),
    .B1(net51),
    .Y(_05982_));
 sky130_fd_sc_hd__o2bb2a_1 _12805_ (.A1_N(net50),
    .A2_N(_05958_),
    .B1(_05977_),
    .B2(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__mux4_1 _12806_ (.A0(net52),
    .A1(net41),
    .A2(net40),
    .A3(_05319_),
    .S0(_05944_),
    .S1(_05946_),
    .X(_05984_));
 sky130_fd_sc_hd__a221o_1 _12807_ (.A1(net43),
    .A2(_05955_),
    .B1(_05956_),
    .B2(net46),
    .C1(net31),
    .X(_05985_));
 sky130_fd_sc_hd__o21ai_1 _12808_ (.A1(_05948_),
    .A2(_05984_),
    .B1(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__o22a_1 _12809_ (.A1(_05983_),
    .A2(_05980_),
    .B1(_05986_),
    .B2(net30),
    .X(_05987_));
 sky130_fd_sc_hd__nor2_1 _12810_ (.A(_05981_),
    .B(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__a22o_1 _12811_ (.A1(net56),
    .A2(_05958_),
    .B1(_05956_),
    .B2(net54),
    .X(_05989_));
 sky130_fd_sc_hd__a21oi_1 _12812_ (.A1(net53),
    .A2(_05955_),
    .B1(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__nor2_1 _12813_ (.A(_05980_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__nand2_1 _12814_ (.A(_05955_),
    .B(_05959_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand3_1 _12815_ (.A(net3),
    .B(_05956_),
    .C(_05959_),
    .Y(_05993_));
 sky130_fd_sc_hd__nand2_1 _12816_ (.A(_05992_),
    .B(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__and4_1 _12817_ (.A(_05944_),
    .B(_05946_),
    .C(\gpout4.clk_div[1] ),
    .D(_05959_),
    .X(_05995_));
 sky130_fd_sc_hd__a31o_2 _12818_ (.A1(clknet_1_0__leaf__05825_),
    .A2(_05958_),
    .A3(_05959_),
    .B1(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__o31a_2 _12819_ (.A1(_05991_),
    .A2(_05994_),
    .A3(_05996_),
    .B1(_05978_),
    .X(_05997_));
 sky130_fd_sc_hd__or4_2 _12820_ (.A(_05969_),
    .B(_05976_),
    .C(_05988_),
    .D(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__a31o_2 _12821_ (.A1(_05954_),
    .A2(net33),
    .A3(_05962_),
    .B1(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__or3b_1 _12822_ (.A(_05992_),
    .B(_05629_),
    .C_N(_05978_),
    .X(_06000_));
 sky130_fd_sc_hd__o21a_2 _12823_ (.A1(_05953_),
    .A2(_05999_),
    .B1(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__mux2_2 _12824_ (.A0(\reg_gpout[4] ),
    .A1(clknet_1_1__leaf__06001_),
    .S(net45),
    .X(_06002_));
 sky130_fd_sc_hd__buf_1 _12825_ (.A(_06002_),
    .X(net61));
 sky130_fd_sc_hd__or2_1 _12826_ (.A(net38),
    .B(net39),
    .X(_06003_));
 sky130_fd_sc_hd__clkbuf_4 _12827_ (.A(net34),
    .X(_06004_));
 sky130_fd_sc_hd__nor2_1 _12828_ (.A(net35),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__or4b_1 _12829_ (.A(net37),
    .B(net36),
    .C(_05710_),
    .D_N(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__inv_2 _12830_ (.A(net35),
    .Y(_06007_));
 sky130_fd_sc_hd__clkinv_2 _12831_ (.A(net36),
    .Y(_06008_));
 sky130_fd_sc_hd__or2_1 _12832_ (.A(_06004_),
    .B(_05102_),
    .X(_06009_));
 sky130_fd_sc_hd__nand2_1 _12833_ (.A(_06004_),
    .B(_05363_),
    .Y(_06010_));
 sky130_fd_sc_hd__inv_2 _12834_ (.A(net37),
    .Y(_06011_));
 sky130_fd_sc_hd__nor2_1 _12835_ (.A(_06011_),
    .B(net38),
    .Y(_06012_));
 sky130_fd_sc_hd__mux4_1 _12836_ (.A0(_05450_),
    .A1(_05539_),
    .A2(_05629_),
    .A3(_05710_),
    .S0(_06004_),
    .S1(net37),
    .X(_06013_));
 sky130_fd_sc_hd__a32o_1 _12837_ (.A1(_06009_),
    .A2(_06010_),
    .A3(_06012_),
    .B1(_06013_),
    .B2(net38),
    .X(_06014_));
 sky130_fd_sc_hd__or3b_1 _12838_ (.A(_06007_),
    .B(_06008_),
    .C_N(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__mux4_1 _12839_ (.A0(_05752_),
    .A1(_05753_),
    .A2(_05755_),
    .A3(_05756_),
    .S0(_06004_),
    .S1(net36),
    .X(_06016_));
 sky130_fd_sc_hd__mux4_1 _12840_ (.A0(_05758_),
    .A1(_04704_),
    .A2(_05761_),
    .A3(_05762_),
    .S0(_06004_),
    .S1(net36),
    .X(_06017_));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(_06016_),
    .A1(_06017_),
    .S(net35),
    .X(_06018_));
 sky130_fd_sc_hd__mux4_1 _12842_ (.A0(_04643_),
    .A1(_04033_),
    .A2(_05105_),
    .A3(_04034_),
    .S0(net36),
    .S1(_06004_),
    .X(_06019_));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(_04481_),
    .A1(_04032_),
    .S(_06004_),
    .X(_06020_));
 sky130_fd_sc_hd__mux2_1 _12844_ (.A0(_05760_),
    .A1(_04744_),
    .S(net34),
    .X(_06021_));
 sky130_fd_sc_hd__and3_1 _12845_ (.A(net35),
    .B(net36),
    .C(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__a31o_1 _12846_ (.A1(net35),
    .A2(_06008_),
    .A3(_06020_),
    .B1(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__a211o_1 _12847_ (.A1(_06007_),
    .A2(_06019_),
    .B1(_06023_),
    .C1(net37),
    .X(_06024_));
 sky130_fd_sc_hd__o21ai_1 _12848_ (.A1(_06011_),
    .A2(_06018_),
    .B1(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__a211o_1 _12849_ (.A1(net43),
    .A2(_06005_),
    .B1(net36),
    .C1(net37),
    .X(_06026_));
 sky130_fd_sc_hd__and2_1 _12850_ (.A(net35),
    .B(net34),
    .X(_06027_));
 sky130_fd_sc_hd__and2_1 _12851_ (.A(_06007_),
    .B(net34),
    .X(_06028_));
 sky130_fd_sc_hd__nor2_1 _12852_ (.A(_06007_),
    .B(net34),
    .Y(_06029_));
 sky130_fd_sc_hd__a22o_1 _12853_ (.A1(net46),
    .A2(_06028_),
    .B1(_06029_),
    .B2(net44),
    .X(_06030_));
 sky130_fd_sc_hd__a21o_1 _12854_ (.A1(_05098_),
    .A2(_06027_),
    .B1(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__a22o_1 _12855_ (.A1(net40),
    .A2(_06028_),
    .B1(_06005_),
    .B2(net52),
    .X(_06032_));
 sky130_fd_sc_hd__a21o_1 _12856_ (.A1(_06008_),
    .A2(_06032_),
    .B1(_06011_),
    .X(_06033_));
 sky130_fd_sc_hd__a221o_1 _12857_ (.A1(net50),
    .A2(_06029_),
    .B1(_06027_),
    .B2(net51),
    .C1(_06008_),
    .X(_06034_));
 sky130_fd_sc_hd__a221o_1 _12858_ (.A1(net72),
    .A2(_06028_),
    .B1(_06005_),
    .B2(_05100_),
    .C1(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__o211a_1 _12859_ (.A1(_06026_),
    .A2(_06031_),
    .B1(_06033_),
    .C1(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__mux4_1 _12860_ (.A0(\gpout0.hpos[0] ),
    .A1(_04507_),
    .A2(_04506_),
    .A3(_04513_),
    .S0(_06004_),
    .S1(net35),
    .X(_06037_));
 sky130_fd_sc_hd__a221o_1 _12861_ (.A1(net41),
    .A2(_06029_),
    .B1(_06027_),
    .B2(_05319_),
    .C1(net36),
    .X(_06038_));
 sky130_fd_sc_hd__o211a_1 _12862_ (.A1(_06008_),
    .A2(_06037_),
    .B1(_06038_),
    .C1(net37),
    .X(_06039_));
 sky130_fd_sc_hd__o31a_1 _12863_ (.A1(net38),
    .A2(_06036_),
    .A3(_06039_),
    .B1(net39),
    .X(_06040_));
 sky130_fd_sc_hd__a21bo_1 _12864_ (.A1(net38),
    .A2(_06025_),
    .B1_N(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__nand2_1 _12865_ (.A(net54),
    .B(_06028_),
    .Y(_06042_));
 sky130_fd_sc_hd__a22o_1 _12866_ (.A1(net53),
    .A2(_06005_),
    .B1(_06029_),
    .B2(net56),
    .X(_06043_));
 sky130_fd_sc_hd__a21oi_1 _12867_ (.A1(_05734_),
    .A2(_06027_),
    .B1(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__a21o_2 _12868_ (.A1(net127),
    .A2(net35),
    .B1(_06004_),
    .X(_06045_));
 sky130_fd_sc_hd__nand2_1 _12869_ (.A(\gpout5.clk_div[1] ),
    .B(_06027_),
    .Y(_06046_));
 sky130_fd_sc_hd__a311o_2 _12870_ (.A1(_06008_),
    .A2(_06045_),
    .A3(_06046_),
    .B1(_06003_),
    .C1(net37),
    .X(_06047_));
 sky130_fd_sc_hd__a31o_2 _12871_ (.A1(net36),
    .A2(_06042_),
    .A3(_06044_),
    .B1(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__o211a_2 _12872_ (.A1(net39),
    .A2(_06015_),
    .B1(_06041_),
    .C1(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__o21ba_2 _12873_ (.A1(_06003_),
    .A2(_06006_),
    .B1_N(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__mux2_2 _12874_ (.A0(\reg_gpout[5] ),
    .A1(clknet_1_1__leaf__06050_),
    .S(net45),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _12875_ (.A(_06051_),
    .X(net62));
 sky130_fd_sc_hd__clkinv_2 _12876_ (.A(\rbzero.map_rom.i_row[4] ),
    .Y(_06052_));
 sky130_fd_sc_hd__inv_2 _12877_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .Y(_06053_));
 sky130_fd_sc_hd__nand2_1 _12878_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_06054_));
 sky130_fd_sc_hd__or2_1 _12879_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_06055_));
 sky130_fd_sc_hd__nand2_1 _12880_ (.A(_06054_),
    .B(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__nand2_2 _12881_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06057_));
 sky130_fd_sc_hd__or2_1 _12882_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_06058_));
 sky130_fd_sc_hd__nand2_1 _12883_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__nor2_1 _12884_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06060_));
 sky130_fd_sc_hd__and2_1 _12885_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_06061_));
 sky130_fd_sc_hd__nor2_1 _12886_ (.A(_06060_),
    .B(_06061_),
    .Y(_06062_));
 sky130_fd_sc_hd__or3b_1 _12887_ (.A(_06056_),
    .B(_06059_),
    .C_N(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__or2_1 _12888_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06064_));
 sky130_fd_sc_hd__xor2_2 _12889_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06065_));
 sky130_fd_sc_hd__and2_1 _12890_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06066_));
 sky130_fd_sc_hd__a31o_1 _12891_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_06065_),
    .B1(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__and2_1 _12892_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06068_));
 sky130_fd_sc_hd__a221o_1 _12893_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_06064_),
    .B2(_06067_),
    .C1(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__or2_2 _12894_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_06070_));
 sky130_fd_sc_hd__nand2_1 _12895_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_06071_));
 sky130_fd_sc_hd__or2_1 _12896_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_06072_));
 sky130_fd_sc_hd__and2_1 _12897_ (.A(_06071_),
    .B(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__nand4b_2 _12898_ (.A_N(_06063_),
    .B(_06069_),
    .C(_06070_),
    .D(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__nor2_1 _12899_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_06075_));
 sky130_fd_sc_hd__nand2_1 _12900_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06076_));
 sky130_fd_sc_hd__a2111o_1 _12901_ (.A1(_06071_),
    .A2(_06076_),
    .B1(_06060_),
    .C1(_06059_),
    .D1(_06056_),
    .X(_06077_));
 sky130_fd_sc_hd__o211a_1 _12902_ (.A1(_06075_),
    .A2(_06057_),
    .B1(_06077_),
    .C1(_06054_),
    .X(_06078_));
 sky130_fd_sc_hd__and2_1 _12903_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_06079_));
 sky130_fd_sc_hd__nor2_1 _12904_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_06080_));
 sky130_fd_sc_hd__or2_1 _12905_ (.A(_06079_),
    .B(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__a21oi_2 _12906_ (.A1(_06074_),
    .A2(_06078_),
    .B1(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand2_1 _12907_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_06083_));
 sky130_fd_sc_hd__or2b_1 _12908_ (.A(_06079_),
    .B_N(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__or2_1 _12909_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_06085_));
 sky130_fd_sc_hd__o221a_1 _12910_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(\rbzero.wall_tracer.rayAddendY[9] ),
    .B1(_06082_),
    .B2(_06084_),
    .C1(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__or2_1 _12911_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_06087_));
 sky130_fd_sc_hd__nand2_1 _12912_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06088_));
 sky130_fd_sc_hd__nand2_1 _12913_ (.A(_06087_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__nand2_1 _12914_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_06090_));
 sky130_fd_sc_hd__o21a_1 _12915_ (.A1(_06086_),
    .A2(_06089_),
    .B1(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__nand3_1 _12916_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .C(_06085_),
    .Y(_06092_));
 sky130_fd_sc_hd__nand2_1 _12917_ (.A(_06085_),
    .B(_06083_),
    .Y(_06093_));
 sky130_fd_sc_hd__a211o_1 _12918_ (.A1(_06074_),
    .A2(_06078_),
    .B1(_06093_),
    .C1(_06081_),
    .X(_06094_));
 sky130_fd_sc_hd__nor2_1 _12919_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06095_));
 sky130_fd_sc_hd__a41o_1 _12920_ (.A1(_06083_),
    .A2(_06092_),
    .A3(_06094_),
    .A4(_06088_),
    .B1(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__nand2_1 _12921_ (.A(_06087_),
    .B(_06090_),
    .Y(_06097_));
 sky130_fd_sc_hd__xor2_2 _12922_ (.A(_06096_),
    .B(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__and2b_1 _12923_ (.A_N(_06095_),
    .B(_06088_),
    .X(_06099_));
 sky130_fd_sc_hd__nand2_1 _12924_ (.A(_06083_),
    .B(_06092_),
    .Y(_06100_));
 sky130_fd_sc_hd__or3b_1 _12925_ (.A(_06099_),
    .B(_06100_),
    .C_N(_06094_),
    .X(_06101_));
 sky130_fd_sc_hd__o211ai_1 _12926_ (.A1(_06082_),
    .A2(_06084_),
    .B1(_06099_),
    .C1(_06085_),
    .Y(_06102_));
 sky130_fd_sc_hd__and2_1 _12927_ (.A(_06101_),
    .B(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__o21bai_1 _12928_ (.A1(_06079_),
    .A2(_06082_),
    .B1_N(_06093_),
    .Y(_06104_));
 sky130_fd_sc_hd__or3b_1 _12929_ (.A(_06079_),
    .B(_06082_),
    .C_N(_06093_),
    .X(_06105_));
 sky130_fd_sc_hd__and2_1 _12930_ (.A(_06104_),
    .B(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__nand3_1 _12931_ (.A(_06070_),
    .B(_06069_),
    .C(_06073_),
    .Y(_06107_));
 sky130_fd_sc_hd__a311o_2 _12932_ (.A1(_06071_),
    .A2(_06107_),
    .A3(_06076_),
    .B1(_06060_),
    .C1(_06059_),
    .X(_06108_));
 sky130_fd_sc_hd__inv_2 _12933_ (.A(_06060_),
    .Y(_06109_));
 sky130_fd_sc_hd__a32o_1 _12934_ (.A1(_06070_),
    .A2(_06069_),
    .A3(_06073_),
    .B1(\rbzero.wall_tracer.rayAddendY[3] ),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .X(_06110_));
 sky130_fd_sc_hd__a221o_1 _12935_ (.A1(_06057_),
    .A2(_06058_),
    .B1(_06109_),
    .B2(_06110_),
    .C1(_06061_),
    .X(_06111_));
 sky130_fd_sc_hd__and2_1 _12936_ (.A(_06108_),
    .B(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__and3_1 _12937_ (.A(_06081_),
    .B(_06074_),
    .C(_06078_),
    .X(_06113_));
 sky130_fd_sc_hd__nor2_1 _12938_ (.A(_06082_),
    .B(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__xor2_2 _12939_ (.A(_06062_),
    .B(_06110_),
    .X(_06115_));
 sky130_fd_sc_hd__a21o_1 _12940_ (.A1(_06070_),
    .A2(_06069_),
    .B1(_06073_),
    .X(_06116_));
 sky130_fd_sc_hd__and2_1 _12941_ (.A(_06107_),
    .B(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__nand2_1 _12942_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_06118_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(_06070_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__a21o_1 _12944_ (.A1(_06064_),
    .A2(_06067_),
    .B1(_06068_),
    .X(_06120_));
 sky130_fd_sc_hd__xnor2_2 _12945_ (.A(_06119_),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__or2b_1 _12946_ (.A(_06068_),
    .B_N(_06064_),
    .X(_06122_));
 sky130_fd_sc_hd__xnor2_2 _12947_ (.A(_06122_),
    .B(_06067_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _12948_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_06124_));
 sky130_fd_sc_hd__xnor2_2 _12949_ (.A(_06124_),
    .B(_06065_),
    .Y(_06125_));
 sky130_fd_sc_hd__xor2_2 _12950_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_06126_));
 sky130_fd_sc_hd__or4_1 _12951_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C(_06125_),
    .D(_06126_),
    .X(_06127_));
 sky130_fd_sc_hd__or4_1 _12952_ (.A(_06117_),
    .B(_06121_),
    .C(_06123_),
    .D(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__or3_1 _12953_ (.A(_06114_),
    .B(_06115_),
    .C(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__or3_1 _12954_ (.A(_06106_),
    .B(_06112_),
    .C(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__a21oi_1 _12955_ (.A1(_06057_),
    .A2(_06108_),
    .B1(_06056_),
    .Y(_06131_));
 sky130_fd_sc_hd__and3_1 _12956_ (.A(_06056_),
    .B(_06057_),
    .C(_06108_),
    .X(_06132_));
 sky130_fd_sc_hd__nor2_1 _12957_ (.A(_06131_),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__or4_1 _12958_ (.A(_06098_),
    .B(_06103_),
    .C(_06130_),
    .D(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__and2_1 _12959_ (.A(_06091_),
    .B(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__clkbuf_4 _12960_ (.A(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__buf_4 _12961_ (.A(_06136_),
    .X(_06137_));
 sky130_fd_sc_hd__a21oi_2 _12962_ (.A1(_06052_),
    .A2(_06053_),
    .B1(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__xnor2_1 _12963_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .B(_06137_),
    .Y(_06139_));
 sky130_fd_sc_hd__xnor2_1 _12964_ (.A(\rbzero.map_rom.i_row[4] ),
    .B(_06137_),
    .Y(_06140_));
 sky130_fd_sc_hd__inv_2 _12965_ (.A(\rbzero.map_rom.a6 ),
    .Y(_06141_));
 sky130_fd_sc_hd__nand2_1 _12966_ (.A(_06141_),
    .B(_06137_),
    .Y(_06142_));
 sky130_fd_sc_hd__clkinv_2 _12967_ (.A(\rbzero.map_rom.b6 ),
    .Y(_06143_));
 sky130_fd_sc_hd__clkinv_2 _12968_ (.A(\rbzero.map_rom.c6 ),
    .Y(_06144_));
 sky130_fd_sc_hd__nor2_1 _12969_ (.A(_06144_),
    .B(_06136_),
    .Y(_06145_));
 sky130_fd_sc_hd__nand2_1 _12970_ (.A(_06091_),
    .B(_06134_),
    .Y(_06146_));
 sky130_fd_sc_hd__clkbuf_4 _12971_ (.A(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__nor2_1 _12972_ (.A(\rbzero.map_rom.c6 ),
    .B(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__nor2_1 _12973_ (.A(_06145_),
    .B(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__and2_1 _12974_ (.A(\rbzero.map_rom.d6 ),
    .B(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__buf_2 _12975_ (.A(\rbzero.map_rom.b6 ),
    .X(_06151_));
 sky130_fd_sc_hd__xnor2_1 _12976_ (.A(_06151_),
    .B(_06137_),
    .Y(_06152_));
 sky130_fd_sc_hd__o21ai_1 _12977_ (.A1(_06145_),
    .A2(_06150_),
    .B1(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__o21ai_1 _12978_ (.A1(_06143_),
    .A2(_06137_),
    .B1(_06153_),
    .Y(_06154_));
 sky130_fd_sc_hd__nand2_1 _12979_ (.A(\rbzero.map_rom.a6 ),
    .B(_06147_),
    .Y(_06155_));
 sky130_fd_sc_hd__or2b_1 _12980_ (.A(_06154_),
    .B_N(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__and3_1 _12981_ (.A(_06140_),
    .B(_06142_),
    .C(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__and2_1 _12982_ (.A(_06139_),
    .B(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__xnor2_1 _12983_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_06137_),
    .Y(_06159_));
 sky130_fd_sc_hd__o21a_1 _12984_ (.A1(_06138_),
    .A2(_06158_),
    .B1(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__or3b_1 _12985_ (.A(_04486_),
    .B(_04487_),
    .C_N(\rbzero.trace_state[3] ),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_4 _12986_ (.A(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__buf_6 _12987_ (.A(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__buf_6 _12988_ (.A(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__inv_2 _12989_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .Y(_06165_));
 sky130_fd_sc_hd__nor2_1 _12990_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__inv_2 _12991_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .Y(_06167_));
 sky130_fd_sc_hd__inv_2 _12992_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .Y(_06168_));
 sky130_fd_sc_hd__o22a_1 _12993_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(_06167_),
    .B1(\rbzero.wall_tracer.trackDistX[-1] ),
    .B2(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__inv_2 _12994_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .Y(_06170_));
 sky130_fd_sc_hd__o2bb2a_1 _12995_ (.A1_N(\rbzero.wall_tracer.trackDistX[-1] ),
    .A2_N(_06168_),
    .B1(_06170_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_06171_));
 sky130_fd_sc_hd__nand2_1 _12996_ (.A(_06169_),
    .B(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__inv_2 _12997_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .Y(_06173_));
 sky130_fd_sc_hd__inv_2 _12998_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .Y(_06174_));
 sky130_fd_sc_hd__a22o_1 _12999_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_06173_),
    .B1(\rbzero.wall_tracer.trackDistX[2] ),
    .B2(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__inv_2 _13000_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .Y(_06176_));
 sky130_fd_sc_hd__a2bb2o_1 _13001_ (.A1_N(_06176_),
    .A2_N(\rbzero.wall_tracer.trackDistX[-3] ),
    .B1(_06170_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_06177_));
 sky130_fd_sc_hd__inv_2 _13002_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .Y(_06178_));
 sky130_fd_sc_hd__inv_2 _13003_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .Y(_06179_));
 sky130_fd_sc_hd__o22a_1 _13004_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(_06179_),
    .B1(\rbzero.wall_tracer.trackDistX[3] ),
    .B2(_06173_),
    .X(_06180_));
 sky130_fd_sc_hd__o221ai_1 _13005_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_06174_),
    .B1(_06178_),
    .B2(\rbzero.wall_tracer.trackDistX[1] ),
    .C1(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__and2_1 _13006_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(_06179_),
    .X(_06182_));
 sky130_fd_sc_hd__a22o_1 _13007_ (.A1(_06178_),
    .A2(\rbzero.wall_tracer.trackDistX[1] ),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_06167_),
    .X(_06183_));
 sky130_fd_sc_hd__a2111o_1 _13008_ (.A1(_06176_),
    .A2(\rbzero.wall_tracer.trackDistX[-3] ),
    .B1(_06181_),
    .C1(_06182_),
    .D1(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__or4_1 _13009_ (.A(_06172_),
    .B(_06175_),
    .C(_06177_),
    .D(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__inv_2 _13010_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .Y(_06186_));
 sky130_fd_sc_hd__nor2_1 _13011_ (.A(_06186_),
    .B(\rbzero.wall_tracer.trackDistY[9] ),
    .Y(_06187_));
 sky130_fd_sc_hd__inv_2 _13012_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .Y(_06188_));
 sky130_fd_sc_hd__nor2_1 _13013_ (.A(_06188_),
    .B(\rbzero.wall_tracer.trackDistY[-9] ),
    .Y(_06189_));
 sky130_fd_sc_hd__inv_2 _13014_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .Y(_06190_));
 sky130_fd_sc_hd__and2_1 _13015_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__or4_1 _13016_ (.A(_06166_),
    .B(_06187_),
    .C(_06189_),
    .D(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__a22o_1 _13017_ (.A1(\rbzero.wall_tracer.trackDistY[10] ),
    .A2(_06165_),
    .B1(_06186_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .X(_06193_));
 sky130_fd_sc_hd__inv_2 _13018_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .Y(_06194_));
 sky130_fd_sc_hd__o22a_1 _13019_ (.A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .A2(_06194_),
    .B1(\rbzero.wall_tracer.trackDistX[-5] ),
    .B2(_06190_),
    .X(_06195_));
 sky130_fd_sc_hd__inv_2 _13020_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .Y(_06196_));
 sky130_fd_sc_hd__inv_2 _13021_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .Y(_06197_));
 sky130_fd_sc_hd__o22a_1 _13022_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(_06196_),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .B2(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__a21bo_1 _13023_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(_06196_),
    .B1_N(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__inv_2 _13024_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .Y(_06200_));
 sky130_fd_sc_hd__nor2_1 _13025_ (.A(_06200_),
    .B(\rbzero.wall_tracer.trackDistY[-6] ),
    .Y(_06201_));
 sky130_fd_sc_hd__a221o_1 _13026_ (.A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .A2(_06194_),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .B2(_06197_),
    .C1(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__nor2_1 _13027_ (.A(_06199_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__or4bb_1 _13028_ (.A(_06192_),
    .B(_06193_),
    .C_N(_06195_),
    .D_N(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__inv_2 _13029_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .Y(_06205_));
 sky130_fd_sc_hd__inv_2 _13030_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .Y(_06206_));
 sky130_fd_sc_hd__a22o_1 _13031_ (.A1(_06205_),
    .A2(\rbzero.wall_tracer.trackDistY[6] ),
    .B1(\rbzero.wall_tracer.trackDistY[5] ),
    .B2(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__inv_2 _13032_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .Y(_06208_));
 sky130_fd_sc_hd__or2_1 _13033_ (.A(_06208_),
    .B(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_06209_));
 sky130_fd_sc_hd__o21ai_1 _13034_ (.A1(\rbzero.wall_tracer.trackDistY[5] ),
    .A2(_06206_),
    .B1(_06209_),
    .Y(_06210_));
 sky130_fd_sc_hd__inv_2 _13035_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .Y(_06211_));
 sky130_fd_sc_hd__a22o_1 _13036_ (.A1(_06208_),
    .A2(\rbzero.wall_tracer.trackDistY[8] ),
    .B1(_06211_),
    .B2(\rbzero.wall_tracer.trackDistY[7] ),
    .X(_06212_));
 sky130_fd_sc_hd__o22a_1 _13037_ (.A1(_06211_),
    .A2(\rbzero.wall_tracer.trackDistY[7] ),
    .B1(_06205_),
    .B2(\rbzero.wall_tracer.trackDistY[6] ),
    .X(_06213_));
 sky130_fd_sc_hd__or4b_1 _13038_ (.A(_06207_),
    .B(_06210_),
    .C(_06212_),
    .D_N(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__inv_2 _13039_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .Y(_06215_));
 sky130_fd_sc_hd__nor2_1 _13040_ (.A(_06215_),
    .B(\rbzero.wall_tracer.trackDistY[-8] ),
    .Y(_06216_));
 sky130_fd_sc_hd__inv_2 _13041_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .Y(_06217_));
 sky130_fd_sc_hd__nor2_1 _13042_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__a22o_1 _13043_ (.A1(_06200_),
    .A2(\rbzero.wall_tracer.trackDistY[-6] ),
    .B1(\rbzero.wall_tracer.trackDistY[-7] ),
    .B2(_06217_),
    .X(_06219_));
 sky130_fd_sc_hd__a22o_1 _13044_ (.A1(_06215_),
    .A2(\rbzero.wall_tracer.trackDistY[-8] ),
    .B1(_06188_),
    .B2(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(_06220_));
 sky130_fd_sc_hd__or4_1 _13045_ (.A(_06216_),
    .B(_06218_),
    .C(_06219_),
    .D(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__or3_1 _13046_ (.A(_06204_),
    .B(_06214_),
    .C(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__a21boi_1 _13047_ (.A1(_06171_),
    .A2(_06177_),
    .B1_N(_06169_),
    .Y(_06223_));
 sky130_fd_sc_hd__o21ba_1 _13048_ (.A1(_06183_),
    .A2(_06223_),
    .B1_N(_06181_),
    .X(_06224_));
 sky130_fd_sc_hd__a211o_1 _13049_ (.A1(_06175_),
    .A2(_06180_),
    .B1(_06182_),
    .C1(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__o21a_1 _13050_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(_06196_),
    .B1(_06199_),
    .X(_06226_));
 sky130_fd_sc_hd__o21ba_1 _13051_ (.A1(_06189_),
    .A2(_06226_),
    .B1_N(_06220_),
    .X(_06227_));
 sky130_fd_sc_hd__inv_2 _13052_ (.A(_06219_),
    .Y(_06228_));
 sky130_fd_sc_hd__o31a_1 _13053_ (.A1(_06216_),
    .A2(_06218_),
    .A3(_06227_),
    .B1(_06228_),
    .X(_06229_));
 sky130_fd_sc_hd__or3_1 _13054_ (.A(_06191_),
    .B(_06201_),
    .C(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__a221o_1 _13055_ (.A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .A2(_06194_),
    .B1(_06195_),
    .B2(_06230_),
    .C1(_06185_),
    .X(_06231_));
 sky130_fd_sc_hd__a21o_1 _13056_ (.A1(_06225_),
    .A2(_06231_),
    .B1(_06214_),
    .X(_06232_));
 sky130_fd_sc_hd__o221a_1 _13057_ (.A1(_06211_),
    .A2(\rbzero.wall_tracer.trackDistY[7] ),
    .B1(_06205_),
    .B2(\rbzero.wall_tracer.trackDistY[6] ),
    .C1(_06207_),
    .X(_06233_));
 sky130_fd_sc_hd__o21ai_1 _13058_ (.A1(_06212_),
    .A2(_06233_),
    .B1(_06209_),
    .Y(_06234_));
 sky130_fd_sc_hd__a21oi_1 _13059_ (.A1(_06232_),
    .A2(_06234_),
    .B1(_06187_),
    .Y(_06235_));
 sky130_fd_sc_hd__o22ai_2 _13060_ (.A1(_06185_),
    .A2(_06222_),
    .B1(_06235_),
    .B2(_06193_),
    .Y(_06236_));
 sky130_fd_sc_hd__nor2_2 _13061_ (.A(_06166_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__inv_2 _13062_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .Y(_06238_));
 sky130_fd_sc_hd__buf_2 _13063_ (.A(\rbzero.map_rom.f2 ),
    .X(_06239_));
 sky130_fd_sc_hd__inv_2 _13064_ (.A(_06239_),
    .Y(_06240_));
 sky130_fd_sc_hd__inv_2 _13065_ (.A(\rbzero.map_rom.i_col[4] ),
    .Y(_06241_));
 sky130_fd_sc_hd__o2bb2a_1 _13066_ (.A1_N(\rbzero.debug_overlay.playerX[2] ),
    .A2_N(_06240_),
    .B1(_06241_),
    .B2(\rbzero.debug_overlay.playerX[4] ),
    .X(_06242_));
 sky130_fd_sc_hd__o221a_1 _13067_ (.A1(_04734_),
    .A2(_06144_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(_06238_),
    .C1(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__clkinv_2 _13068_ (.A(\rbzero.map_rom.f4 ),
    .Y(_06244_));
 sky130_fd_sc_hd__inv_2 _13069_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .Y(_06245_));
 sky130_fd_sc_hd__o22a_1 _13070_ (.A1(_04735_),
    .A2(\rbzero.map_rom.f3 ),
    .B1(_06151_),
    .B2(_04736_),
    .X(_06246_));
 sky130_fd_sc_hd__o221a_1 _13071_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_06244_),
    .B1(\rbzero.wall_tracer.mapY[5] ),
    .B2(_06245_),
    .C1(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__inv_2 _13072_ (.A(\rbzero.map_rom.d6 ),
    .Y(_06248_));
 sky130_fd_sc_hd__o22a_1 _13073_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_06248_),
    .B1(_06052_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .X(_06249_));
 sky130_fd_sc_hd__o22a_1 _13074_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_06141_),
    .B1(_06053_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .X(_06250_));
 sky130_fd_sc_hd__o221a_1 _13075_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_06143_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_04725_),
    .C1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__o211a_1 _13076_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_06240_),
    .B1(_06249_),
    .C1(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__and3_1 _13077_ (.A(_06243_),
    .B(_06247_),
    .C(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__nand2_1 _13078_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(\rbzero.wall_tracer.mapX[5] ),
    .Y(_06254_));
 sky130_fd_sc_hd__or2_1 _13079_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(\rbzero.wall_tracer.mapX[5] ),
    .X(_06255_));
 sky130_fd_sc_hd__or4_1 _13080_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(\rbzero.wall_tracer.mapY[9] ),
    .C(\rbzero.wall_tracer.mapY[8] ),
    .D(\rbzero.wall_tracer.mapY[10] ),
    .X(_06256_));
 sky130_fd_sc_hd__or4_1 _13081_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(\rbzero.wall_tracer.mapX[8] ),
    .C(\rbzero.wall_tracer.mapX[10] ),
    .D(\rbzero.wall_tracer.mapY[7] ),
    .X(_06257_));
 sky130_fd_sc_hd__a211o_1 _13082_ (.A1(_06254_),
    .A2(_06255_),
    .B1(_06256_),
    .C1(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__clkbuf_4 _13083_ (.A(\rbzero.map_rom.f1 ),
    .X(_06259_));
 sky130_fd_sc_hd__a22o_1 _13084_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_06241_),
    .B1(_06248_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .X(_06260_));
 sky130_fd_sc_hd__a221o_1 _13085_ (.A1(_04730_),
    .A2(_06259_),
    .B1(_06144_),
    .B2(_04734_),
    .C1(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__buf_2 _13086_ (.A(\rbzero.map_rom.f3 ),
    .X(_06262_));
 sky130_fd_sc_hd__inv_2 _13087_ (.A(\rbzero.map_rom.f1 ),
    .Y(_06263_));
 sky130_fd_sc_hd__a211o_1 _13088_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_06244_),
    .B1(\rbzero.wall_tracer.mapX[7] ),
    .C1(\rbzero.wall_tracer.mapX[6] ),
    .X(_06264_));
 sky130_fd_sc_hd__a221o_1 _13089_ (.A1(_04735_),
    .A2(_06262_),
    .B1(_06263_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .C1(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__nor3_1 _13090_ (.A(_06258_),
    .B(_06261_),
    .C(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__or4_1 _13091_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(\rbzero.wall_tracer.visualWallDist[6] ),
    .C(\rbzero.wall_tracer.visualWallDist[5] ),
    .D(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_06267_));
 sky130_fd_sc_hd__or4_1 _13092_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(\rbzero.wall_tracer.visualWallDist[2] ),
    .C(\rbzero.wall_tracer.visualWallDist[1] ),
    .D(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_06268_));
 sky130_fd_sc_hd__or4_1 _13093_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(\rbzero.wall_tracer.visualWallDist[-2] ),
    .C(\rbzero.wall_tracer.visualWallDist[-3] ),
    .D(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__clkinv_4 _13094_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .Y(_06270_));
 sky130_fd_sc_hd__o41a_2 _13095_ (.A1(\rbzero.wall_tracer.visualWallDist[9] ),
    .A2(\rbzero.wall_tracer.visualWallDist[8] ),
    .A3(_06267_),
    .A4(_06269_),
    .B1(_06270_),
    .X(_06271_));
 sky130_fd_sc_hd__a21bo_1 _13096_ (.A1(_06253_),
    .A2(_06266_),
    .B1_N(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__xor2_1 _13097_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(_06151_),
    .X(_06273_));
 sky130_fd_sc_hd__a221o_1 _13098_ (.A1(\rbzero.map_overlay.i_mapdy[1] ),
    .A2(_06144_),
    .B1(_06052_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__xnor2_1 _13099_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_rom.a6 ),
    .Y(_06275_));
 sky130_fd_sc_hd__o221a_1 _13100_ (.A1(_04776_),
    .A2(\rbzero.map_rom.d6 ),
    .B1(_06052_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__o221a_1 _13101_ (.A1(\rbzero.map_overlay.i_mapdy[0] ),
    .A2(_06248_),
    .B1(_06144_),
    .B2(\rbzero.map_overlay.i_mapdy[1] ),
    .C1(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__or2_1 _13102_ (.A(\rbzero.map_rom.d6 ),
    .B(\rbzero.map_rom.c6 ),
    .X(_06278_));
 sky130_fd_sc_hd__or4_1 _13103_ (.A(_06151_),
    .B(\rbzero.map_rom.a6 ),
    .C(\rbzero.map_rom.i_row[4] ),
    .D(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__and4bb_2 _13104_ (.A_N(_06272_),
    .B_N(_06274_),
    .C(_06277_),
    .D(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__a22o_1 _13105_ (.A1(\rbzero.map_overlay.i_mapdx[2] ),
    .A2(_06240_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .B2(_04783_),
    .X(_06281_));
 sky130_fd_sc_hd__inv_2 _13106_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .Y(_06282_));
 sky130_fd_sc_hd__buf_2 _13107_ (.A(\rbzero.map_rom.f4 ),
    .X(_06283_));
 sky130_fd_sc_hd__nor2_1 _13108_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__and2_1 _13109_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06283_),
    .X(_06285_));
 sky130_fd_sc_hd__inv_2 _13110_ (.A(\rbzero.map_rom.f3 ),
    .Y(_06286_));
 sky130_fd_sc_hd__xnor2_1 _13111_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_06259_),
    .Y(_06287_));
 sky130_fd_sc_hd__o221a_1 _13112_ (.A1(\rbzero.map_overlay.i_mapdx[1] ),
    .A2(_06286_),
    .B1(_06240_),
    .B2(\rbzero.map_overlay.i_mapdx[2] ),
    .C1(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__o221a_1 _13113_ (.A1(_06282_),
    .A2(_06262_),
    .B1(_06284_),
    .B2(_06285_),
    .C1(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__a21o_1 _13114_ (.A1(_04783_),
    .A2(_04782_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .X(_06290_));
 sky130_fd_sc_hd__and4bb_4 _13115_ (.A_N(_06272_),
    .B_N(_06281_),
    .C(_06289_),
    .D(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__nand2_1 _13116_ (.A(\rbzero.map_rom.d6 ),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_1 _13117_ (.A(_06278_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__a22o_1 _13118_ (.A1(_06244_),
    .A2(_06248_),
    .B1(_06293_),
    .B2(_06262_),
    .X(_06294_));
 sky130_fd_sc_hd__and4_1 _13119_ (.A(_06283_),
    .B(_06262_),
    .C(_06239_),
    .D(\rbzero.map_rom.i_col[4] ),
    .X(_06295_));
 sky130_fd_sc_hd__a32o_1 _13120_ (.A1(_06239_),
    .A2(_06151_),
    .A3(_06294_),
    .B1(_06295_),
    .B2(_06259_),
    .X(_06296_));
 sky130_fd_sc_hd__or4_1 _13121_ (.A(_06283_),
    .B(_06262_),
    .C(_06239_),
    .D(\rbzero.map_rom.i_col[4] ),
    .X(_06297_));
 sky130_fd_sc_hd__a22o_1 _13122_ (.A1(_06244_),
    .A2(_06248_),
    .B1(\rbzero.map_rom.c6 ),
    .B2(\rbzero.map_rom.f3 ),
    .X(_06298_));
 sky130_fd_sc_hd__a22o_1 _13123_ (.A1(_06286_),
    .A2(_06144_),
    .B1(_06151_),
    .B2(_06239_),
    .X(_06299_));
 sky130_fd_sc_hd__a2111o_1 _13124_ (.A1(_06240_),
    .A2(_06143_),
    .B1(\rbzero.map_rom.a6 ),
    .C1(_06298_),
    .D1(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__a221o_1 _13125_ (.A1(_06283_),
    .A2(\rbzero.map_rom.d6 ),
    .B1(_06297_),
    .B2(_06300_),
    .C1(_06259_),
    .X(_06301_));
 sky130_fd_sc_hd__nand2_1 _13126_ (.A(_06151_),
    .B(\rbzero.map_rom.i_row[4] ),
    .Y(_06302_));
 sky130_fd_sc_hd__or4_1 _13127_ (.A(_06283_),
    .B(_06239_),
    .C(\rbzero.map_rom.d6 ),
    .D(_06151_),
    .X(_06303_));
 sky130_fd_sc_hd__o31a_1 _13128_ (.A1(_06141_),
    .A2(_06292_),
    .A3(_06302_),
    .B1(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__and4b_1 _13129_ (.A_N(_06296_),
    .B(_06301_),
    .C(_06279_),
    .D(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__nand2_1 _13130_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06306_));
 sky130_fd_sc_hd__or2_1 _13131_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(\rbzero.map_rom.c6 ),
    .X(_06307_));
 sky130_fd_sc_hd__or2_1 _13132_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .B(_06239_),
    .X(_06308_));
 sky130_fd_sc_hd__nand2_1 _13133_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .B(_06239_),
    .Y(_06309_));
 sky130_fd_sc_hd__xor2_1 _13134_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(_06283_),
    .X(_06310_));
 sky130_fd_sc_hd__a221o_1 _13135_ (.A1(_04792_),
    .A2(_06262_),
    .B1(_06143_),
    .B2(\rbzero.map_overlay.i_othery[2] ),
    .C1(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__a221o_1 _13136_ (.A1(_06306_),
    .A2(_06307_),
    .B1(_06308_),
    .B2(_06309_),
    .C1(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__o2bb2a_1 _13137_ (.A1_N(\rbzero.map_overlay.i_othery[0] ),
    .A2_N(_06248_),
    .B1(_06143_),
    .B2(\rbzero.map_overlay.i_othery[2] ),
    .X(_06313_));
 sky130_fd_sc_hd__o221a_1 _13138_ (.A1(_04793_),
    .A2(_06259_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_04791_),
    .C1(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__inv_2 _13139_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .Y(_06315_));
 sky130_fd_sc_hd__o22a_1 _13140_ (.A1(\rbzero.map_overlay.i_otherx[4] ),
    .A2(_06241_),
    .B1(_06141_),
    .B2(\rbzero.map_overlay.i_othery[3] ),
    .X(_06316_));
 sky130_fd_sc_hd__o221a_1 _13141_ (.A1(\rbzero.map_overlay.i_otherx[3] ),
    .A2(_06263_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .B2(_06315_),
    .C1(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__o22a_1 _13142_ (.A1(_04792_),
    .A2(_06262_),
    .B1(_06248_),
    .B2(\rbzero.map_overlay.i_othery[0] ),
    .X(_06318_));
 sky130_fd_sc_hd__o221a_1 _13143_ (.A1(_04797_),
    .A2(\rbzero.map_rom.a6 ),
    .B1(_06052_),
    .B2(\rbzero.map_overlay.i_othery[4] ),
    .C1(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__and3_1 _13144_ (.A(_06314_),
    .B(_06317_),
    .C(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__or2b_1 _13145_ (.A(_06312_),
    .B_N(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__a22o_1 _13146_ (.A1(_06259_),
    .A2(\rbzero.map_rom.c6 ),
    .B1(_06143_),
    .B2(_06244_),
    .X(_06322_));
 sky130_fd_sc_hd__a221o_1 _13147_ (.A1(_06286_),
    .A2(_06248_),
    .B1(_06144_),
    .B2(_06263_),
    .C1(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__xnor2_1 _13148_ (.A(_06239_),
    .B(\rbzero.map_rom.a6 ),
    .Y(_06324_));
 sky130_fd_sc_hd__a221o_1 _13149_ (.A1(_06262_),
    .A2(\rbzero.map_rom.d6 ),
    .B1(_06151_),
    .B2(_06283_),
    .C1(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__and4_1 _13150_ (.A(_06259_),
    .B(\rbzero.map_rom.c6 ),
    .C(\rbzero.map_rom.a6 ),
    .D(_06052_),
    .X(_06326_));
 sky130_fd_sc_hd__or4b_1 _13151_ (.A(_06262_),
    .B(\rbzero.map_rom.i_col[4] ),
    .C(_06303_),
    .D_N(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__o21a_1 _13152_ (.A1(_06323_),
    .A2(_06325_),
    .B1(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a31o_2 _13153_ (.A1(_06305_),
    .A2(_06321_),
    .A3(_06328_),
    .B1(_06272_),
    .X(_06329_));
 sky130_fd_sc_hd__or3b_4 _13154_ (.A(_06280_),
    .B(_06291_),
    .C_N(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__nor2_4 _13155_ (.A(_06162_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__nand2_2 _13156_ (.A(_06237_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__nor3_1 _13157_ (.A(_06162_),
    .B(_06280_),
    .C(_06291_),
    .Y(_06333_));
 sky130_fd_sc_hd__clkinv_2 _13158_ (.A(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__and2b_1 _13159_ (.A_N(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .X(_06335_));
 sky130_fd_sc_hd__nand2_2 _13160_ (.A(\rbzero.trace_state[1] ),
    .B(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__or2_1 _13161_ (.A(_04494_),
    .B(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__buf_4 _13162_ (.A(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__buf_8 _13163_ (.A(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__buf_8 _13164_ (.A(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__o21ai_2 _13165_ (.A1(_06334_),
    .A2(_06329_),
    .B1(_04490_),
    .Y(_06341_));
 sky130_fd_sc_hd__a21oi_1 _13166_ (.A1(_06334_),
    .A2(_06340_),
    .B1(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__nand2_2 _13167_ (.A(_06332_),
    .B(_06342_),
    .Y(_06343_));
 sky130_fd_sc_hd__nor2_2 _13168_ (.A(_06164_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__o31ai_1 _13169_ (.A1(_06159_),
    .A2(_06138_),
    .A3(_06158_),
    .B1(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__clkbuf_4 _13170_ (.A(_06343_),
    .X(_06346_));
 sky130_fd_sc_hd__a2bb2o_1 _13171_ (.A1_N(_06160_),
    .A2_N(_06345_),
    .B1(\rbzero.wall_tracer.mapY[6] ),
    .B2(_06346_),
    .X(_00386_));
 sky130_fd_sc_hd__xnor2_1 _13172_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .B(_06137_),
    .Y(_06347_));
 sky130_fd_sc_hd__a21oi_1 _13173_ (.A1(\rbzero.wall_tracer.mapY[6] ),
    .A2(_06147_),
    .B1(_06160_),
    .Y(_06348_));
 sky130_fd_sc_hd__xnor2_1 _13174_ (.A(_06347_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__a22o_1 _13175_ (.A1(\rbzero.wall_tracer.mapY[7] ),
    .A2(_06346_),
    .B1(_06344_),
    .B2(_06349_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _13176_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06147_),
    .X(_06350_));
 sky130_fd_sc_hd__nor2_1 _13177_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06147_),
    .Y(_06351_));
 sky130_fd_sc_hd__nor2_1 _13178_ (.A(_06350_),
    .B(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__o41a_1 _13179_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(\rbzero.wall_tracer.mapY[5] ),
    .A3(\rbzero.wall_tracer.mapY[7] ),
    .A4(\rbzero.wall_tracer.mapY[6] ),
    .B1(_06147_),
    .X(_06353_));
 sky130_fd_sc_hd__a31o_1 _13180_ (.A1(_06159_),
    .A2(_06158_),
    .A3(_06347_),
    .B1(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__xor2_1 _13181_ (.A(_06352_),
    .B(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__a22o_1 _13182_ (.A1(\rbzero.wall_tracer.mapY[8] ),
    .A2(_06346_),
    .B1(_06344_),
    .B2(_06355_),
    .X(_00388_));
 sky130_fd_sc_hd__a21o_1 _13183_ (.A1(_06352_),
    .A2(_06354_),
    .B1(_06350_),
    .X(_06356_));
 sky130_fd_sc_hd__xnor2_1 _13184_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(_06137_),
    .Y(_06357_));
 sky130_fd_sc_hd__nand2_1 _13185_ (.A(_06356_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__or2_1 _13186_ (.A(_06356_),
    .B(_06357_),
    .X(_06359_));
 sky130_fd_sc_hd__a32o_1 _13187_ (.A1(_06344_),
    .A2(_06358_),
    .A3(_06359_),
    .B1(_06346_),
    .B2(\rbzero.wall_tracer.mapY[9] ),
    .X(_00389_));
 sky130_fd_sc_hd__o21a_1 _13188_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06147_),
    .B1(_06356_),
    .X(_06360_));
 sky130_fd_sc_hd__a21o_1 _13189_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06147_),
    .B1(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__xnor2_1 _13190_ (.A(\rbzero.wall_tracer.mapY[10] ),
    .B(_06147_),
    .Y(_06362_));
 sky130_fd_sc_hd__xnor2_1 _13191_ (.A(_06361_),
    .B(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__a22o_1 _13192_ (.A1(\rbzero.wall_tracer.mapY[10] ),
    .A2(_06346_),
    .B1(_06344_),
    .B2(_06363_),
    .X(_00390_));
 sky130_fd_sc_hd__o211a_2 _13193_ (.A1(_06086_),
    .A2(_06089_),
    .B1(_04484_),
    .C1(_06090_),
    .X(_06364_));
 sky130_fd_sc_hd__nor2_1 _13194_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_04485_),
    .Y(_06365_));
 sky130_fd_sc_hd__inv_2 _13195_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06366_));
 sky130_fd_sc_hd__o21a_1 _13196_ (.A1(_06364_),
    .A2(_06365_),
    .B1(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nand2_1 _13197_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_06368_));
 sky130_fd_sc_hd__or2_1 _13198_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_06369_));
 sky130_fd_sc_hd__and2_1 _13199_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_06370_));
 sky130_fd_sc_hd__nor2_1 _13200_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_06371_));
 sky130_fd_sc_hd__nor2_1 _13201_ (.A(_06370_),
    .B(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__and2_1 _13202_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06373_));
 sky130_fd_sc_hd__nor2_1 _13203_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_06374_));
 sky130_fd_sc_hd__nor2_1 _13204_ (.A(_06373_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__xor2_1 _13205_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06376_));
 sky130_fd_sc_hd__o21a_1 _13206_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_06373_),
    .X(_06377_));
 sky130_fd_sc_hd__a21o_1 _13207_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__a21o_1 _13208_ (.A1(_06375_),
    .A2(_06376_),
    .B1(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__and2_1 _13209_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_06380_));
 sky130_fd_sc_hd__nor2_1 _13210_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_06381_));
 sky130_fd_sc_hd__nor2_1 _13211_ (.A(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__nor2_1 _13212_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06383_));
 sky130_fd_sc_hd__nor2_1 _13213_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06384_));
 sky130_fd_sc_hd__nand2_2 _13214_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_06385_));
 sky130_fd_sc_hd__nor2_1 _13215_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06386_));
 sky130_fd_sc_hd__nand2_1 _13216_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06387_));
 sky130_fd_sc_hd__nand2_1 _13217_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06388_));
 sky130_fd_sc_hd__o211a_1 _13218_ (.A1(_06385_),
    .A2(_06386_),
    .B1(_06387_),
    .C1(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nand2_1 _13219_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06390_));
 sky130_fd_sc_hd__o31ai_4 _13220_ (.A1(_06383_),
    .A2(_06384_),
    .A3(_06389_),
    .B1(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__xor2_1 _13221_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_06392_));
 sky130_fd_sc_hd__o21a_1 _13222_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[4] ),
    .B1(_06380_),
    .X(_06393_));
 sky130_fd_sc_hd__a21o_1 _13223_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[4] ),
    .B1(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__a311o_1 _13224_ (.A1(_06382_),
    .A2(_06391_),
    .A3(_06392_),
    .B1(_06394_),
    .C1(_06378_),
    .X(_06395_));
 sky130_fd_sc_hd__nand2_1 _13225_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_06396_));
 sky130_fd_sc_hd__or2b_1 _13226_ (.A(_06370_),
    .B_N(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__a31o_1 _13227_ (.A1(_06372_),
    .A2(_06379_),
    .A3(_06395_),
    .B1(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__or2_1 _13228_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_06399_));
 sky130_fd_sc_hd__and2_1 _13229_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_06400_));
 sky130_fd_sc_hd__a31o_1 _13230_ (.A1(_06369_),
    .A2(_06398_),
    .A3(_06399_),
    .B1(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__nor2_1 _13231_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_06402_));
 sky130_fd_sc_hd__a21o_1 _13232_ (.A1(_06368_),
    .A2(_06401_),
    .B1(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__a21oi_1 _13233_ (.A1(_04504_),
    .A2(_06403_),
    .B1(_06367_),
    .Y(_06404_));
 sky130_fd_sc_hd__nor2_2 _13234_ (.A(_04504_),
    .B(_06364_),
    .Y(_06405_));
 sky130_fd_sc_hd__or2_1 _13235_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_04485_),
    .X(_06406_));
 sky130_fd_sc_hd__nor2_2 _13236_ (.A(_06366_),
    .B(_06403_),
    .Y(_06407_));
 sky130_fd_sc_hd__a21o_1 _13237_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__inv_2 _13238_ (.A(_04484_),
    .Y(_06409_));
 sky130_fd_sc_hd__clkbuf_4 _13239_ (.A(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__a21o_1 _13240_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_06410_),
    .B1(_04503_),
    .X(_06411_));
 sky130_fd_sc_hd__a21o_1 _13241_ (.A1(_04485_),
    .A2(_06098_),
    .B1(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__and2b_1 _13242_ (.A_N(_06402_),
    .B(_06368_),
    .X(_06413_));
 sky130_fd_sc_hd__xnor2_2 _13243_ (.A(_06401_),
    .B(_06413_),
    .Y(_06414_));
 sky130_fd_sc_hd__nand2_1 _13244_ (.A(_04504_),
    .B(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__nand2_1 _13245_ (.A(_06369_),
    .B(_06398_),
    .Y(_06416_));
 sky130_fd_sc_hd__nand2_1 _13246_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_06417_));
 sky130_fd_sc_hd__nand2_1 _13247_ (.A(_06399_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__xnor2_2 _13248_ (.A(_06416_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__clkinv_4 _13249_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .Y(_06420_));
 sky130_fd_sc_hd__nor2_1 _13250_ (.A(_06420_),
    .B(_04484_),
    .Y(_06421_));
 sky130_fd_sc_hd__a311o_1 _13251_ (.A1(_04484_),
    .A2(_06101_),
    .A3(_06102_),
    .B1(_06421_),
    .C1(_04503_),
    .X(_06422_));
 sky130_fd_sc_hd__a21bo_1 _13252_ (.A1(_04504_),
    .A2(_06419_),
    .B1_N(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__a21bo_1 _13253_ (.A1(_06412_),
    .A2(_06415_),
    .B1_N(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__a31o_1 _13254_ (.A1(_06382_),
    .A2(_06391_),
    .A3(_06392_),
    .B1(_06394_),
    .X(_06425_));
 sky130_fd_sc_hd__a21o_1 _13255_ (.A1(_06375_),
    .A2(_06425_),
    .B1(_06373_),
    .X(_06426_));
 sky130_fd_sc_hd__xnor2_1 _13256_ (.A(_06376_),
    .B(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__and2_1 _13257_ (.A(_04503_),
    .B(_06427_),
    .X(_06428_));
 sky130_fd_sc_hd__a21oi_1 _13258_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_06410_),
    .B1(_04503_),
    .Y(_06429_));
 sky130_fd_sc_hd__o31a_1 _13259_ (.A1(_06410_),
    .A2(_06131_),
    .A3(_06132_),
    .B1(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__xnor2_1 _13260_ (.A(_06375_),
    .B(_06425_),
    .Y(_06431_));
 sky130_fd_sc_hd__a21o_1 _13261_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_06410_),
    .B1(_04502_),
    .X(_06432_));
 sky130_fd_sc_hd__a31o_1 _13262_ (.A1(_04484_),
    .A2(_06108_),
    .A3(_06111_),
    .B1(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__a21bo_1 _13263_ (.A1(_04503_),
    .A2(_06431_),
    .B1_N(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__a21o_1 _13264_ (.A1(_06382_),
    .A2(_06391_),
    .B1(_06380_),
    .X(_06435_));
 sky130_fd_sc_hd__xnor2_1 _13265_ (.A(_06392_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _13266_ (.A(_04484_),
    .B(_06115_),
    .Y(_06437_));
 sky130_fd_sc_hd__a21oi_1 _13267_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_06410_),
    .B1(_04503_),
    .Y(_06438_));
 sky130_fd_sc_hd__a22o_2 _13268_ (.A1(_04503_),
    .A2(_06436_),
    .B1(_06437_),
    .B2(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__xnor2_1 _13269_ (.A(_06382_),
    .B(_06391_),
    .Y(_06440_));
 sky130_fd_sc_hd__a21o_1 _13270_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_06409_),
    .B1(_04502_),
    .X(_06441_));
 sky130_fd_sc_hd__and3_1 _13271_ (.A(_04484_),
    .B(_06107_),
    .C(_06116_),
    .X(_06442_));
 sky130_fd_sc_hd__o2bb2a_2 _13272_ (.A1_N(_04502_),
    .A2_N(_06440_),
    .B1(_06441_),
    .B2(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__nor2_1 _13273_ (.A(_06410_),
    .B(_06121_),
    .Y(_06444_));
 sky130_fd_sc_hd__inv_2 _13274_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .Y(_06445_));
 sky130_fd_sc_hd__a21o_1 _13275_ (.A1(_06445_),
    .A2(_06409_),
    .B1(_04502_),
    .X(_06446_));
 sky130_fd_sc_hd__o21ai_1 _13276_ (.A1(_06385_),
    .A2(_06386_),
    .B1(_06387_),
    .Y(_06447_));
 sky130_fd_sc_hd__and2b_1 _13277_ (.A_N(_06384_),
    .B(_06388_),
    .X(_06448_));
 sky130_fd_sc_hd__xnor2_2 _13278_ (.A(_06447_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__nand2_1 _13279_ (.A(_04502_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__a21o_1 _13280_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_06409_),
    .B1(_04502_),
    .X(_06451_));
 sky130_fd_sc_hd__a21o_1 _13281_ (.A1(_04484_),
    .A2(_06123_),
    .B1(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__or2b_1 _13282_ (.A(_06386_),
    .B_N(_06387_),
    .X(_06453_));
 sky130_fd_sc_hd__xor2_4 _13283_ (.A(_06385_),
    .B(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__or2_1 _13284_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_04484_),
    .X(_06455_));
 sky130_fd_sc_hd__o211a_1 _13285_ (.A1(_06409_),
    .A2(_06125_),
    .B1(_06455_),
    .C1(_06366_),
    .X(_06456_));
 sky130_fd_sc_hd__mux2_1 _13286_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06457_));
 sky130_fd_sc_hd__mux2_2 _13287_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_06457_),
    .S(_06366_),
    .X(_06458_));
 sky130_fd_sc_hd__mux2_1 _13288_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06459_));
 sky130_fd_sc_hd__mux2_2 _13289_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_06459_),
    .S(_06366_),
    .X(_06460_));
 sky130_fd_sc_hd__or2_1 _13290_ (.A(_06458_),
    .B(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__or2_1 _13291_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_06462_));
 sky130_fd_sc_hd__and2_1 _13292_ (.A(_06385_),
    .B(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__mux2_1 _13293_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_06126_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06464_));
 sky130_fd_sc_hd__mux2_2 _13294_ (.A0(_06463_),
    .A1(_06464_),
    .S(_06366_),
    .X(_06465_));
 sky130_fd_sc_hd__a2111o_2 _13295_ (.A1(_04502_),
    .A2(_06454_),
    .B1(_06456_),
    .C1(_06461_),
    .D1(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__a21oi_1 _13296_ (.A1(_06450_),
    .A2(_06452_),
    .B1(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__nor2_1 _13297_ (.A(_06384_),
    .B(_06389_),
    .Y(_06468_));
 sky130_fd_sc_hd__or2b_1 _13298_ (.A(_06383_),
    .B_N(_06390_),
    .X(_06469_));
 sky130_fd_sc_hd__xnor2_2 _13299_ (.A(_06468_),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__nand2_1 _13300_ (.A(_04502_),
    .B(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__o211a_1 _13301_ (.A1(_06444_),
    .A2(_06446_),
    .B1(_06467_),
    .C1(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__and2b_1 _13302_ (.A_N(_06443_),
    .B(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__o2111a_1 _13303_ (.A1(_06428_),
    .A2(_06430_),
    .B1(_06434_),
    .C1(_06439_),
    .D1(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__nand2_1 _13304_ (.A(_06369_),
    .B(_06396_),
    .Y(_06475_));
 sky130_fd_sc_hd__a31o_1 _13305_ (.A1(_06372_),
    .A2(_06379_),
    .A3(_06395_),
    .B1(_06370_),
    .X(_06476_));
 sky130_fd_sc_hd__xor2_2 _13306_ (.A(_06475_),
    .B(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__nand2_1 _13307_ (.A(_04504_),
    .B(_06477_),
    .Y(_06478_));
 sky130_fd_sc_hd__a21o_1 _13308_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_06410_),
    .B1(_04503_),
    .X(_06479_));
 sky130_fd_sc_hd__a31o_1 _13309_ (.A1(_04485_),
    .A2(_06104_),
    .A3(_06105_),
    .B1(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__or3_1 _13310_ (.A(_06410_),
    .B(_06082_),
    .C(_06113_),
    .X(_06481_));
 sky130_fd_sc_hd__a21oi_1 _13311_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_06410_),
    .B1(_04502_),
    .Y(_06482_));
 sky130_fd_sc_hd__nand2_1 _13312_ (.A(_06379_),
    .B(_06395_),
    .Y(_06483_));
 sky130_fd_sc_hd__xor2_1 _13313_ (.A(_06372_),
    .B(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__a22o_2 _13314_ (.A1(_06481_),
    .A2(_06482_),
    .B1(_06484_),
    .B2(_04503_),
    .X(_06485_));
 sky130_fd_sc_hd__a21boi_1 _13315_ (.A1(_06478_),
    .A2(_06480_),
    .B1_N(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__nor2_1 _13316_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_04485_),
    .Y(_06487_));
 sky130_fd_sc_hd__a211o_2 _13317_ (.A1(_06368_),
    .A2(_06401_),
    .B1(_06366_),
    .C1(_06402_),
    .X(_06488_));
 sky130_fd_sc_hd__o31a_2 _13318_ (.A1(_04504_),
    .A2(_06364_),
    .A3(_06487_),
    .B1(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__nand3_1 _13319_ (.A(_06474_),
    .B(_06486_),
    .C(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__or2_1 _13320_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_04485_),
    .X(_06491_));
 sky130_fd_sc_hd__nor2_1 _13321_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_04485_),
    .Y(_06492_));
 sky130_fd_sc_hd__o31a_1 _13322_ (.A1(_04504_),
    .A2(_06364_),
    .A3(_06492_),
    .B1(_06488_),
    .X(_06493_));
 sky130_fd_sc_hd__a21bo_1 _13323_ (.A1(_06405_),
    .A2(_06491_),
    .B1_N(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__nor4_2 _13324_ (.A(_06408_),
    .B(_06424_),
    .C(_06490_),
    .D(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__o21a_1 _13325_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_04485_),
    .B1(_06405_),
    .X(_06496_));
 sky130_fd_sc_hd__or2_1 _13326_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_04485_),
    .X(_06497_));
 sky130_fd_sc_hd__a21oi_1 _13327_ (.A1(_06405_),
    .A2(_06497_),
    .B1(_06407_),
    .Y(_06498_));
 sky130_fd_sc_hd__and2b_1 _13328_ (.A_N(_06496_),
    .B(_06498_),
    .X(_06499_));
 sky130_fd_sc_hd__a211o_1 _13329_ (.A1(_06270_),
    .A2(_06410_),
    .B1(_04504_),
    .C1(_06364_),
    .X(_06500_));
 sky130_fd_sc_hd__and2_2 _13330_ (.A(_06488_),
    .B(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__buf_2 _13331_ (.A(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__a21o_1 _13332_ (.A1(_06495_),
    .A2(_06499_),
    .B1(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__mux2_1 _13333_ (.A0(_06367_),
    .A1(_06404_),
    .S(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__and4b_1 _13334_ (.A_N(_06500_),
    .B(_06495_),
    .C(_06499_),
    .D(_06365_),
    .X(_06505_));
 sky130_fd_sc_hd__nand2_2 _13335_ (.A(_06488_),
    .B(_06500_),
    .Y(_06506_));
 sky130_fd_sc_hd__or4_1 _13336_ (.A(_06408_),
    .B(_06424_),
    .C(_06490_),
    .D(_06494_),
    .X(_06507_));
 sky130_fd_sc_hd__and3_1 _13337_ (.A(_06506_),
    .B(_06507_),
    .C(_06498_),
    .X(_06508_));
 sky130_fd_sc_hd__a21oi_1 _13338_ (.A1(_06506_),
    .A2(_06507_),
    .B1(_06498_),
    .Y(_06509_));
 sky130_fd_sc_hd__a2111oi_1 _13339_ (.A1(_06495_),
    .A2(_06498_),
    .B1(_06496_),
    .C1(_06407_),
    .D1(_06502_),
    .Y(_06510_));
 sky130_fd_sc_hd__or2_1 _13340_ (.A(_06501_),
    .B(_06498_),
    .X(_06511_));
 sky130_fd_sc_hd__o221a_1 _13341_ (.A1(_06501_),
    .A2(_06495_),
    .B1(_06496_),
    .B2(_06407_),
    .C1(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__or4_1 _13342_ (.A(_06508_),
    .B(_06509_),
    .C(_06510_),
    .D(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__a21oi_2 _13343_ (.A1(_06405_),
    .A2(_06491_),
    .B1(_06407_),
    .Y(_06514_));
 sky130_fd_sc_hd__a21oi_2 _13344_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06407_),
    .Y(_06515_));
 sky130_fd_sc_hd__a21boi_1 _13345_ (.A1(_06412_),
    .A2(_06415_),
    .B1_N(_06423_),
    .Y(_06516_));
 sky130_fd_sc_hd__and3_1 _13346_ (.A(_06474_),
    .B(_06486_),
    .C(_06489_),
    .X(_06517_));
 sky130_fd_sc_hd__a31o_1 _13347_ (.A1(_06515_),
    .A2(_06516_),
    .A3(_06517_),
    .B1(_06501_),
    .X(_06518_));
 sky130_fd_sc_hd__a21oi_1 _13348_ (.A1(_06514_),
    .A2(_06518_),
    .B1(_06502_),
    .Y(_06519_));
 sky130_fd_sc_hd__xnor2_1 _13349_ (.A(_06493_),
    .B(_06519_),
    .Y(_06520_));
 sky130_fd_sc_hd__or4_4 _13350_ (.A(_06504_),
    .B(_06505_),
    .C(_06513_),
    .D(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__a21oi_1 _13351_ (.A1(_06516_),
    .A2(_06517_),
    .B1(_06502_),
    .Y(_06522_));
 sky130_fd_sc_hd__xnor2_2 _13352_ (.A(_06515_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__xor2_2 _13353_ (.A(_06514_),
    .B(_06518_),
    .X(_06524_));
 sky130_fd_sc_hd__or2_1 _13354_ (.A(_06523_),
    .B(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__or2_1 _13355_ (.A(_06521_),
    .B(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__or2_2 _13356_ (.A(_06501_),
    .B(_06474_),
    .X(_06527_));
 sky130_fd_sc_hd__xnor2_2 _13357_ (.A(_06485_),
    .B(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__and2_1 _13358_ (.A(_06474_),
    .B(_06486_),
    .X(_06529_));
 sky130_fd_sc_hd__or2_1 _13359_ (.A(_06502_),
    .B(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__xnor2_2 _13360_ (.A(_06423_),
    .B(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_1 _13361_ (.A(_06478_),
    .B(_06480_),
    .Y(_06532_));
 sky130_fd_sc_hd__a21o_1 _13362_ (.A1(_06485_),
    .A2(_06474_),
    .B1(_06502_),
    .X(_06533_));
 sky130_fd_sc_hd__xnor2_2 _13363_ (.A(_06532_),
    .B(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__nand2_1 _13364_ (.A(_06531_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__a21o_2 _13365_ (.A1(_06529_),
    .A2(_06516_),
    .B1(_06502_),
    .X(_06536_));
 sky130_fd_sc_hd__xnor2_1 _13366_ (.A(_06489_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__nand2_1 _13367_ (.A(_06412_),
    .B(_06415_),
    .Y(_06538_));
 sky130_fd_sc_hd__a21o_1 _13368_ (.A1(_06423_),
    .A2(_06529_),
    .B1(_06502_),
    .X(_06539_));
 sky130_fd_sc_hd__xnor2_2 _13369_ (.A(_06538_),
    .B(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand2_1 _13370_ (.A(_06537_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__nor2_1 _13371_ (.A(_06535_),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__nand2_1 _13372_ (.A(_06528_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__or2_2 _13373_ (.A(_06526_),
    .B(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__buf_4 _13374_ (.A(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__or2_1 _13375_ (.A(_06525_),
    .B(_06541_),
    .X(_06546_));
 sky130_fd_sc_hd__or3_4 _13376_ (.A(_06535_),
    .B(_06521_),
    .C(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__and2_2 _13377_ (.A(_06450_),
    .B(_06452_),
    .X(_06548_));
 sky130_fd_sc_hd__and2_2 _13378_ (.A(_06466_),
    .B(_06506_),
    .X(_06549_));
 sky130_fd_sc_hd__xor2_4 _13379_ (.A(_06548_),
    .B(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__or2_2 _13380_ (.A(_06501_),
    .B(_06472_),
    .X(_06551_));
 sky130_fd_sc_hd__xnor2_4 _13381_ (.A(_06443_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__nor2_2 _13382_ (.A(_06502_),
    .B(_06473_),
    .Y(_06553_));
 sky130_fd_sc_hd__xnor2_4 _13383_ (.A(_06439_),
    .B(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__o21ai_1 _13384_ (.A1(_06444_),
    .A2(_06446_),
    .B1(_06471_),
    .Y(_06555_));
 sky130_fd_sc_hd__or2_1 _13385_ (.A(_06501_),
    .B(_06467_),
    .X(_06556_));
 sky130_fd_sc_hd__xnor2_2 _13386_ (.A(_06555_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__or3_1 _13387_ (.A(_06552_),
    .B(_06554_),
    .C(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__a21o_1 _13388_ (.A1(_06439_),
    .A2(_06473_),
    .B1(_06502_),
    .X(_06559_));
 sky130_fd_sc_hd__xor2_1 _13389_ (.A(_06434_),
    .B(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__xor2_2 _13390_ (.A(_06485_),
    .B(_06527_),
    .X(_06561_));
 sky130_fd_sc_hd__nor2_1 _13391_ (.A(_06428_),
    .B(_06430_),
    .Y(_06562_));
 sky130_fd_sc_hd__a31o_1 _13392_ (.A1(_06434_),
    .A2(_06439_),
    .A3(_06473_),
    .B1(_06501_),
    .X(_06563_));
 sky130_fd_sc_hd__xnor2_2 _13393_ (.A(_06562_),
    .B(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__or3_1 _13394_ (.A(_06560_),
    .B(_06561_),
    .C(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__or3_4 _13395_ (.A(_06550_),
    .B(_06558_),
    .C(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__nor3_4 _13396_ (.A(_06466_),
    .B(_06547_),
    .C(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__a21o_2 _13397_ (.A1(_04504_),
    .A2(_06454_),
    .B1(_06456_),
    .X(_06568_));
 sky130_fd_sc_hd__o21a_2 _13398_ (.A1(_06461_),
    .A2(_06465_),
    .B1(_06506_),
    .X(_06569_));
 sky130_fd_sc_hd__xor2_2 _13399_ (.A(_06568_),
    .B(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__and2_1 _13400_ (.A(_06461_),
    .B(_06506_),
    .X(_06571_));
 sky130_fd_sc_hd__xor2_4 _13401_ (.A(_06465_),
    .B(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__nor2_1 _13402_ (.A(_06570_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__inv_2 _13403_ (.A(_06458_),
    .Y(_06574_));
 sky130_fd_sc_hd__nand2_2 _13404_ (.A(_06458_),
    .B(_06506_),
    .Y(_06575_));
 sky130_fd_sc_hd__xnor2_2 _13405_ (.A(_06460_),
    .B(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__nor2_1 _13406_ (.A(_06574_),
    .B(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__and4bb_1 _13407_ (.A_N(_06547_),
    .B_N(_06566_),
    .C(_06573_),
    .D(_06577_),
    .X(_06578_));
 sky130_fd_sc_hd__or3_1 _13408_ (.A(_06523_),
    .B(_06524_),
    .C(_06520_),
    .X(_06579_));
 sky130_fd_sc_hd__xor2_4 _13409_ (.A(_06489_),
    .B(_06536_),
    .X(_06580_));
 sky130_fd_sc_hd__and3b_1 _13410_ (.A_N(_06565_),
    .B(_06542_),
    .C(_06554_),
    .X(_06581_));
 sky130_fd_sc_hd__and4b_1 _13411_ (.A_N(_06566_),
    .B(_06542_),
    .C(_06573_),
    .D(_06576_),
    .X(_06582_));
 sky130_fd_sc_hd__nor3_1 _13412_ (.A(_06504_),
    .B(_06505_),
    .C(_06513_),
    .Y(_06583_));
 sky130_fd_sc_hd__o41a_1 _13413_ (.A1(_06579_),
    .A2(_06580_),
    .A3(_06581_),
    .A4(_06582_),
    .B1(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__or3_2 _13414_ (.A(_06567_),
    .B(_06578_),
    .C(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__or2b_1 _13415_ (.A(_06534_),
    .B_N(_06531_),
    .X(_06586_));
 sky130_fd_sc_hd__a21o_1 _13416_ (.A1(_06540_),
    .A2(_06586_),
    .B1(_06580_),
    .X(_06587_));
 sky130_fd_sc_hd__or4_4 _13417_ (.A(_06535_),
    .B(_06521_),
    .C(_06546_),
    .D(_06528_),
    .X(_06588_));
 sky130_fd_sc_hd__or3_1 _13418_ (.A(_06531_),
    .B(_06521_),
    .C(_06546_),
    .X(_06589_));
 sky130_fd_sc_hd__o211ai_4 _13419_ (.A1(_06526_),
    .A2(_06587_),
    .B1(_06588_),
    .C1(_06589_),
    .Y(_06590_));
 sky130_fd_sc_hd__or4_2 _13420_ (.A(_06535_),
    .B(_06521_),
    .C(_06546_),
    .D(_06565_),
    .X(_06591_));
 sky130_fd_sc_hd__inv_2 _13421_ (.A(_06554_),
    .Y(_06592_));
 sky130_fd_sc_hd__nand2_1 _13422_ (.A(_06552_),
    .B(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__nor2_2 _13423_ (.A(_06591_),
    .B(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__nand2_1 _13424_ (.A(_06528_),
    .B(_06564_),
    .Y(_06595_));
 sky130_fd_sc_hd__or3b_1 _13425_ (.A(_06561_),
    .B(_06564_),
    .C_N(_06560_),
    .X(_06596_));
 sky130_fd_sc_hd__or4_1 _13426_ (.A(_06535_),
    .B(_06521_),
    .C(_06546_),
    .D(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__o21ai_1 _13427_ (.A1(_06547_),
    .A2(_06595_),
    .B1(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__nor2_1 _13428_ (.A(_06592_),
    .B(_06591_),
    .Y(_06599_));
 sky130_fd_sc_hd__nor4_2 _13429_ (.A(_06590_),
    .B(_06594_),
    .C(_06598_),
    .D(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__a21oi_1 _13430_ (.A1(_06585_),
    .A2(_06600_),
    .B1(_06590_),
    .Y(_06601_));
 sky130_fd_sc_hd__clkbuf_4 _13431_ (.A(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__or2_1 _13432_ (.A(_06594_),
    .B(_06598_),
    .X(_06603_));
 sky130_fd_sc_hd__nor2_4 _13433_ (.A(_06585_),
    .B(_06603_),
    .Y(_06604_));
 sky130_fd_sc_hd__buf_2 _13434_ (.A(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__buf_2 _13435_ (.A(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__nor2_2 _13436_ (.A(_06547_),
    .B(_06566_),
    .Y(_06607_));
 sky130_fd_sc_hd__xnor2_4 _13437_ (.A(_06568_),
    .B(_06569_),
    .Y(_06608_));
 sky130_fd_sc_hd__a31oi_4 _13438_ (.A1(_06607_),
    .A2(_06608_),
    .A3(_06572_),
    .B1(_06594_),
    .Y(_06609_));
 sky130_fd_sc_hd__xor2_2 _13439_ (.A(_06460_),
    .B(_06575_),
    .X(_06610_));
 sky130_fd_sc_hd__nand2_1 _13440_ (.A(_06573_),
    .B(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__or4_1 _13441_ (.A(_06574_),
    .B(_06547_),
    .C(_06566_),
    .D(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__and2_1 _13442_ (.A(_06588_),
    .B(_06589_),
    .X(_06613_));
 sky130_fd_sc_hd__xnor2_1 _13443_ (.A(_06548_),
    .B(_06549_),
    .Y(_06614_));
 sky130_fd_sc_hd__or3_1 _13444_ (.A(_06614_),
    .B(_06558_),
    .C(_06591_),
    .X(_06615_));
 sky130_fd_sc_hd__inv_2 _13445_ (.A(_06524_),
    .Y(_06616_));
 sky130_fd_sc_hd__or3_1 _13446_ (.A(_06521_),
    .B(_06525_),
    .C(_06537_),
    .X(_06617_));
 sky130_fd_sc_hd__or2_1 _13447_ (.A(_06508_),
    .B(_06509_),
    .X(_06618_));
 sky130_fd_sc_hd__nor2_1 _13448_ (.A(_06510_),
    .B(_06512_),
    .Y(_06619_));
 sky130_fd_sc_hd__a21oi_1 _13449_ (.A1(_06618_),
    .A2(_06619_),
    .B1(_06504_),
    .Y(_06620_));
 sky130_fd_sc_hd__o2111a_1 _13450_ (.A1(_06616_),
    .A2(_06521_),
    .B1(_06617_),
    .C1(_06597_),
    .D1(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__and4_1 _13451_ (.A(_06612_),
    .B(_06613_),
    .C(_06615_),
    .D(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__nand2_4 _13452_ (.A(_06609_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__clkbuf_4 _13453_ (.A(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__buf_2 _13454_ (.A(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__buf_2 _13455_ (.A(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__or2_1 _13456_ (.A(_06585_),
    .B(_06603_),
    .X(_06627_));
 sky130_fd_sc_hd__buf_2 _13457_ (.A(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__buf_2 _13458_ (.A(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__a31o_2 _13459_ (.A1(_06607_),
    .A2(_06608_),
    .A3(_06572_),
    .B1(_06594_),
    .X(_06630_));
 sky130_fd_sc_hd__or3_1 _13460_ (.A(_06466_),
    .B(_06547_),
    .C(_06566_),
    .X(_06631_));
 sky130_fd_sc_hd__buf_4 _13461_ (.A(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__nor2_1 _13462_ (.A(_06541_),
    .B(_06586_),
    .Y(_06633_));
 sky130_fd_sc_hd__and3b_1 _13463_ (.A_N(_06566_),
    .B(_06542_),
    .C(_06570_),
    .X(_06634_));
 sky130_fd_sc_hd__nor2_1 _13464_ (.A(_06524_),
    .B(_06521_),
    .Y(_06635_));
 sky130_fd_sc_hd__o31ai_1 _13465_ (.A1(_06523_),
    .A2(_06633_),
    .A3(_06634_),
    .B1(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__or3b_1 _13466_ (.A(_06504_),
    .B(_06505_),
    .C_N(_06513_),
    .X(_06637_));
 sky130_fd_sc_hd__o211a_1 _13467_ (.A1(_06592_),
    .A2(_06591_),
    .B1(_06588_),
    .C1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__nand4_2 _13468_ (.A(_06632_),
    .B(_06617_),
    .C(_06636_),
    .D(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__nor2_2 _13469_ (.A(_06630_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__clkbuf_4 _13470_ (.A(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__clkbuf_4 _13471_ (.A(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__buf_2 _13472_ (.A(_06609_),
    .X(_06643_));
 sky130_fd_sc_hd__buf_2 _13473_ (.A(_06622_),
    .X(_06644_));
 sky130_fd_sc_hd__and3_1 _13474_ (.A(_06531_),
    .B(_06643_),
    .C(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__a21oi_1 _13475_ (.A1(_06534_),
    .A2(_06624_),
    .B1(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__a21o_1 _13476_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06564_),
    .X(_06647_));
 sky130_fd_sc_hd__and4_2 _13477_ (.A(_06632_),
    .B(_06617_),
    .C(_06636_),
    .D(_06638_),
    .X(_06648_));
 sky130_fd_sc_hd__nand2_2 _13478_ (.A(_06609_),
    .B(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__buf_2 _13479_ (.A(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__o211a_1 _13480_ (.A1(_06561_),
    .A2(_06623_),
    .B1(_06647_),
    .C1(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__a21o_1 _13481_ (.A1(_06642_),
    .A2(_06646_),
    .B1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__nand4_4 _13482_ (.A(_06612_),
    .B(_06613_),
    .C(_06615_),
    .D(_06621_),
    .Y(_06653_));
 sky130_fd_sc_hd__or3_1 _13483_ (.A(_06552_),
    .B(_06630_),
    .C(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__a21o_1 _13484_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06557_),
    .X(_06655_));
 sky130_fd_sc_hd__a21oi_1 _13485_ (.A1(_06654_),
    .A2(_06655_),
    .B1(_06640_),
    .Y(_06656_));
 sky130_fd_sc_hd__a21o_1 _13486_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06554_),
    .X(_06657_));
 sky130_fd_sc_hd__or3_1 _13487_ (.A(_06560_),
    .B(_06630_),
    .C(_06653_),
    .X(_06658_));
 sky130_fd_sc_hd__a21oi_1 _13488_ (.A1(_06657_),
    .A2(_06658_),
    .B1(_06649_),
    .Y(_06659_));
 sky130_fd_sc_hd__a21o_1 _13489_ (.A1(_06585_),
    .A2(_06600_),
    .B1(_06590_),
    .X(_06660_));
 sky130_fd_sc_hd__buf_4 _13490_ (.A(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__o31a_1 _13491_ (.A1(_06629_),
    .A2(_06656_),
    .A3(_06659_),
    .B1(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__a21bo_1 _13492_ (.A1(_06629_),
    .A2(_06652_),
    .B1_N(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__nand2_1 _13493_ (.A(_06600_),
    .B(_06605_),
    .Y(_06664_));
 sky130_fd_sc_hd__inv_2 _13494_ (.A(_06540_),
    .Y(_06665_));
 sky130_fd_sc_hd__mux2_1 _13495_ (.A0(_06580_),
    .A1(_06665_),
    .S(_06623_),
    .X(_06666_));
 sky130_fd_sc_hd__nor2_1 _13496_ (.A(_06630_),
    .B(_06653_),
    .Y(_06667_));
 sky130_fd_sc_hd__clkbuf_4 _13497_ (.A(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__mux2_1 _13498_ (.A0(_06523_),
    .A1(_06524_),
    .S(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__mux2_1 _13499_ (.A0(_06666_),
    .A1(_06669_),
    .S(_06641_),
    .X(_06670_));
 sky130_fd_sc_hd__o21a_1 _13500_ (.A1(_06664_),
    .A2(_06670_),
    .B1(_06545_),
    .X(_06671_));
 sky130_fd_sc_hd__a21o_4 _13501_ (.A1(_06639_),
    .A2(_06653_),
    .B1(_06630_),
    .X(_06672_));
 sky130_fd_sc_hd__xnor2_4 _13502_ (.A(_06604_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nor2_1 _13503_ (.A(_06526_),
    .B(_06543_),
    .Y(_06674_));
 sky130_fd_sc_hd__o311a_4 _13504_ (.A1(_06629_),
    .A2(_06641_),
    .A3(_06668_),
    .B1(_06602_),
    .C1(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__nand2_1 _13505_ (.A(_06673_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__inv_2 _13506_ (.A(_06572_),
    .Y(_06677_));
 sky130_fd_sc_hd__mux2_1 _13507_ (.A0(_06608_),
    .A1(_06677_),
    .S(_06668_),
    .X(_06678_));
 sky130_fd_sc_hd__o21ai_1 _13508_ (.A1(_06550_),
    .A2(_06624_),
    .B1(_06655_),
    .Y(_06679_));
 sky130_fd_sc_hd__a21o_1 _13509_ (.A1(_06648_),
    .A2(_06668_),
    .B1(_06672_),
    .X(_06680_));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(_06678_),
    .A1(_06679_),
    .S(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__a21oi_4 _13511_ (.A1(_06648_),
    .A2(_06667_),
    .B1(_06672_),
    .Y(_06682_));
 sky130_fd_sc_hd__a21o_1 _13512_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06576_),
    .X(_06683_));
 sky130_fd_sc_hd__o21ai_1 _13513_ (.A1(_06458_),
    .A2(_06624_),
    .B1(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__or4_1 _13514_ (.A(_06544_),
    .B(_06673_),
    .C(_06682_),
    .D(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__o21ai_2 _13515_ (.A1(_06676_),
    .A2(_06681_),
    .B1(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__a21oi_4 _13516_ (.A1(_06663_),
    .A2(_06671_),
    .B1(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__clkbuf_4 _13517_ (.A(_06687_),
    .X(_06688_));
 sky130_fd_sc_hd__or3_1 _13518_ (.A(_06605_),
    .B(_06656_),
    .C(_06659_),
    .X(_06689_));
 sky130_fd_sc_hd__o211ai_1 _13519_ (.A1(_06572_),
    .A2(_06623_),
    .B1(_06683_),
    .C1(_06650_),
    .Y(_06690_));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(_06614_),
    .A1(_06608_),
    .S(_06623_),
    .X(_06691_));
 sky130_fd_sc_hd__nand2_2 _13521_ (.A(_06604_),
    .B(_06640_),
    .Y(_06692_));
 sky130_fd_sc_hd__o221a_1 _13522_ (.A1(_06629_),
    .A2(_06690_),
    .B1(_06691_),
    .B2(_06692_),
    .C1(_06660_),
    .X(_06693_));
 sky130_fd_sc_hd__a211oi_1 _13523_ (.A1(_06641_),
    .A2(_06646_),
    .B1(_06651_),
    .C1(_06664_),
    .Y(_06694_));
 sky130_fd_sc_hd__buf_4 _13524_ (.A(_06674_),
    .X(_06695_));
 sky130_fd_sc_hd__a211o_4 _13525_ (.A1(_06689_),
    .A2(_06693_),
    .B1(_06694_),
    .C1(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__a211o_4 _13526_ (.A1(_06604_),
    .A2(_06672_),
    .B1(_06660_),
    .C1(_06544_),
    .X(_06697_));
 sky130_fd_sc_hd__xnor2_4 _13527_ (.A(_06628_),
    .B(_06672_),
    .Y(_06698_));
 sky130_fd_sc_hd__or3_1 _13528_ (.A(_06698_),
    .B(_06682_),
    .C(_06684_),
    .X(_06699_));
 sky130_fd_sc_hd__or2_4 _13529_ (.A(_06697_),
    .B(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__or3_1 _13530_ (.A(_06554_),
    .B(_06630_),
    .C(_06653_),
    .X(_06701_));
 sky130_fd_sc_hd__a21o_1 _13531_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06552_),
    .X(_06702_));
 sky130_fd_sc_hd__a21o_1 _13532_ (.A1(_06701_),
    .A2(_06702_),
    .B1(_06649_),
    .X(_06703_));
 sky130_fd_sc_hd__and3_1 _13533_ (.A(_06557_),
    .B(_06609_),
    .C(_06622_),
    .X(_06704_));
 sky130_fd_sc_hd__a211o_1 _13534_ (.A1(_06550_),
    .A2(_06623_),
    .B1(_06704_),
    .C1(_06640_),
    .X(_06705_));
 sky130_fd_sc_hd__a21oi_1 _13535_ (.A1(_06703_),
    .A2(_06705_),
    .B1(_06605_),
    .Y(_06706_));
 sky130_fd_sc_hd__nand2_1 _13536_ (.A(_06458_),
    .B(_06624_),
    .Y(_06707_));
 sky130_fd_sc_hd__nor2_2 _13537_ (.A(_06628_),
    .B(_06640_),
    .Y(_06708_));
 sky130_fd_sc_hd__o211a_1 _13538_ (.A1(_06610_),
    .A2(_06624_),
    .B1(_06707_),
    .C1(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__mux2_1 _13539_ (.A0(_06570_),
    .A1(_06572_),
    .S(_06623_),
    .X(_06710_));
 sky130_fd_sc_hd__nor2_1 _13540_ (.A(_06692_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__o31a_4 _13541_ (.A1(_06706_),
    .A2(_06709_),
    .A3(_06711_),
    .B1(_06661_),
    .X(_06712_));
 sky130_fd_sc_hd__and3_1 _13542_ (.A(_06665_),
    .B(_06643_),
    .C(_06644_),
    .X(_06713_));
 sky130_fd_sc_hd__a21oi_1 _13543_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06531_),
    .Y(_06714_));
 sky130_fd_sc_hd__or3_1 _13544_ (.A(_06640_),
    .B(_06713_),
    .C(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__and3_1 _13545_ (.A(_06523_),
    .B(_06643_),
    .C(_06644_),
    .X(_06716_));
 sky130_fd_sc_hd__a211o_1 _13546_ (.A1(_06580_),
    .A2(_06623_),
    .B1(_06716_),
    .C1(_06649_),
    .X(_06717_));
 sky130_fd_sc_hd__and3_1 _13547_ (.A(_06629_),
    .B(_06715_),
    .C(_06717_),
    .X(_06718_));
 sky130_fd_sc_hd__a21o_1 _13548_ (.A1(_06643_),
    .A2(_06644_),
    .B1(_06560_),
    .X(_06719_));
 sky130_fd_sc_hd__or3_1 _13549_ (.A(_06564_),
    .B(_06630_),
    .C(_06653_),
    .X(_06720_));
 sky130_fd_sc_hd__a21oi_1 _13550_ (.A1(_06719_),
    .A2(_06720_),
    .B1(_06641_),
    .Y(_06721_));
 sky130_fd_sc_hd__or3_1 _13551_ (.A(_06534_),
    .B(_06630_),
    .C(_06653_),
    .X(_06722_));
 sky130_fd_sc_hd__o211a_1 _13552_ (.A1(_06528_),
    .A2(_06668_),
    .B1(_06722_),
    .C1(_06641_),
    .X(_06723_));
 sky130_fd_sc_hd__nor3_1 _13553_ (.A(_06629_),
    .B(_06721_),
    .C(_06723_),
    .Y(_06724_));
 sky130_fd_sc_hd__nor3_4 _13554_ (.A(_06661_),
    .B(_06718_),
    .C(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__a211o_4 _13555_ (.A1(_06696_),
    .A2(_06700_),
    .B1(_06712_),
    .C1(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__and3_1 _13556_ (.A(_06640_),
    .B(_06719_),
    .C(_06720_),
    .X(_06727_));
 sky130_fd_sc_hd__a31o_1 _13557_ (.A1(_06650_),
    .A2(_06701_),
    .A3(_06702_),
    .B1(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__nor2_1 _13558_ (.A(_06628_),
    .B(_06649_),
    .Y(_06729_));
 sky130_fd_sc_hd__a21o_1 _13559_ (.A1(_06550_),
    .A2(_06623_),
    .B1(_06704_),
    .X(_06730_));
 sky130_fd_sc_hd__a221o_1 _13560_ (.A1(_06729_),
    .A2(_06730_),
    .B1(_06710_),
    .B2(_06708_),
    .C1(_06601_),
    .X(_06731_));
 sky130_fd_sc_hd__a21o_1 _13561_ (.A1(_06629_),
    .A2(_06728_),
    .B1(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__o21a_1 _13562_ (.A1(_06528_),
    .A2(_06668_),
    .B1(_06722_),
    .X(_06733_));
 sky130_fd_sc_hd__or3_1 _13563_ (.A(_06649_),
    .B(_06713_),
    .C(_06714_),
    .X(_06734_));
 sky130_fd_sc_hd__a21bo_1 _13564_ (.A1(_06650_),
    .A2(_06733_),
    .B1_N(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__nand2_1 _13565_ (.A(_06605_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__nor2_1 _13566_ (.A(_06698_),
    .B(_06697_),
    .Y(_06737_));
 sky130_fd_sc_hd__mux2_1 _13567_ (.A0(_06572_),
    .A1(_06576_),
    .S(_06668_),
    .X(_06738_));
 sky130_fd_sc_hd__clkbuf_4 _13568_ (.A(_06680_),
    .X(_06739_));
 sky130_fd_sc_hd__a2bb2o_1 _13569_ (.A1_N(_06650_),
    .A2_N(_06707_),
    .B1(_06738_),
    .B2(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__a32oi_4 _13570_ (.A1(_06545_),
    .A2(_06732_),
    .A3(_06736_),
    .B1(_06737_),
    .B2(_06740_),
    .Y(_06741_));
 sky130_fd_sc_hd__nor2_1 _13571_ (.A(_06721_),
    .B(_06723_),
    .Y(_06742_));
 sky130_fd_sc_hd__a31o_1 _13572_ (.A1(_06605_),
    .A2(_06703_),
    .A3(_06705_),
    .B1(_06602_),
    .X(_06743_));
 sky130_fd_sc_hd__a21o_1 _13573_ (.A1(_06629_),
    .A2(_06742_),
    .B1(_06743_),
    .X(_06744_));
 sky130_fd_sc_hd__a21o_1 _13574_ (.A1(_06715_),
    .A2(_06717_),
    .B1(_06664_),
    .X(_06745_));
 sky130_fd_sc_hd__mux2_1 _13575_ (.A0(_06550_),
    .A1(_06570_),
    .S(_06668_),
    .X(_06746_));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(_06746_),
    .A1(_06738_),
    .S(_06682_),
    .X(_06747_));
 sky130_fd_sc_hd__or4_1 _13577_ (.A(_06605_),
    .B(_06641_),
    .C(_06697_),
    .D(_06707_),
    .X(_06748_));
 sky130_fd_sc_hd__a21bo_1 _13578_ (.A1(_06737_),
    .A2(_06747_),
    .B1_N(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__a31oi_4 _13579_ (.A1(_06545_),
    .A2(_06744_),
    .A3(_06745_),
    .B1(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__buf_2 _13580_ (.A(_06629_),
    .X(_06751_));
 sky130_fd_sc_hd__o211a_1 _13581_ (.A1(_06561_),
    .A2(_06624_),
    .B1(_06647_),
    .C1(_06641_),
    .X(_06752_));
 sky130_fd_sc_hd__a31o_1 _13582_ (.A1(_06650_),
    .A2(_06657_),
    .A3(_06658_),
    .B1(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__nand2_1 _13583_ (.A(_06605_),
    .B(_06650_),
    .Y(_06754_));
 sky130_fd_sc_hd__nand2_1 _13584_ (.A(_06654_),
    .B(_06655_),
    .Y(_06755_));
 sky130_fd_sc_hd__o221a_1 _13585_ (.A1(_06754_),
    .A2(_06691_),
    .B1(_06692_),
    .B2(_06755_),
    .C1(_06660_),
    .X(_06756_));
 sky130_fd_sc_hd__a21boi_1 _13586_ (.A1(_06751_),
    .A2(_06753_),
    .B1_N(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__mux2_1 _13587_ (.A0(_06666_),
    .A1(_06646_),
    .S(_06650_),
    .X(_06758_));
 sky130_fd_sc_hd__nor2_1 _13588_ (.A(_06664_),
    .B(_06758_),
    .Y(_06759_));
 sky130_fd_sc_hd__mux4_2 _13589_ (.A0(_06574_),
    .A1(_06608_),
    .A2(_06677_),
    .A3(_06610_),
    .S0(_06624_),
    .S1(_06641_),
    .X(_06760_));
 sky130_fd_sc_hd__o32a_4 _13590_ (.A1(_06695_),
    .A2(_06757_),
    .A3(_06759_),
    .B1(_06676_),
    .B2(_06760_),
    .X(_06761_));
 sky130_fd_sc_hd__a2111o_4 _13591_ (.A1(_06726_),
    .A2(_06741_),
    .B1(_06750_),
    .C1(_06761_),
    .D1(_06687_),
    .X(_06762_));
 sky130_fd_sc_hd__nor2_1 _13592_ (.A(_06629_),
    .B(_06728_),
    .Y(_06763_));
 sky130_fd_sc_hd__a211o_1 _13593_ (.A1(_06751_),
    .A2(_06735_),
    .B1(_06763_),
    .C1(_06602_),
    .X(_06764_));
 sky130_fd_sc_hd__a21oi_1 _13594_ (.A1(_06552_),
    .A2(_06624_),
    .B1(_06704_),
    .Y(_06765_));
 sky130_fd_sc_hd__nor2_1 _13595_ (.A(_06682_),
    .B(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__a211o_1 _13596_ (.A1(_06682_),
    .A2(_06746_),
    .B1(_06766_),
    .C1(_06698_),
    .X(_06767_));
 sky130_fd_sc_hd__o211ai_1 _13597_ (.A1(_06673_),
    .A2(_06740_),
    .B1(_06767_),
    .C1(_06675_),
    .Y(_06768_));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(_06524_),
    .A1(_06520_),
    .S(_06668_),
    .X(_06769_));
 sky130_fd_sc_hd__a21oi_1 _13599_ (.A1(_06580_),
    .A2(_06625_),
    .B1(_06716_),
    .Y(_06770_));
 sky130_fd_sc_hd__o2bb2a_1 _13600_ (.A1_N(_06769_),
    .A2_N(_06729_),
    .B1(_06754_),
    .B2(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__and3_1 _13601_ (.A(_06764_),
    .B(_06768_),
    .C(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__clkbuf_4 _13602_ (.A(_06772_),
    .X(_06773_));
 sky130_fd_sc_hd__mux2_1 _13603_ (.A0(_06758_),
    .A1(_06753_),
    .S(_06605_),
    .X(_06774_));
 sky130_fd_sc_hd__and3b_1 _13604_ (.A_N(_06760_),
    .B(_06698_),
    .C(_06695_),
    .X(_06775_));
 sky130_fd_sc_hd__mux2_1 _13605_ (.A0(_06618_),
    .A1(_06520_),
    .S(_06624_),
    .X(_06776_));
 sky130_fd_sc_hd__mux2_1 _13606_ (.A0(_06669_),
    .A1(_06776_),
    .S(_06642_),
    .X(_06777_));
 sky130_fd_sc_hd__mux4_1 _13607_ (.A0(_06550_),
    .A1(_06552_),
    .A2(_06554_),
    .A3(_06557_),
    .S0(_06641_),
    .S1(_06625_),
    .X(_06778_));
 sky130_fd_sc_hd__and3_1 _13608_ (.A(_06673_),
    .B(_06675_),
    .C(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__or3_2 _13609_ (.A(_06775_),
    .B(_06777_),
    .C(_06779_),
    .X(_06780_));
 sky130_fd_sc_hd__a21oi_4 _13610_ (.A1(_06661_),
    .A2(_06774_),
    .B1(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__a21o_1 _13611_ (.A1(_06762_),
    .A2(_06773_),
    .B1(_06781_),
    .X(_06782_));
 sky130_fd_sc_hd__buf_6 _13612_ (.A(_06782_),
    .X(_06783_));
 sky130_fd_sc_hd__nand3_4 _13613_ (.A(_06781_),
    .B(_06762_),
    .C(_06773_),
    .Y(_06784_));
 sky130_fd_sc_hd__and2_1 _13614_ (.A(_06783_),
    .B(_06784_),
    .X(_06785_));
 sky130_fd_sc_hd__or2_1 _13615_ (.A(_06688_),
    .B(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__xnor2_4 _13616_ (.A(_06762_),
    .B(_06773_),
    .Y(_06787_));
 sky130_fd_sc_hd__or2_1 _13617_ (.A(_06750_),
    .B(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__buf_2 _13618_ (.A(_06761_),
    .X(_06789_));
 sky130_fd_sc_hd__or2_1 _13619_ (.A(_06718_),
    .B(_06724_),
    .X(_06790_));
 sky130_fd_sc_hd__and2_1 _13620_ (.A(_06618_),
    .B(_06625_),
    .X(_06791_));
 sky130_fd_sc_hd__buf_2 _13621_ (.A(_06650_),
    .X(_06792_));
 sky130_fd_sc_hd__mux2_1 _13622_ (.A0(_06791_),
    .A1(_06769_),
    .S(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__a211o_1 _13623_ (.A1(_06661_),
    .A2(_06790_),
    .B1(_06793_),
    .C1(_06695_),
    .X(_06794_));
 sky130_fd_sc_hd__nand2_4 _13624_ (.A(_06607_),
    .B(_06608_),
    .Y(_06795_));
 sky130_fd_sc_hd__a31o_1 _13625_ (.A1(_06458_),
    .A2(_06605_),
    .A3(_06672_),
    .B1(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__nand2_1 _13626_ (.A(_06719_),
    .B(_06701_),
    .Y(_06797_));
 sky130_fd_sc_hd__mux2_1 _13627_ (.A0(_06797_),
    .A1(_06765_),
    .S(_06682_),
    .X(_06798_));
 sky130_fd_sc_hd__nor2_1 _13628_ (.A(_06698_),
    .B(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__a211o_1 _13629_ (.A1(_06698_),
    .A2(_06747_),
    .B1(_06799_),
    .C1(_06697_),
    .X(_06800_));
 sky130_fd_sc_hd__and3_2 _13630_ (.A(_06794_),
    .B(_06796_),
    .C(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__clkbuf_4 _13631_ (.A(_06801_),
    .X(_06802_));
 sky130_fd_sc_hd__xnor2_4 _13632_ (.A(_06802_),
    .B(_06783_),
    .Y(_06803_));
 sky130_fd_sc_hd__nor2_1 _13633_ (.A(_06688_),
    .B(_06787_),
    .Y(_06804_));
 sky130_fd_sc_hd__a21oi_1 _13634_ (.A1(_06783_),
    .A2(_06784_),
    .B1(_06750_),
    .Y(_06805_));
 sky130_fd_sc_hd__xnor2_1 _13635_ (.A(_06804_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__or3_1 _13636_ (.A(_06789_),
    .B(_06803_),
    .C(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__o21ai_1 _13637_ (.A1(_06786_),
    .A2(_06788_),
    .B1(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__clkinv_2 _13638_ (.A(_06801_),
    .Y(_06809_));
 sky130_fd_sc_hd__a211oi_4 _13639_ (.A1(_06696_),
    .A2(_06700_),
    .B1(_06712_),
    .C1(_06725_),
    .Y(_06810_));
 sky130_fd_sc_hd__nand2_1 _13640_ (.A(_06741_),
    .B(_06761_),
    .Y(_06811_));
 sky130_fd_sc_hd__a21o_1 _13641_ (.A1(_06726_),
    .A2(_06741_),
    .B1(_06761_),
    .X(_06812_));
 sky130_fd_sc_hd__o21a_2 _13642_ (.A1(_06810_),
    .A2(_06811_),
    .B1(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__clkbuf_4 _13643_ (.A(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__nor2_1 _13644_ (.A(_06809_),
    .B(_06814_),
    .Y(_06815_));
 sky130_fd_sc_hd__clkbuf_4 _13645_ (.A(_06781_),
    .X(_06816_));
 sky130_fd_sc_hd__xor2_1 _13646_ (.A(_06750_),
    .B(_06812_),
    .X(_06817_));
 sky130_fd_sc_hd__clkbuf_4 _13647_ (.A(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__nor2_1 _13648_ (.A(_06816_),
    .B(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__clkbuf_4 _13649_ (.A(_06773_),
    .X(_06820_));
 sky130_fd_sc_hd__nand2_1 _13650_ (.A(_06726_),
    .B(_06741_),
    .Y(_06821_));
 sky130_fd_sc_hd__nor2_2 _13651_ (.A(_06750_),
    .B(_06761_),
    .Y(_06822_));
 sky130_fd_sc_hd__nand2_4 _13652_ (.A(_06821_),
    .B(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__xor2_4 _13653_ (.A(_06823_),
    .B(_06687_),
    .X(_06824_));
 sky130_fd_sc_hd__nor2_1 _13654_ (.A(_06820_),
    .B(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__o21ai_2 _13655_ (.A1(_06810_),
    .A2(_06811_),
    .B1(_06812_),
    .Y(_06826_));
 sky130_fd_sc_hd__nand2_1 _13656_ (.A(_06802_),
    .B(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__xnor2_1 _13657_ (.A(_06827_),
    .B(_06819_),
    .Y(_06828_));
 sky130_fd_sc_hd__a22o_1 _13658_ (.A1(_06815_),
    .A2(_06819_),
    .B1(_06825_),
    .B2(_06828_),
    .X(_06829_));
 sky130_fd_sc_hd__buf_2 _13659_ (.A(_06750_),
    .X(_06830_));
 sky130_fd_sc_hd__nor2_1 _13660_ (.A(_06830_),
    .B(_06803_),
    .Y(_06831_));
 sky130_fd_sc_hd__nor2_2 _13661_ (.A(_06823_),
    .B(_06687_),
    .Y(_06832_));
 sky130_fd_sc_hd__nor2_1 _13662_ (.A(_06832_),
    .B(_06820_),
    .Y(_06833_));
 sky130_fd_sc_hd__xnor2_1 _13663_ (.A(_06786_),
    .B(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__xnor2_1 _13664_ (.A(_06831_),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__xnor2_1 _13665_ (.A(_06829_),
    .B(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__and2b_1 _13666_ (.A_N(_06835_),
    .B(_06829_),
    .X(_06837_));
 sky130_fd_sc_hd__a21o_1 _13667_ (.A1(_06808_),
    .A2(_06836_),
    .B1(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__nor2_4 _13668_ (.A(_06809_),
    .B(_06783_),
    .Y(_06839_));
 sky130_fd_sc_hd__inv_2 _13669_ (.A(_06699_),
    .Y(_06840_));
 sky130_fd_sc_hd__nand2_1 _13670_ (.A(_06657_),
    .B(_06654_),
    .Y(_06841_));
 sky130_fd_sc_hd__nand2_1 _13671_ (.A(_06647_),
    .B(_06658_),
    .Y(_06842_));
 sky130_fd_sc_hd__mux4_1 _13672_ (.A0(_06678_),
    .A1(_06841_),
    .A2(_06679_),
    .A3(_06842_),
    .S0(_06673_),
    .S1(_06739_),
    .X(_06843_));
 sky130_fd_sc_hd__inv_2 _13673_ (.A(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__buf_2 _13674_ (.A(_06668_),
    .X(_06845_));
 sky130_fd_sc_hd__nor2_1 _13675_ (.A(_06619_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__a211o_1 _13676_ (.A1(_06650_),
    .A2(_06776_),
    .B1(_06846_),
    .C1(_06695_),
    .X(_06847_));
 sky130_fd_sc_hd__a221o_1 _13677_ (.A1(_06590_),
    .A2(_06652_),
    .B1(_06670_),
    .B2(_06751_),
    .C1(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__o221a_1 _13678_ (.A1(_06795_),
    .A2(_06840_),
    .B1(_06844_),
    .B2(_06697_),
    .C1(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__clkbuf_4 _13679_ (.A(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__a21o_2 _13680_ (.A1(_06839_),
    .A2(_06850_),
    .B1(_06567_),
    .X(_06851_));
 sky130_fd_sc_hd__or2_1 _13681_ (.A(_06789_),
    .B(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__clkbuf_4 _13682_ (.A(_06741_),
    .X(_06853_));
 sky130_fd_sc_hd__xor2_4 _13683_ (.A(_06839_),
    .B(_06850_),
    .X(_06854_));
 sky130_fd_sc_hd__or2_1 _13684_ (.A(_06853_),
    .B(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__or2_1 _13685_ (.A(_06852_),
    .B(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__or2_1 _13686_ (.A(_06789_),
    .B(_06854_),
    .X(_06857_));
 sky130_fd_sc_hd__or2_1 _13687_ (.A(_06830_),
    .B(_06851_),
    .X(_06858_));
 sky130_fd_sc_hd__nor2_1 _13688_ (.A(_06857_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__o21a_1 _13689_ (.A1(_06830_),
    .A2(_06854_),
    .B1(_06852_),
    .X(_06860_));
 sky130_fd_sc_hd__nor2_1 _13690_ (.A(_06859_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__xnor2_1 _13691_ (.A(_06856_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__nand2_8 _13692_ (.A(_06696_),
    .B(_06700_),
    .Y(_06863_));
 sky130_fd_sc_hd__clkinv_4 _13693_ (.A(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__or2_1 _13694_ (.A(_06864_),
    .B(_06854_),
    .X(_06865_));
 sky130_fd_sc_hd__or4b_1 _13695_ (.A(_06853_),
    .B(_06851_),
    .C(_06865_),
    .D_N(_06857_),
    .X(_06866_));
 sky130_fd_sc_hd__xnor2_1 _13696_ (.A(_06838_),
    .B(_06862_),
    .Y(_06867_));
 sky130_fd_sc_hd__nor2_1 _13697_ (.A(_06866_),
    .B(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__a21o_1 _13698_ (.A1(_06838_),
    .A2(_06862_),
    .B1(_06868_),
    .X(_06869_));
 sky130_fd_sc_hd__xnor2_4 _13699_ (.A(_06810_),
    .B(_06741_),
    .Y(_06870_));
 sky130_fd_sc_hd__nor2_8 _13700_ (.A(_06712_),
    .B(_06725_),
    .Y(_06871_));
 sky130_fd_sc_hd__xnor2_4 _13701_ (.A(_06863_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__and4_1 _13702_ (.A(_06632_),
    .B(_06850_),
    .C(_06870_),
    .D(_06872_),
    .X(_06873_));
 sky130_fd_sc_hd__a22o_1 _13703_ (.A1(_06850_),
    .A2(_06870_),
    .B1(_06872_),
    .B2(_06632_),
    .X(_06874_));
 sky130_fd_sc_hd__or2b_1 _13704_ (.A(_06873_),
    .B_N(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__and2_1 _13705_ (.A(_06871_),
    .B(_06849_),
    .X(_06876_));
 sky130_fd_sc_hd__xnor2_4 _13706_ (.A(_06726_),
    .B(_06741_),
    .Y(_06877_));
 sky130_fd_sc_hd__or2_1 _13707_ (.A(_06712_),
    .B(_06725_),
    .X(_06878_));
 sky130_fd_sc_hd__clkbuf_4 _13708_ (.A(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__mux2_1 _13709_ (.A0(_06879_),
    .A1(_06863_),
    .S(_06849_),
    .X(_06880_));
 sky130_fd_sc_hd__or3b_1 _13710_ (.A(_06877_),
    .B(_06880_),
    .C_N(_06801_),
    .X(_06881_));
 sky130_fd_sc_hd__a21bo_1 _13711_ (.A1(_06863_),
    .A2(_06876_),
    .B1_N(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__and2b_1 _13712_ (.A_N(_06875_),
    .B(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__xor2_1 _13713_ (.A(_06875_),
    .B(_06882_),
    .X(_06884_));
 sky130_fd_sc_hd__xnor2_1 _13714_ (.A(_06825_),
    .B(_06828_),
    .Y(_06885_));
 sky130_fd_sc_hd__nor2_1 _13715_ (.A(_06884_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__or2_1 _13716_ (.A(_06877_),
    .B(_06873_),
    .X(_06887_));
 sky130_fd_sc_hd__nor2_1 _13717_ (.A(_06816_),
    .B(_06824_),
    .Y(_06888_));
 sky130_fd_sc_hd__nand2b_2 _13718_ (.A_N(_06818_),
    .B(_06850_),
    .Y(_06889_));
 sky130_fd_sc_hd__a2bb2o_1 _13719_ (.A1_N(_06809_),
    .A2_N(_06818_),
    .B1(_06826_),
    .B2(_06850_),
    .X(_06890_));
 sky130_fd_sc_hd__o21a_1 _13720_ (.A1(_06827_),
    .A2(_06889_),
    .B1(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__xor2_1 _13721_ (.A(_06888_),
    .B(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__xnor2_1 _13722_ (.A(_06887_),
    .B(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__o21ai_2 _13723_ (.A1(_06883_),
    .A2(_06886_),
    .B1(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__or3_1 _13724_ (.A(_06893_),
    .B(_06883_),
    .C(_06886_),
    .X(_06895_));
 sky130_fd_sc_hd__and2_1 _13725_ (.A(_06894_),
    .B(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__xor2_1 _13726_ (.A(_06808_),
    .B(_06836_),
    .X(_06897_));
 sky130_fd_sc_hd__nand2_1 _13727_ (.A(_06896_),
    .B(_06897_),
    .Y(_06898_));
 sky130_fd_sc_hd__nor2_1 _13728_ (.A(_06813_),
    .B(_06889_),
    .Y(_06899_));
 sky130_fd_sc_hd__o21ai_1 _13729_ (.A1(_06567_),
    .A2(_06813_),
    .B1(_06889_),
    .Y(_06900_));
 sky130_fd_sc_hd__and2b_1 _13730_ (.A_N(_06899_),
    .B(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__nand2_1 _13731_ (.A(_06823_),
    .B(_06688_),
    .Y(_06902_));
 sky130_fd_sc_hd__nand2_2 _13732_ (.A(_06762_),
    .B(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand2_1 _13733_ (.A(_06802_),
    .B(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__xnor2_1 _13734_ (.A(_06901_),
    .B(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__a21oi_1 _13735_ (.A1(_06870_),
    .A2(_06892_),
    .B1(_06873_),
    .Y(_06906_));
 sky130_fd_sc_hd__xnor2_1 _13736_ (.A(_06905_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__or3_1 _13737_ (.A(_06832_),
    .B(_06820_),
    .C(_06786_),
    .X(_06908_));
 sky130_fd_sc_hd__a21bo_1 _13738_ (.A1(_06831_),
    .A2(_06834_),
    .B1_N(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__o2bb2a_1 _13739_ (.A1_N(_06888_),
    .A2_N(_06890_),
    .B1(_06889_),
    .B2(_06827_),
    .X(_06910_));
 sky130_fd_sc_hd__xnor2_1 _13740_ (.A(_06809_),
    .B(_06782_),
    .Y(_06911_));
 sky130_fd_sc_hd__clkbuf_4 _13741_ (.A(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__or2_1 _13742_ (.A(_06688_),
    .B(_06803_),
    .X(_06913_));
 sky130_fd_sc_hd__or2_1 _13743_ (.A(_06816_),
    .B(_06762_),
    .X(_06914_));
 sky130_fd_sc_hd__mux2_1 _13744_ (.A0(_06912_),
    .A1(_06913_),
    .S(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__xnor2_1 _13745_ (.A(_06910_),
    .B(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__xnor2_1 _13746_ (.A(_06909_),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__xnor2_1 _13747_ (.A(_06907_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__a21o_1 _13748_ (.A1(_06894_),
    .A2(_06898_),
    .B1(_06918_),
    .X(_06919_));
 sky130_fd_sc_hd__nand3_1 _13749_ (.A(_06894_),
    .B(_06898_),
    .C(_06918_),
    .Y(_06920_));
 sky130_fd_sc_hd__nand2_1 _13750_ (.A(_06919_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__and2_1 _13751_ (.A(_06866_),
    .B(_06867_),
    .X(_06922_));
 sky130_fd_sc_hd__nor2_1 _13752_ (.A(_06868_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__or2b_1 _13753_ (.A(_06921_),
    .B_N(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__or2b_1 _13754_ (.A(_06906_),
    .B_N(_06905_),
    .X(_06925_));
 sky130_fd_sc_hd__a21bo_1 _13755_ (.A1(_06907_),
    .A2(_06917_),
    .B1_N(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__nand2_1 _13756_ (.A(_06632_),
    .B(_06903_),
    .Y(_06927_));
 sky130_fd_sc_hd__or2_1 _13757_ (.A(_06889_),
    .B(_06927_),
    .X(_06928_));
 sky130_fd_sc_hd__a2bb2o_1 _13758_ (.A1_N(_06567_),
    .A2_N(_06818_),
    .B1(_06903_),
    .B2(_06850_),
    .X(_06929_));
 sky130_fd_sc_hd__and2_1 _13759_ (.A(_06928_),
    .B(_06929_),
    .X(_06930_));
 sky130_fd_sc_hd__a31o_1 _13760_ (.A1(_06802_),
    .A2(_06903_),
    .A3(_06901_),
    .B1(_06899_),
    .X(_06931_));
 sky130_fd_sc_hd__inv_2 _13761_ (.A(_06787_),
    .Y(_06932_));
 sky130_fd_sc_hd__o2bb2a_1 _13762_ (.A1_N(_06820_),
    .A2_N(_06912_),
    .B1(_06932_),
    .B2(_06809_),
    .X(_06933_));
 sky130_fd_sc_hd__xnor2_1 _13763_ (.A(_06931_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__nor2_1 _13764_ (.A(_06802_),
    .B(_06762_),
    .Y(_06935_));
 sky130_fd_sc_hd__nor2_1 _13765_ (.A(_06783_),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__xnor2_1 _13766_ (.A(_06934_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__nand2_1 _13767_ (.A(_06930_),
    .B(_06937_),
    .Y(_06938_));
 sky130_fd_sc_hd__or2_1 _13768_ (.A(_06930_),
    .B(_06937_),
    .X(_06939_));
 sky130_fd_sc_hd__nand2_1 _13769_ (.A(_06938_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__xnor2_1 _13770_ (.A(_06926_),
    .B(_06940_),
    .Y(_06941_));
 sky130_fd_sc_hd__nor2_1 _13771_ (.A(_06830_),
    .B(_06854_),
    .Y(_06942_));
 sky130_fd_sc_hd__or3_1 _13772_ (.A(_06852_),
    .B(_06855_),
    .C(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__or2_1 _13773_ (.A(_06910_),
    .B(_06915_),
    .X(_06944_));
 sky130_fd_sc_hd__or2b_1 _13774_ (.A(_06916_),
    .B_N(_06909_),
    .X(_06945_));
 sky130_fd_sc_hd__nor2_1 _13775_ (.A(_06688_),
    .B(_06854_),
    .Y(_06946_));
 sky130_fd_sc_hd__xnor2_1 _13776_ (.A(_06858_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__xnor2_1 _13777_ (.A(_06859_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__a21o_1 _13778_ (.A1(_06944_),
    .A2(_06945_),
    .B1(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__nand3_1 _13779_ (.A(_06944_),
    .B(_06945_),
    .C(_06948_),
    .Y(_06950_));
 sky130_fd_sc_hd__nand2_1 _13780_ (.A(_06949_),
    .B(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__xor2_1 _13781_ (.A(_06943_),
    .B(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__xnor2_1 _13782_ (.A(_06941_),
    .B(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__a21o_1 _13783_ (.A1(_06919_),
    .A2(_06924_),
    .B1(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__nand3_1 _13784_ (.A(_06919_),
    .B(_06924_),
    .C(_06953_),
    .Y(_06955_));
 sky130_fd_sc_hd__and2_1 _13785_ (.A(_06954_),
    .B(_06955_),
    .X(_06956_));
 sky130_fd_sc_hd__xnor2_1 _13786_ (.A(_06869_),
    .B(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__or2_1 _13787_ (.A(_06864_),
    .B(_06851_),
    .X(_06958_));
 sky130_fd_sc_hd__o21ai_1 _13788_ (.A1(_06853_),
    .A2(_06851_),
    .B1(_06857_),
    .Y(_06959_));
 sky130_fd_sc_hd__a2bb2o_1 _13789_ (.A1_N(_06855_),
    .A2_N(_06958_),
    .B1(_06959_),
    .B2(_06856_),
    .X(_06960_));
 sky130_fd_sc_hd__and2_1 _13790_ (.A(_06866_),
    .B(_06960_),
    .X(_06961_));
 sky130_fd_sc_hd__o22ai_2 _13791_ (.A1(_06773_),
    .A2(_06817_),
    .B1(_06813_),
    .B2(_06816_),
    .Y(_06962_));
 sky130_fd_sc_hd__or4_1 _13792_ (.A(_06781_),
    .B(_06773_),
    .C(_06817_),
    .D(_06813_),
    .X(_06963_));
 sky130_fd_sc_hd__a21bo_1 _13793_ (.A1(_06832_),
    .A2(_06962_),
    .B1_N(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__nor2_1 _13794_ (.A(_06761_),
    .B(_06803_),
    .Y(_06965_));
 sky130_fd_sc_hd__xnor2_1 _13795_ (.A(_06965_),
    .B(_06806_),
    .Y(_06966_));
 sky130_fd_sc_hd__xnor2_1 _13796_ (.A(_06964_),
    .B(_06966_),
    .Y(_06967_));
 sky130_fd_sc_hd__inv_2 _13797_ (.A(_06853_),
    .Y(_06968_));
 sky130_fd_sc_hd__nand2_1 _13798_ (.A(_06968_),
    .B(_06911_),
    .Y(_06969_));
 sky130_fd_sc_hd__a21o_1 _13799_ (.A1(_06783_),
    .A2(_06784_),
    .B1(_06761_),
    .X(_06970_));
 sky130_fd_sc_hd__xnor2_1 _13800_ (.A(_06788_),
    .B(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__or2_1 _13801_ (.A(_06788_),
    .B(_06970_),
    .X(_06972_));
 sky130_fd_sc_hd__o21ai_1 _13802_ (.A1(_06969_),
    .A2(_06971_),
    .B1(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__or2b_1 _13803_ (.A(_06967_),
    .B_N(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__a21bo_1 _13804_ (.A1(_06964_),
    .A2(_06966_),
    .B1_N(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__clkbuf_4 _13805_ (.A(_06879_),
    .X(_06976_));
 sky130_fd_sc_hd__or2_1 _13806_ (.A(_06976_),
    .B(_06854_),
    .X(_06977_));
 sky130_fd_sc_hd__or3b_1 _13807_ (.A(_06958_),
    .B(_06977_),
    .C_N(_06855_),
    .X(_06978_));
 sky130_fd_sc_hd__xor2_1 _13808_ (.A(_06961_),
    .B(_06975_),
    .X(_06979_));
 sky130_fd_sc_hd__and2b_1 _13809_ (.A_N(_06978_),
    .B(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__a21o_1 _13810_ (.A1(_06961_),
    .A2(_06975_),
    .B1(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__xor2_1 _13811_ (.A(_06884_),
    .B(_06885_),
    .X(_06982_));
 sky130_fd_sc_hd__a21bo_1 _13812_ (.A1(_06801_),
    .A2(_06870_),
    .B1_N(_06880_),
    .X(_06983_));
 sky130_fd_sc_hd__nand2_1 _13813_ (.A(_06881_),
    .B(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__nor2_1 _13814_ (.A(_06816_),
    .B(_06877_),
    .Y(_06985_));
 sky130_fd_sc_hd__a21o_1 _13815_ (.A1(_06801_),
    .A2(_06872_),
    .B1(_06876_),
    .X(_06986_));
 sky130_fd_sc_hd__nand3_1 _13816_ (.A(_06802_),
    .B(_06872_),
    .C(_06876_),
    .Y(_06987_));
 sky130_fd_sc_hd__a21boi_1 _13817_ (.A1(_06985_),
    .A2(_06986_),
    .B1_N(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__xnor2_1 _13818_ (.A(_06984_),
    .B(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__and3_1 _13819_ (.A(_06832_),
    .B(_06963_),
    .C(_06962_),
    .X(_06990_));
 sky130_fd_sc_hd__a21oi_1 _13820_ (.A1(_06963_),
    .A2(_06962_),
    .B1(_06832_),
    .Y(_06991_));
 sky130_fd_sc_hd__nor3_1 _13821_ (.A(_06989_),
    .B(_06990_),
    .C(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__o21ba_1 _13822_ (.A1(_06984_),
    .A2(_06988_),
    .B1_N(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__xnor2_1 _13823_ (.A(_06982_),
    .B(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__xnor2_1 _13824_ (.A(_06973_),
    .B(_06967_),
    .Y(_06995_));
 sky130_fd_sc_hd__or2b_1 _13825_ (.A(_06993_),
    .B_N(_06982_),
    .X(_06996_));
 sky130_fd_sc_hd__a21bo_1 _13826_ (.A1(_06994_),
    .A2(_06995_),
    .B1_N(_06996_),
    .X(_06997_));
 sky130_fd_sc_hd__xnor2_1 _13827_ (.A(_06896_),
    .B(_06897_),
    .Y(_06998_));
 sky130_fd_sc_hd__xor2_1 _13828_ (.A(_06997_),
    .B(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__xor2_1 _13829_ (.A(_06978_),
    .B(_06979_),
    .X(_07000_));
 sky130_fd_sc_hd__and2b_1 _13830_ (.A_N(_06998_),
    .B(_06997_),
    .X(_07001_));
 sky130_fd_sc_hd__o21ba_1 _13831_ (.A1(_06999_),
    .A2(_07000_),
    .B1_N(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__xnor2_1 _13832_ (.A(_06921_),
    .B(_06923_),
    .Y(_07003_));
 sky130_fd_sc_hd__xnor2_1 _13833_ (.A(_07002_),
    .B(_07003_),
    .Y(_07004_));
 sky130_fd_sc_hd__or2b_1 _13834_ (.A(_07002_),
    .B_N(_07003_),
    .X(_07005_));
 sky130_fd_sc_hd__a21boi_1 _13835_ (.A1(_06981_),
    .A2(_07004_),
    .B1_N(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__xor2_1 _13836_ (.A(_06957_),
    .B(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__xnor2_1 _13837_ (.A(_06981_),
    .B(_07004_),
    .Y(_07008_));
 sky130_fd_sc_hd__nor2_1 _13838_ (.A(_06830_),
    .B(_06824_),
    .Y(_07009_));
 sky130_fd_sc_hd__nor4_1 _13839_ (.A(_06688_),
    .B(_06820_),
    .C(_06818_),
    .D(_06813_),
    .Y(_07010_));
 sky130_fd_sc_hd__o22a_1 _13840_ (.A1(_06688_),
    .A2(_06818_),
    .B1(_06813_),
    .B2(_06820_),
    .X(_07011_));
 sky130_fd_sc_hd__nor2_1 _13841_ (.A(_07010_),
    .B(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__a21oi_1 _13842_ (.A1(_07009_),
    .A2(_07012_),
    .B1(_07010_),
    .Y(_07013_));
 sky130_fd_sc_hd__xnor2_1 _13843_ (.A(_06969_),
    .B(_06971_),
    .Y(_07014_));
 sky130_fd_sc_hd__nand2_1 _13844_ (.A(_06863_),
    .B(_06912_),
    .Y(_07015_));
 sky130_fd_sc_hd__or2_1 _13845_ (.A(_06761_),
    .B(_06787_),
    .X(_07016_));
 sky130_fd_sc_hd__a21oi_1 _13846_ (.A1(_06783_),
    .A2(_06784_),
    .B1(_06853_),
    .Y(_07017_));
 sky130_fd_sc_hd__xnor2_1 _13847_ (.A(_07016_),
    .B(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__or2b_1 _13848_ (.A(_07015_),
    .B_N(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__o31a_1 _13849_ (.A1(_06853_),
    .A2(_06787_),
    .A3(_06970_),
    .B1(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__xor2_1 _13850_ (.A(_07013_),
    .B(_07014_),
    .X(_07021_));
 sky130_fd_sc_hd__and2b_1 _13851_ (.A_N(_07020_),
    .B(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__o21ba_1 _13852_ (.A1(_07013_),
    .A2(_07014_),
    .B1_N(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__or2_1 _13853_ (.A(_06958_),
    .B(_06977_),
    .X(_07024_));
 sky130_fd_sc_hd__xor2_1 _13854_ (.A(_06855_),
    .B(_06958_),
    .X(_07025_));
 sky130_fd_sc_hd__xnor2_1 _13855_ (.A(_07024_),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__and2b_1 _13856_ (.A_N(_07023_),
    .B(_07026_),
    .X(_07027_));
 sky130_fd_sc_hd__xnor2_1 _13857_ (.A(_06994_),
    .B(_06995_),
    .Y(_07028_));
 sky130_fd_sc_hd__o21a_1 _13858_ (.A1(_06990_),
    .A2(_06991_),
    .B1(_06989_),
    .X(_07029_));
 sky130_fd_sc_hd__or2_1 _13859_ (.A(_06992_),
    .B(_07029_),
    .X(_07030_));
 sky130_fd_sc_hd__and3_1 _13860_ (.A(_06987_),
    .B(_06985_),
    .C(_06986_),
    .X(_07031_));
 sky130_fd_sc_hd__a21oi_1 _13861_ (.A1(_06987_),
    .A2(_06986_),
    .B1(_06985_),
    .Y(_07032_));
 sky130_fd_sc_hd__nor2_1 _13862_ (.A(_07031_),
    .B(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__nor2_1 _13863_ (.A(_06820_),
    .B(_06877_),
    .Y(_07034_));
 sky130_fd_sc_hd__xnor2_2 _13864_ (.A(_06863_),
    .B(_06879_),
    .Y(_07035_));
 sky130_fd_sc_hd__a2bb2o_1 _13865_ (.A1_N(_06781_),
    .A2_N(_07035_),
    .B1(_06871_),
    .B2(_06801_),
    .X(_07036_));
 sky130_fd_sc_hd__nor2_1 _13866_ (.A(_06781_),
    .B(_06879_),
    .Y(_07037_));
 sky130_fd_sc_hd__and3_1 _13867_ (.A(_06801_),
    .B(_06872_),
    .C(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__a21o_1 _13868_ (.A1(_07034_),
    .A2(_07036_),
    .B1(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__xor2_1 _13869_ (.A(_07033_),
    .B(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__xor2_1 _13870_ (.A(_07009_),
    .B(_07012_),
    .X(_07041_));
 sky130_fd_sc_hd__and2_1 _13871_ (.A(_07033_),
    .B(_07039_),
    .X(_07042_));
 sky130_fd_sc_hd__a21o_1 _13872_ (.A1(_07040_),
    .A2(_07041_),
    .B1(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__xnor2_1 _13873_ (.A(_07030_),
    .B(_07043_),
    .Y(_07044_));
 sky130_fd_sc_hd__xnor2_1 _13874_ (.A(_07020_),
    .B(_07021_),
    .Y(_07045_));
 sky130_fd_sc_hd__or2b_1 _13875_ (.A(_07030_),
    .B_N(_07043_),
    .X(_07046_));
 sky130_fd_sc_hd__a21bo_1 _13876_ (.A1(_07044_),
    .A2(_07045_),
    .B1_N(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__and2b_1 _13877_ (.A_N(_07028_),
    .B(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__xor2_1 _13878_ (.A(_07047_),
    .B(_07028_),
    .X(_07049_));
 sky130_fd_sc_hd__xnor2_1 _13879_ (.A(_07023_),
    .B(_07026_),
    .Y(_07050_));
 sky130_fd_sc_hd__and2b_1 _13880_ (.A_N(_07049_),
    .B(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__nor2_1 _13881_ (.A(_07048_),
    .B(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__xor2_1 _13882_ (.A(_06999_),
    .B(_07000_),
    .X(_07053_));
 sky130_fd_sc_hd__xnor2_1 _13883_ (.A(_07052_),
    .B(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__and2b_1 _13884_ (.A_N(_07052_),
    .B(_07053_),
    .X(_07055_));
 sky130_fd_sc_hd__a21oi_1 _13885_ (.A1(_07027_),
    .A2(_07054_),
    .B1(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__nor2_1 _13886_ (.A(_07008_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__and2_1 _13887_ (.A(_07007_),
    .B(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__nand2_1 _13888_ (.A(_06869_),
    .B(_06956_),
    .Y(_07059_));
 sky130_fd_sc_hd__nand2_1 _13889_ (.A(_06954_),
    .B(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__o21a_1 _13890_ (.A1(_06943_),
    .A2(_06951_),
    .B1(_06949_),
    .X(_07061_));
 sky130_fd_sc_hd__a32o_1 _13891_ (.A1(_06926_),
    .A2(_06938_),
    .A3(_06939_),
    .B1(_06941_),
    .B2(_06952_),
    .X(_07062_));
 sky130_fd_sc_hd__inv_2 _13892_ (.A(_06839_),
    .Y(_07063_));
 sky130_fd_sc_hd__nor2_1 _13893_ (.A(_06816_),
    .B(_06803_),
    .Y(_07064_));
 sky130_fd_sc_hd__nand2_1 _13894_ (.A(_06850_),
    .B(_06932_),
    .Y(_07065_));
 sky130_fd_sc_hd__nand2_2 _13895_ (.A(_06783_),
    .B(_06784_),
    .Y(_07066_));
 sky130_fd_sc_hd__nand2_1 _13896_ (.A(_06802_),
    .B(_07066_),
    .Y(_07067_));
 sky130_fd_sc_hd__xor2_1 _13897_ (.A(_07065_),
    .B(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__xnor2_1 _13898_ (.A(_07064_),
    .B(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__xnor2_1 _13899_ (.A(_06928_),
    .B(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__xnor2_1 _13900_ (.A(_07063_),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__xnor2_1 _13901_ (.A(_06927_),
    .B(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__or2_1 _13902_ (.A(_06938_),
    .B(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__nand2_1 _13903_ (.A(_06938_),
    .B(_07072_),
    .Y(_07074_));
 sky130_fd_sc_hd__and2_1 _13904_ (.A(_07073_),
    .B(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__nand2_1 _13905_ (.A(_06859_),
    .B(_06947_),
    .Y(_07076_));
 sky130_fd_sc_hd__nand2_1 _13906_ (.A(_06931_),
    .B(_06933_),
    .Y(_07077_));
 sky130_fd_sc_hd__o31ai_2 _13907_ (.A1(_06783_),
    .A2(_06934_),
    .A3(_06935_),
    .B1(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__nor2_1 _13908_ (.A(_06820_),
    .B(_06854_),
    .Y(_07079_));
 sky130_fd_sc_hd__or2_1 _13909_ (.A(_06688_),
    .B(_06851_),
    .X(_07080_));
 sky130_fd_sc_hd__or3b_1 _13910_ (.A(_07079_),
    .B(_07080_),
    .C_N(_06942_),
    .X(_07081_));
 sky130_fd_sc_hd__inv_2 _13911_ (.A(_07080_),
    .Y(_07082_));
 sky130_fd_sc_hd__xnor2_1 _13912_ (.A(_07080_),
    .B(_07079_),
    .Y(_07083_));
 sky130_fd_sc_hd__a21o_1 _13913_ (.A1(_06942_),
    .A2(_07082_),
    .B1(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__and2_1 _13914_ (.A(_07081_),
    .B(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__xnor2_1 _13915_ (.A(_07078_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__nor2_1 _13916_ (.A(_07076_),
    .B(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__and2_1 _13917_ (.A(_07076_),
    .B(_07086_),
    .X(_07088_));
 sky130_fd_sc_hd__nor2_1 _13918_ (.A(_07087_),
    .B(_07088_),
    .Y(_07089_));
 sky130_fd_sc_hd__nand2_1 _13919_ (.A(_07075_),
    .B(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__or2_1 _13920_ (.A(_07075_),
    .B(_07089_),
    .X(_07091_));
 sky130_fd_sc_hd__nand2_1 _13921_ (.A(_07090_),
    .B(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__xnor2_1 _13922_ (.A(_07062_),
    .B(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__or2b_1 _13923_ (.A(_07061_),
    .B_N(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__or2b_1 _13924_ (.A(_07093_),
    .B_N(_07061_),
    .X(_07095_));
 sky130_fd_sc_hd__nand2_1 _13925_ (.A(_07094_),
    .B(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__xnor2_1 _13926_ (.A(_07060_),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__nor2_1 _13927_ (.A(_06957_),
    .B(_07006_),
    .Y(_07098_));
 sky130_fd_sc_hd__nor2_1 _13928_ (.A(_07098_),
    .B(_07058_),
    .Y(_07099_));
 sky130_fd_sc_hd__xnor2_1 _13929_ (.A(_07097_),
    .B(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__xnor2_2 _13930_ (.A(_07027_),
    .B(_07054_),
    .Y(_07101_));
 sky130_fd_sc_hd__xnor2_1 _13931_ (.A(_07040_),
    .B(_07041_),
    .Y(_07102_));
 sky130_fd_sc_hd__and2b_1 _13932_ (.A_N(_07038_),
    .B(_07036_),
    .X(_07103_));
 sky130_fd_sc_hd__xnor2_2 _13933_ (.A(_07034_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__or2_1 _13934_ (.A(_06687_),
    .B(_06877_),
    .X(_07105_));
 sky130_fd_sc_hd__or3b_1 _13935_ (.A(_06773_),
    .B(_07035_),
    .C_N(_07037_),
    .X(_07106_));
 sky130_fd_sc_hd__o21bai_1 _13936_ (.A1(_06773_),
    .A2(_07035_),
    .B1_N(_07037_),
    .Y(_07107_));
 sky130_fd_sc_hd__nand2_1 _13937_ (.A(_07106_),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__o21a_1 _13938_ (.A1(_07105_),
    .A2(_07108_),
    .B1(_07106_),
    .X(_07109_));
 sky130_fd_sc_hd__xnor2_1 _13939_ (.A(_07104_),
    .B(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__mux2_1 _13940_ (.A0(_06813_),
    .A1(_06789_),
    .S(_06688_),
    .X(_07111_));
 sky130_fd_sc_hd__o22ai_2 _13941_ (.A1(_07104_),
    .A2(_07109_),
    .B1(_07110_),
    .B2(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__xnor2_1 _13942_ (.A(_07102_),
    .B(_07112_),
    .Y(_07113_));
 sky130_fd_sc_hd__nor2_2 _13943_ (.A(_06853_),
    .B(_06787_),
    .Y(_07114_));
 sky130_fd_sc_hd__a21oi_4 _13944_ (.A1(_06783_),
    .A2(_06784_),
    .B1(_06864_),
    .Y(_07115_));
 sky130_fd_sc_hd__xor2_2 _13945_ (.A(_07114_),
    .B(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__a32oi_4 _13946_ (.A1(_06871_),
    .A2(_06912_),
    .A3(_07116_),
    .B1(_07115_),
    .B2(_07114_),
    .Y(_07117_));
 sky130_fd_sc_hd__xnor2_1 _13947_ (.A(_07015_),
    .B(_07018_),
    .Y(_07118_));
 sky130_fd_sc_hd__xnor2_1 _13948_ (.A(_06762_),
    .B(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__xnor2_1 _13949_ (.A(_07117_),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__or2b_1 _13950_ (.A(_07102_),
    .B_N(_07112_),
    .X(_07121_));
 sky130_fd_sc_hd__a21boi_1 _13951_ (.A1(_07113_),
    .A2(_07120_),
    .B1_N(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__xnor2_1 _13952_ (.A(_07044_),
    .B(_07045_),
    .Y(_07123_));
 sky130_fd_sc_hd__xor2_1 _13953_ (.A(_07122_),
    .B(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__nand2_1 _13954_ (.A(_06832_),
    .B(_07118_),
    .Y(_07125_));
 sky130_fd_sc_hd__or2b_1 _13955_ (.A(_07117_),
    .B_N(_07119_),
    .X(_07126_));
 sky130_fd_sc_hd__o21ai_1 _13956_ (.A1(_06976_),
    .A2(_06851_),
    .B1(_06865_),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_1 _13957_ (.A(_07024_),
    .B(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__a21oi_2 _13958_ (.A1(_07125_),
    .A2(_07126_),
    .B1(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__and3_1 _13959_ (.A(_07125_),
    .B(_07126_),
    .C(_07128_),
    .X(_07130_));
 sky130_fd_sc_hd__nor2_1 _13960_ (.A(_07129_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__nor2_1 _13961_ (.A(_07122_),
    .B(_07123_),
    .Y(_07132_));
 sky130_fd_sc_hd__a21o_1 _13962_ (.A1(_07124_),
    .A2(_07131_),
    .B1(_07132_),
    .X(_07133_));
 sky130_fd_sc_hd__xnor2_1 _13963_ (.A(_07049_),
    .B(_07050_),
    .Y(_07134_));
 sky130_fd_sc_hd__xor2_1 _13964_ (.A(_07133_),
    .B(_07134_),
    .X(_07135_));
 sky130_fd_sc_hd__and2_1 _13965_ (.A(_07129_),
    .B(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__a21oi_2 _13966_ (.A1(_07133_),
    .A2(_07134_),
    .B1(_07136_),
    .Y(_07137_));
 sky130_fd_sc_hd__nor2_1 _13967_ (.A(_07101_),
    .B(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__inv_2 _13968_ (.A(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__xnor2_1 _13969_ (.A(_07008_),
    .B(_07056_),
    .Y(_07140_));
 sky130_fd_sc_hd__nor2_1 _13970_ (.A(_07139_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__xnor2_1 _13971_ (.A(_07129_),
    .B(_07135_),
    .Y(_07142_));
 sky130_fd_sc_hd__clkbuf_4 _13972_ (.A(_06854_),
    .X(_07143_));
 sky130_fd_sc_hd__clkinv_2 _13973_ (.A(_07143_),
    .Y(_07144_));
 sky130_fd_sc_hd__nand2_1 _13974_ (.A(_06871_),
    .B(_06912_),
    .Y(_07145_));
 sky130_fd_sc_hd__xnor2_1 _13975_ (.A(_07145_),
    .B(_07116_),
    .Y(_07146_));
 sky130_fd_sc_hd__xor2_1 _13976_ (.A(_06823_),
    .B(_07146_),
    .X(_07147_));
 sky130_fd_sc_hd__nor2_1 _13977_ (.A(_06879_),
    .B(_06787_),
    .Y(_07148_));
 sky130_fd_sc_hd__and2_1 _13978_ (.A(_07115_),
    .B(_07148_),
    .X(_07149_));
 sky130_fd_sc_hd__and2b_1 _13979_ (.A_N(_07147_),
    .B(_07149_),
    .X(_07150_));
 sky130_fd_sc_hd__a31o_1 _13980_ (.A1(_06821_),
    .A2(_06822_),
    .A3(_07146_),
    .B1(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__and3_1 _13981_ (.A(_06871_),
    .B(_07144_),
    .C(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__xor2_1 _13982_ (.A(_07110_),
    .B(_07111_),
    .X(_07153_));
 sky130_fd_sc_hd__xnor2_1 _13983_ (.A(_07105_),
    .B(_07108_),
    .Y(_07154_));
 sky130_fd_sc_hd__nor2_1 _13984_ (.A(_06879_),
    .B(_06820_),
    .Y(_07155_));
 sky130_fd_sc_hd__nor2_1 _13985_ (.A(_06687_),
    .B(_07035_),
    .Y(_07156_));
 sky130_fd_sc_hd__nor2_1 _13986_ (.A(_06830_),
    .B(_06877_),
    .Y(_07157_));
 sky130_fd_sc_hd__xor2_1 _13987_ (.A(_07155_),
    .B(_07156_),
    .X(_07158_));
 sky130_fd_sc_hd__a22oi_2 _13988_ (.A1(_07155_),
    .A2(_07156_),
    .B1(_07157_),
    .B2(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__xnor2_1 _13989_ (.A(_07154_),
    .B(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__and2_1 _13990_ (.A(_06830_),
    .B(_06789_),
    .X(_07161_));
 sky130_fd_sc_hd__o32a_1 _13991_ (.A1(_06821_),
    .A2(_06822_),
    .A3(_07161_),
    .B1(_06824_),
    .B2(_06853_),
    .X(_07162_));
 sky130_fd_sc_hd__or2_1 _13992_ (.A(_07154_),
    .B(_07159_),
    .X(_07163_));
 sky130_fd_sc_hd__o21ai_1 _13993_ (.A1(_07160_),
    .A2(_07162_),
    .B1(_07163_),
    .Y(_07164_));
 sky130_fd_sc_hd__xor2_1 _13994_ (.A(_07153_),
    .B(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__xnor2_1 _13995_ (.A(_07147_),
    .B(_07149_),
    .Y(_07166_));
 sky130_fd_sc_hd__and2_1 _13996_ (.A(_07153_),
    .B(_07164_),
    .X(_07167_));
 sky130_fd_sc_hd__a21oi_1 _13997_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__xor2_1 _13998_ (.A(_07113_),
    .B(_07120_),
    .X(_07169_));
 sky130_fd_sc_hd__xnor2_1 _13999_ (.A(_07168_),
    .B(_07169_),
    .Y(_07170_));
 sky130_fd_sc_hd__xnor2_1 _14000_ (.A(_06977_),
    .B(_07151_),
    .Y(_07171_));
 sky130_fd_sc_hd__or2b_1 _14001_ (.A(_07168_),
    .B_N(_07169_),
    .X(_07172_));
 sky130_fd_sc_hd__a21boi_1 _14002_ (.A1(_07170_),
    .A2(_07171_),
    .B1_N(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__xnor2_1 _14003_ (.A(_07124_),
    .B(_07131_),
    .Y(_07174_));
 sky130_fd_sc_hd__xor2_1 _14004_ (.A(_07173_),
    .B(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__nor2_1 _14005_ (.A(_07173_),
    .B(_07174_),
    .Y(_07176_));
 sky130_fd_sc_hd__a21oi_1 _14006_ (.A1(_07152_),
    .A2(_07175_),
    .B1(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__nor2_1 _14007_ (.A(_07142_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__xor2_2 _14008_ (.A(_07101_),
    .B(_07137_),
    .X(_07179_));
 sky130_fd_sc_hd__nand2_1 _14009_ (.A(_07178_),
    .B(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__xnor2_1 _14010_ (.A(_07152_),
    .B(_07175_),
    .Y(_07181_));
 sky130_fd_sc_hd__xnor2_1 _14011_ (.A(_07157_),
    .B(_07158_),
    .Y(_07182_));
 sky130_fd_sc_hd__nor2_1 _14012_ (.A(_06879_),
    .B(_06688_),
    .Y(_07183_));
 sky130_fd_sc_hd__nor2_1 _14013_ (.A(_06750_),
    .B(_07035_),
    .Y(_07184_));
 sky130_fd_sc_hd__xnor2_1 _14014_ (.A(_07183_),
    .B(_07184_),
    .Y(_07185_));
 sky130_fd_sc_hd__nand2_1 _14015_ (.A(_07183_),
    .B(_07184_),
    .Y(_07186_));
 sky130_fd_sc_hd__o31a_1 _14016_ (.A1(_06789_),
    .A2(_06877_),
    .A3(_07185_),
    .B1(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__or2_1 _14017_ (.A(_07182_),
    .B(_07187_),
    .X(_07188_));
 sky130_fd_sc_hd__nor2_1 _14018_ (.A(_06864_),
    .B(_06824_),
    .Y(_07189_));
 sky130_fd_sc_hd__nor2_1 _14019_ (.A(_06726_),
    .B(_06789_),
    .Y(_07190_));
 sky130_fd_sc_hd__mux2_1 _14020_ (.A0(_06830_),
    .A1(_07190_),
    .S(_06853_),
    .X(_07191_));
 sky130_fd_sc_hd__xnor2_1 _14021_ (.A(_07189_),
    .B(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__xnor2_1 _14022_ (.A(_07182_),
    .B(_07187_),
    .Y(_07193_));
 sky130_fd_sc_hd__or2_1 _14023_ (.A(_07192_),
    .B(_07193_),
    .X(_07194_));
 sky130_fd_sc_hd__xnor2_1 _14024_ (.A(_07160_),
    .B(_07162_),
    .Y(_07195_));
 sky130_fd_sc_hd__a21o_1 _14025_ (.A1(_07188_),
    .A2(_07194_),
    .B1(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__o22a_1 _14026_ (.A1(_06879_),
    .A2(_06785_),
    .B1(_06787_),
    .B2(_06864_),
    .X(_07197_));
 sky130_fd_sc_hd__nor2_1 _14027_ (.A(_07149_),
    .B(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__a22o_1 _14028_ (.A1(_06968_),
    .A2(_06822_),
    .B1(_07189_),
    .B2(_07191_),
    .X(_07199_));
 sky130_fd_sc_hd__nand2_1 _14029_ (.A(_07198_),
    .B(_07199_),
    .Y(_07200_));
 sky130_fd_sc_hd__or2_1 _14030_ (.A(_07198_),
    .B(_07199_),
    .X(_07201_));
 sky130_fd_sc_hd__and2_1 _14031_ (.A(_07200_),
    .B(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__nand3_1 _14032_ (.A(_07195_),
    .B(_07188_),
    .C(_07194_),
    .Y(_07203_));
 sky130_fd_sc_hd__nand3_1 _14033_ (.A(_07196_),
    .B(_07202_),
    .C(_07203_),
    .Y(_07204_));
 sky130_fd_sc_hd__xnor2_1 _14034_ (.A(_07165_),
    .B(_07166_),
    .Y(_07205_));
 sky130_fd_sc_hd__a21oi_1 _14035_ (.A1(_07196_),
    .A2(_07204_),
    .B1(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__and3_1 _14036_ (.A(_07196_),
    .B(_07204_),
    .C(_07205_),
    .X(_07207_));
 sky130_fd_sc_hd__or2_1 _14037_ (.A(_07206_),
    .B(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__nor2_1 _14038_ (.A(_07200_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__xor2_1 _14039_ (.A(_07170_),
    .B(_07171_),
    .X(_07210_));
 sky130_fd_sc_hd__o21ai_1 _14040_ (.A1(_07206_),
    .A2(_07209_),
    .B1(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__nor2_1 _14041_ (.A(_07181_),
    .B(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__xor2_1 _14042_ (.A(_07142_),
    .B(_07177_),
    .X(_07213_));
 sky130_fd_sc_hd__and2_1 _14043_ (.A(_07212_),
    .B(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__xnor2_2 _14044_ (.A(_07212_),
    .B(_07213_),
    .Y(_07215_));
 sky130_fd_sc_hd__or3_1 _14045_ (.A(_07210_),
    .B(_07206_),
    .C(_07209_),
    .X(_07216_));
 sky130_fd_sc_hd__and3b_1 _14046_ (.A_N(_07181_),
    .B(_07211_),
    .C(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__and2_1 _14047_ (.A(_07200_),
    .B(_07208_),
    .X(_07218_));
 sky130_fd_sc_hd__nor2_1 _14048_ (.A(_07209_),
    .B(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__nor2_1 _14049_ (.A(_06853_),
    .B(_06789_),
    .Y(_07220_));
 sky130_fd_sc_hd__nor2_1 _14050_ (.A(_06864_),
    .B(_06818_),
    .Y(_07221_));
 sky130_fd_sc_hd__xor2_1 _14051_ (.A(_07220_),
    .B(_07221_),
    .X(_07222_));
 sky130_fd_sc_hd__clkbuf_4 _14052_ (.A(_06824_),
    .X(_07223_));
 sky130_fd_sc_hd__nor2_1 _14053_ (.A(_06976_),
    .B(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__a22o_1 _14054_ (.A1(_07220_),
    .A2(_07221_),
    .B1(_07222_),
    .B2(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__and2_1 _14055_ (.A(_07148_),
    .B(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__clkbuf_4 _14056_ (.A(_06877_),
    .X(_07227_));
 sky130_fd_sc_hd__nor2_1 _14057_ (.A(_06789_),
    .B(_07227_),
    .Y(_07228_));
 sky130_fd_sc_hd__xnor2_1 _14058_ (.A(_07228_),
    .B(_07185_),
    .Y(_07229_));
 sky130_fd_sc_hd__clkbuf_4 _14059_ (.A(_07035_),
    .X(_07230_));
 sky130_fd_sc_hd__o22ai_1 _14060_ (.A1(_06879_),
    .A2(_06830_),
    .B1(_06789_),
    .B2(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__and2_1 _14061_ (.A(_06810_),
    .B(_06822_),
    .X(_07232_));
 sky130_fd_sc_hd__a31o_1 _14062_ (.A1(_06726_),
    .A2(_06968_),
    .A3(_07231_),
    .B1(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__nand2_1 _14063_ (.A(_07229_),
    .B(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__xnor2_1 _14064_ (.A(_07222_),
    .B(_07224_),
    .Y(_07235_));
 sky130_fd_sc_hd__or2_1 _14065_ (.A(_07229_),
    .B(_07233_),
    .X(_07236_));
 sky130_fd_sc_hd__nand2_1 _14066_ (.A(_07234_),
    .B(_07236_),
    .Y(_07237_));
 sky130_fd_sc_hd__or2_1 _14067_ (.A(_07235_),
    .B(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__nand2_1 _14068_ (.A(_07192_),
    .B(_07193_),
    .Y(_07239_));
 sky130_fd_sc_hd__nand2_1 _14069_ (.A(_07194_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__a21oi_1 _14070_ (.A1(_07234_),
    .A2(_07238_),
    .B1(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__xnor2_1 _14071_ (.A(_07148_),
    .B(_07225_),
    .Y(_07242_));
 sky130_fd_sc_hd__and3_1 _14072_ (.A(_07240_),
    .B(_07234_),
    .C(_07238_),
    .X(_07243_));
 sky130_fd_sc_hd__or2_1 _14073_ (.A(_07241_),
    .B(_07243_),
    .X(_07244_));
 sky130_fd_sc_hd__nor2_1 _14074_ (.A(_07242_),
    .B(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__a21o_1 _14075_ (.A1(_07196_),
    .A2(_07203_),
    .B1(_07202_),
    .X(_07246_));
 sky130_fd_sc_hd__and2_1 _14076_ (.A(_07204_),
    .B(_07246_),
    .X(_07247_));
 sky130_fd_sc_hd__o21a_1 _14077_ (.A1(_07241_),
    .A2(_07245_),
    .B1(_07247_),
    .X(_07248_));
 sky130_fd_sc_hd__nor3_1 _14078_ (.A(_07247_),
    .B(_07241_),
    .C(_07245_),
    .Y(_07249_));
 sky130_fd_sc_hd__nor2_1 _14079_ (.A(_07248_),
    .B(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__a21o_1 _14080_ (.A1(_07226_),
    .A2(_07250_),
    .B1(_07248_),
    .X(_07251_));
 sky130_fd_sc_hd__nand3_2 _14081_ (.A(_07217_),
    .B(_07219_),
    .C(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__xor2_2 _14082_ (.A(_07215_),
    .B(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__and2_1 _14083_ (.A(_07242_),
    .B(_07244_),
    .X(_07254_));
 sky130_fd_sc_hd__or2_1 _14084_ (.A(_07245_),
    .B(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__nand2_1 _14085_ (.A(_07235_),
    .B(_07237_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand2_1 _14086_ (.A(_07238_),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__o22a_1 _14087_ (.A1(_06976_),
    .A2(_06818_),
    .B1(_06814_),
    .B2(_06864_),
    .X(_07258_));
 sky130_fd_sc_hd__a21oi_1 _14088_ (.A1(_06726_),
    .A2(_06968_),
    .B1(_07231_),
    .Y(_07259_));
 sky130_fd_sc_hd__or3_1 _14089_ (.A(_07233_),
    .B(_07258_),
    .C(_07259_),
    .X(_07260_));
 sky130_fd_sc_hd__o2bb2a_1 _14090_ (.A1_N(_06830_),
    .A2_N(_07190_),
    .B1(_07257_),
    .B2(_07260_),
    .X(_07261_));
 sky130_fd_sc_hd__a21oi_1 _14091_ (.A1(_06726_),
    .A2(_07255_),
    .B1(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__o21a_1 _14092_ (.A1(_07226_),
    .A2(_07250_),
    .B1(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__o211a_1 _14093_ (.A1(_07219_),
    .A2(_07251_),
    .B1(_07263_),
    .C1(_07217_),
    .X(_07264_));
 sky130_fd_sc_hd__nor2_1 _14094_ (.A(_07215_),
    .B(_07252_),
    .Y(_07265_));
 sky130_fd_sc_hd__a21o_1 _14095_ (.A1(_07253_),
    .A2(_07264_),
    .B1(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__nor2_1 _14096_ (.A(_07178_),
    .B(_07214_),
    .Y(_07267_));
 sky130_fd_sc_hd__xnor2_1 _14097_ (.A(_07179_),
    .B(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__a22o_1 _14098_ (.A1(_07179_),
    .A2(_07214_),
    .B1(_07266_),
    .B2(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__nand2_1 _14099_ (.A(_07139_),
    .B(_07180_),
    .Y(_07270_));
 sky130_fd_sc_hd__xnor2_1 _14100_ (.A(_07140_),
    .B(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__a2bb2o_1 _14101_ (.A1_N(_07140_),
    .A2_N(_07180_),
    .B1(_07269_),
    .B2(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__nor3_1 _14102_ (.A(_07007_),
    .B(_07057_),
    .C(_07141_),
    .Y(_07273_));
 sky130_fd_sc_hd__a211oi_1 _14103_ (.A1(_07007_),
    .A2(_07141_),
    .B1(_07273_),
    .C1(_07058_),
    .Y(_07274_));
 sky130_fd_sc_hd__a22o_1 _14104_ (.A1(_07007_),
    .A2(_07141_),
    .B1(_07272_),
    .B2(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__a22o_2 _14105_ (.A1(_07058_),
    .A2(_07097_),
    .B1(_07100_),
    .B2(_07275_),
    .X(_07276_));
 sky130_fd_sc_hd__nand2_1 _14106_ (.A(_07098_),
    .B(_07097_),
    .Y(_07277_));
 sky130_fd_sc_hd__a21oi_1 _14107_ (.A1(_06954_),
    .A2(_07059_),
    .B1(_07096_),
    .Y(_07278_));
 sky130_fd_sc_hd__or2b_1 _14108_ (.A(_07092_),
    .B_N(_07062_),
    .X(_07279_));
 sky130_fd_sc_hd__or2_1 _14109_ (.A(_06927_),
    .B(_07071_),
    .X(_07280_));
 sky130_fd_sc_hd__clkbuf_4 _14110_ (.A(_06787_),
    .X(_07281_));
 sky130_fd_sc_hd__nand2_1 _14111_ (.A(_06850_),
    .B(_07066_),
    .Y(_07282_));
 sky130_fd_sc_hd__nor2_1 _14112_ (.A(_07281_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__and2_1 _14113_ (.A(_07281_),
    .B(_07282_),
    .X(_07284_));
 sky130_fd_sc_hd__or2_1 _14114_ (.A(_07283_),
    .B(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__nor2_1 _14115_ (.A(_07280_),
    .B(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__and2_1 _14116_ (.A(_07280_),
    .B(_07285_),
    .X(_07287_));
 sky130_fd_sc_hd__or2_1 _14117_ (.A(_07286_),
    .B(_07287_),
    .X(_07288_));
 sky130_fd_sc_hd__or2_1 _14118_ (.A(_07063_),
    .B(_07070_),
    .X(_07289_));
 sky130_fd_sc_hd__o21ai_1 _14119_ (.A1(_06928_),
    .A2(_07069_),
    .B1(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__or2_1 _14120_ (.A(_06820_),
    .B(_06851_),
    .X(_07291_));
 sky130_fd_sc_hd__nor3_1 _14121_ (.A(_06816_),
    .B(_07143_),
    .C(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__or3b_1 _14122_ (.A(_07292_),
    .B(_07291_),
    .C_N(_06946_),
    .X(_07293_));
 sky130_fd_sc_hd__o21a_1 _14123_ (.A1(_06816_),
    .A2(_07143_),
    .B1(_07291_),
    .X(_07294_));
 sky130_fd_sc_hd__a2bb2o_1 _14124_ (.A1_N(_07292_),
    .A2_N(_07294_),
    .B1(_07082_),
    .B2(_07079_),
    .X(_07295_));
 sky130_fd_sc_hd__and2_1 _14125_ (.A(_07293_),
    .B(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__xnor2_1 _14126_ (.A(_07290_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__xnor2_1 _14127_ (.A(_07081_),
    .B(_07297_),
    .Y(_07298_));
 sky130_fd_sc_hd__xnor2_1 _14128_ (.A(_07288_),
    .B(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__a21oi_1 _14129_ (.A1(_07073_),
    .A2(_07090_),
    .B1(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__and3_1 _14130_ (.A(_07073_),
    .B(_07090_),
    .C(_07299_),
    .X(_07301_));
 sky130_fd_sc_hd__nor2_1 _14131_ (.A(_07300_),
    .B(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__a21oi_1 _14132_ (.A1(_07078_),
    .A2(_07085_),
    .B1(_07087_),
    .Y(_07303_));
 sky130_fd_sc_hd__xor2_1 _14133_ (.A(_07302_),
    .B(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__a21oi_2 _14134_ (.A1(_07279_),
    .A2(_07094_),
    .B1(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__and3_1 _14135_ (.A(_07279_),
    .B(_07094_),
    .C(_07304_),
    .X(_07306_));
 sky130_fd_sc_hd__nor2_1 _14136_ (.A(_07305_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__xor2_1 _14137_ (.A(_07278_),
    .B(_07307_),
    .X(_07308_));
 sky130_fd_sc_hd__xnor2_2 _14138_ (.A(_07277_),
    .B(_07308_),
    .Y(_07309_));
 sky130_fd_sc_hd__xnor2_2 _14139_ (.A(_07276_),
    .B(_07309_),
    .Y(_07310_));
 sky130_fd_sc_hd__xnor2_1 _14140_ (.A(_07272_),
    .B(_07274_),
    .Y(_07311_));
 sky130_fd_sc_hd__xor2_1 _14141_ (.A(_07269_),
    .B(_07271_),
    .X(_07312_));
 sky130_fd_sc_hd__xnor2_1 _14142_ (.A(_07266_),
    .B(_07268_),
    .Y(_07313_));
 sky130_fd_sc_hd__xnor2_2 _14143_ (.A(_07253_),
    .B(_07264_),
    .Y(_07314_));
 sky130_fd_sc_hd__nor2_1 _14144_ (.A(_07313_),
    .B(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__nor2_1 _14145_ (.A(_07312_),
    .B(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__nand2_1 _14146_ (.A(_07311_),
    .B(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__xor2_1 _14147_ (.A(_07275_),
    .B(_07100_),
    .X(_07318_));
 sky130_fd_sc_hd__nor2_1 _14148_ (.A(_07317_),
    .B(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__nand2_2 _14149_ (.A(_07310_),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__nand2_2 _14150_ (.A(_07278_),
    .B(_07307_),
    .Y(_07321_));
 sky130_fd_sc_hd__and2b_1 _14151_ (.A_N(_07303_),
    .B(_07302_),
    .X(_07322_));
 sky130_fd_sc_hd__nor2_1 _14152_ (.A(_07288_),
    .B(_07298_),
    .Y(_07323_));
 sky130_fd_sc_hd__nor2_1 _14153_ (.A(_07063_),
    .B(_07285_),
    .Y(_07324_));
 sky130_fd_sc_hd__a22o_1 _14154_ (.A1(_06850_),
    .A2(_06912_),
    .B1(_07066_),
    .B2(_06632_),
    .X(_07325_));
 sky130_fd_sc_hd__o31a_1 _14155_ (.A1(_06567_),
    .A2(_06803_),
    .A3(_07282_),
    .B1(_07325_),
    .X(_07326_));
 sky130_fd_sc_hd__o21a_1 _14156_ (.A1(_07283_),
    .A2(_07324_),
    .B1(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__nor3_1 _14157_ (.A(_07283_),
    .B(_07324_),
    .C(_07326_),
    .Y(_07328_));
 sky130_fd_sc_hd__nor2_1 _14158_ (.A(_07327_),
    .B(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__buf_2 _14159_ (.A(_06851_),
    .X(_07330_));
 sky130_fd_sc_hd__a2bb2o_1 _14160_ (.A1_N(_06816_),
    .A2_N(_07330_),
    .B1(_07144_),
    .B2(_06802_),
    .X(_07331_));
 sky130_fd_sc_hd__or4_1 _14161_ (.A(_06809_),
    .B(_06816_),
    .C(_07330_),
    .D(_07143_),
    .X(_07332_));
 sky130_fd_sc_hd__nand2_1 _14162_ (.A(_06839_),
    .B(_07285_),
    .Y(_07333_));
 sky130_fd_sc_hd__and4b_1 _14163_ (.A_N(_07292_),
    .B(_07331_),
    .C(_07332_),
    .D(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__xnor2_1 _14164_ (.A(_07293_),
    .B(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__nand2_1 _14165_ (.A(_07329_),
    .B(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__or2_1 _14166_ (.A(_07329_),
    .B(_07335_),
    .X(_07337_));
 sky130_fd_sc_hd__and2_1 _14167_ (.A(_07336_),
    .B(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__o21a_1 _14168_ (.A1(_07286_),
    .A2(_07323_),
    .B1(_07338_),
    .X(_07339_));
 sky130_fd_sc_hd__nor3_1 _14169_ (.A(_07286_),
    .B(_07323_),
    .C(_07338_),
    .Y(_07340_));
 sky130_fd_sc_hd__nor2_1 _14170_ (.A(_07339_),
    .B(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__nor2_1 _14171_ (.A(_07081_),
    .B(_07297_),
    .Y(_07342_));
 sky130_fd_sc_hd__a21oi_1 _14172_ (.A1(_07290_),
    .A2(_07296_),
    .B1(_07342_),
    .Y(_07343_));
 sky130_fd_sc_hd__xnor2_1 _14173_ (.A(_07341_),
    .B(_07343_),
    .Y(_07344_));
 sky130_fd_sc_hd__o21a_1 _14174_ (.A1(_07300_),
    .A2(_07322_),
    .B1(_07344_),
    .X(_07345_));
 sky130_fd_sc_hd__nor3_1 _14175_ (.A(_07300_),
    .B(_07322_),
    .C(_07344_),
    .Y(_07346_));
 sky130_fd_sc_hd__nor2_1 _14176_ (.A(_07345_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__xnor2_2 _14177_ (.A(_07305_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__xnor2_4 _14178_ (.A(_07321_),
    .B(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__or2b_1 _14179_ (.A(_07277_),
    .B_N(_07308_),
    .X(_07350_));
 sky130_fd_sc_hd__a21boi_2 _14180_ (.A1(_07276_),
    .A2(_07309_),
    .B1_N(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__xor2_4 _14181_ (.A(_07349_),
    .B(_07351_),
    .X(_07352_));
 sky130_fd_sc_hd__nand2_1 _14182_ (.A(_07276_),
    .B(_07309_),
    .Y(_07353_));
 sky130_fd_sc_hd__and2b_1 _14183_ (.A_N(_07343_),
    .B(_07341_),
    .X(_07354_));
 sky130_fd_sc_hd__and3_2 _14184_ (.A(_06802_),
    .B(_07327_),
    .C(_07332_),
    .X(_07355_));
 sky130_fd_sc_hd__a21oi_1 _14185_ (.A1(_06802_),
    .A2(_07332_),
    .B1(_07327_),
    .Y(_07356_));
 sky130_fd_sc_hd__nor2_1 _14186_ (.A(_07355_),
    .B(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__or2b_1 _14187_ (.A(_07293_),
    .B_N(_07334_),
    .X(_07358_));
 sky130_fd_sc_hd__o211a_1 _14188_ (.A1(_07292_),
    .A2(_07357_),
    .B1(_07358_),
    .C1(_07333_),
    .X(_07359_));
 sky130_fd_sc_hd__and3_1 _14189_ (.A(_06632_),
    .B(_06912_),
    .C(_07282_),
    .X(_07360_));
 sky130_fd_sc_hd__xnor2_1 _14190_ (.A(_07336_),
    .B(_07360_),
    .Y(_07361_));
 sky130_fd_sc_hd__xnor2_1 _14191_ (.A(_07359_),
    .B(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__or3_1 _14192_ (.A(_07339_),
    .B(_07354_),
    .C(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__o21a_1 _14193_ (.A1(_07065_),
    .A2(_07067_),
    .B1(_07363_),
    .X(_07364_));
 sky130_fd_sc_hd__xnor2_1 _14194_ (.A(_07345_),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__a21oi_1 _14195_ (.A1(_07321_),
    .A2(_07350_),
    .B1(_07348_),
    .Y(_07366_));
 sky130_fd_sc_hd__a21oi_1 _14196_ (.A1(_07305_),
    .A2(_07347_),
    .B1(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__o211a_1 _14197_ (.A1(_07353_),
    .A2(_07349_),
    .B1(_07365_),
    .C1(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__o21ba_2 _14198_ (.A1(_07320_),
    .A2(_07352_),
    .B1_N(_07368_),
    .X(_07369_));
 sky130_fd_sc_hd__buf_2 _14199_ (.A(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__buf_2 _14200_ (.A(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__xor2_4 _14201_ (.A(_07320_),
    .B(_07352_),
    .X(_07372_));
 sky130_fd_sc_hd__buf_2 _14202_ (.A(_07372_),
    .X(_07373_));
 sky130_fd_sc_hd__or2b_1 _14203_ (.A(_07330_),
    .B_N(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__and2_1 _14204_ (.A(_07144_),
    .B(_07371_),
    .X(_07375_));
 sky130_fd_sc_hd__nand2_1 _14205_ (.A(_07374_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__and2_1 _14206_ (.A(_06932_),
    .B(_07369_),
    .X(_07377_));
 sky130_fd_sc_hd__clkbuf_2 _14207_ (.A(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__nand2_1 _14208_ (.A(_07066_),
    .B(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__and2_1 _14209_ (.A(_06912_),
    .B(_07371_),
    .X(_07380_));
 sky130_fd_sc_hd__nand2_1 _14210_ (.A(_07066_),
    .B(_07370_),
    .Y(_07381_));
 sky130_fd_sc_hd__xnor2_2 _14211_ (.A(_07381_),
    .B(_07378_),
    .Y(_07382_));
 sky130_fd_sc_hd__nand2_1 _14212_ (.A(_07380_),
    .B(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__and3_1 _14213_ (.A(_06912_),
    .B(_07066_),
    .C(_07371_),
    .X(_07384_));
 sky130_fd_sc_hd__a21o_1 _14214_ (.A1(_07379_),
    .A2(_07383_),
    .B1(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__and3_1 _14215_ (.A(_07371_),
    .B(_07376_),
    .C(_07385_),
    .X(_07386_));
 sky130_fd_sc_hd__clkbuf_4 _14216_ (.A(_06785_),
    .X(_07387_));
 sky130_fd_sc_hd__or2_2 _14217_ (.A(_06567_),
    .B(_07369_),
    .X(_07388_));
 sky130_fd_sc_hd__o21ba_1 _14218_ (.A1(_07387_),
    .A2(_07388_),
    .B1_N(_07380_),
    .X(_07389_));
 sky130_fd_sc_hd__nor2_1 _14219_ (.A(_07384_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__nor2_1 _14220_ (.A(_07386_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__o21ai_1 _14221_ (.A1(_07281_),
    .A2(_07388_),
    .B1(_07381_),
    .Y(_07392_));
 sky130_fd_sc_hd__or2_1 _14222_ (.A(_07380_),
    .B(_07392_),
    .X(_07393_));
 sky130_fd_sc_hd__a21o_1 _14223_ (.A1(_07385_),
    .A2(_07393_),
    .B1(_06567_),
    .X(_07394_));
 sky130_fd_sc_hd__inv_2 _14224_ (.A(_07355_),
    .Y(_07395_));
 sky130_fd_sc_hd__xnor2_2 _14225_ (.A(_07310_),
    .B(_07319_),
    .Y(_07396_));
 sky130_fd_sc_hd__buf_2 _14226_ (.A(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__a21o_1 _14227_ (.A1(_07375_),
    .A2(_07397_),
    .B1(_07374_),
    .X(_07398_));
 sky130_fd_sc_hd__a21boi_1 _14228_ (.A1(_07395_),
    .A2(_07398_),
    .B1_N(_07376_),
    .Y(_07399_));
 sky130_fd_sc_hd__nand2_1 _14229_ (.A(_07394_),
    .B(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__a21oi_1 _14230_ (.A1(_07386_),
    .A2(_07390_),
    .B1(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__o21a_1 _14231_ (.A1(_07391_),
    .A2(_07401_),
    .B1(_07376_),
    .X(_07402_));
 sky130_fd_sc_hd__and2_1 _14232_ (.A(_07317_),
    .B(_07318_),
    .X(_07403_));
 sky130_fd_sc_hd__or2_1 _14233_ (.A(_07319_),
    .B(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__clkbuf_4 _14234_ (.A(_07404_),
    .X(_07405_));
 sky130_fd_sc_hd__or2_1 _14235_ (.A(_07143_),
    .B(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__or2_1 _14236_ (.A(_07311_),
    .B(_07316_),
    .X(_07407_));
 sky130_fd_sc_hd__nand2_2 _14237_ (.A(_07317_),
    .B(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__clkbuf_4 _14238_ (.A(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__or2_1 _14239_ (.A(_07330_),
    .B(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__nor2_1 _14240_ (.A(_07406_),
    .B(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__or2_1 _14241_ (.A(_07330_),
    .B(_07405_),
    .X(_07412_));
 sky130_fd_sc_hd__nor2_1 _14242_ (.A(_07143_),
    .B(_07397_),
    .Y(_07413_));
 sky130_fd_sc_hd__xnor2_1 _14243_ (.A(_07412_),
    .B(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__or2b_1 _14244_ (.A(_06818_),
    .B_N(_07369_),
    .X(_07415_));
 sky130_fd_sc_hd__o21ai_1 _14245_ (.A1(_06814_),
    .A2(_07388_),
    .B1(_07415_),
    .Y(_07416_));
 sky130_fd_sc_hd__and3_1 _14246_ (.A(_06903_),
    .B(_07371_),
    .C(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__and2_1 _14247_ (.A(_06912_),
    .B(_07373_),
    .X(_07418_));
 sky130_fd_sc_hd__xor2_1 _14248_ (.A(_07382_),
    .B(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__nand2_1 _14249_ (.A(_07417_),
    .B(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__or2_1 _14250_ (.A(_07417_),
    .B(_07419_),
    .X(_07421_));
 sky130_fd_sc_hd__nand2_1 _14251_ (.A(_07420_),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__buf_2 _14252_ (.A(_06803_),
    .X(_07423_));
 sky130_fd_sc_hd__nor2_1 _14253_ (.A(_07423_),
    .B(_07397_),
    .Y(_07424_));
 sky130_fd_sc_hd__and2_1 _14254_ (.A(_07066_),
    .B(_07373_),
    .X(_07425_));
 sky130_fd_sc_hd__xor2_1 _14255_ (.A(_07378_),
    .B(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__nand2_1 _14256_ (.A(_07378_),
    .B(_07425_),
    .Y(_07427_));
 sky130_fd_sc_hd__a21boi_1 _14257_ (.A1(_07424_),
    .A2(_07426_),
    .B1_N(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__o21ai_1 _14258_ (.A1(_07422_),
    .A2(_07428_),
    .B1(_07420_),
    .Y(_07429_));
 sky130_fd_sc_hd__nand2_1 _14259_ (.A(_07144_),
    .B(_07373_),
    .Y(_07430_));
 sky130_fd_sc_hd__or3b_1 _14260_ (.A(_07330_),
    .B(_07397_),
    .C_N(_07406_),
    .X(_07431_));
 sky130_fd_sc_hd__xnor2_1 _14261_ (.A(_07430_),
    .B(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__xnor2_1 _14262_ (.A(_07429_),
    .B(_07432_),
    .Y(_07433_));
 sky130_fd_sc_hd__inv_2 _14263_ (.A(_07432_),
    .Y(_07434_));
 sky130_fd_sc_hd__a32o_1 _14264_ (.A1(_07411_),
    .A2(_07414_),
    .A3(_07433_),
    .B1(_07434_),
    .B2(_07429_),
    .X(_07435_));
 sky130_fd_sc_hd__or2_1 _14265_ (.A(_07394_),
    .B(_07399_),
    .X(_07436_));
 sky130_fd_sc_hd__nand2_1 _14266_ (.A(_07400_),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__nand2_1 _14267_ (.A(_07411_),
    .B(_07414_),
    .Y(_07438_));
 sky130_fd_sc_hd__xnor2_1 _14268_ (.A(_07438_),
    .B(_07433_),
    .Y(_07439_));
 sky130_fd_sc_hd__clkbuf_4 _14269_ (.A(_06818_),
    .X(_07440_));
 sky130_fd_sc_hd__nand2_1 _14270_ (.A(_06903_),
    .B(_07370_),
    .Y(_07441_));
 sky130_fd_sc_hd__o21ai_1 _14271_ (.A1(_07440_),
    .A2(_07371_),
    .B1(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__xor2_1 _14272_ (.A(_07422_),
    .B(_07428_),
    .X(_07443_));
 sky130_fd_sc_hd__nand2_1 _14273_ (.A(_07442_),
    .B(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__nand2_1 _14274_ (.A(_07382_),
    .B(_07418_),
    .Y(_07445_));
 sky130_fd_sc_hd__or2_1 _14275_ (.A(_07380_),
    .B(_07382_),
    .X(_07446_));
 sky130_fd_sc_hd__nand2_1 _14276_ (.A(_07383_),
    .B(_07446_),
    .Y(_07447_));
 sky130_fd_sc_hd__a31o_1 _14277_ (.A1(_07379_),
    .A2(_07445_),
    .A3(_07447_),
    .B1(_07355_),
    .X(_07448_));
 sky130_fd_sc_hd__o21a_1 _14278_ (.A1(_07223_),
    .A2(_07371_),
    .B1(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__xor2_1 _14279_ (.A(_07444_),
    .B(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__nor2_1 _14280_ (.A(_07444_),
    .B(_07449_),
    .Y(_07451_));
 sky130_fd_sc_hd__a21oi_1 _14281_ (.A1(_07439_),
    .A2(_07450_),
    .B1(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__nand2_1 _14282_ (.A(_07437_),
    .B(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__nor2_1 _14283_ (.A(_07437_),
    .B(_07452_),
    .Y(_07454_));
 sky130_fd_sc_hd__a21oi_1 _14284_ (.A1(_07435_),
    .A2(_07453_),
    .B1(_07454_),
    .Y(_07455_));
 sky130_fd_sc_hd__nor2_1 _14285_ (.A(_07402_),
    .B(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__o21ai_1 _14286_ (.A1(_07423_),
    .A2(_07387_),
    .B1(_07371_),
    .Y(_07457_));
 sky130_fd_sc_hd__or2_1 _14287_ (.A(_07423_),
    .B(_07371_),
    .X(_07458_));
 sky130_fd_sc_hd__a21bo_1 _14288_ (.A1(_07386_),
    .A2(_07390_),
    .B1_N(_07385_),
    .X(_07459_));
 sky130_fd_sc_hd__a21o_1 _14289_ (.A1(_07457_),
    .A2(_07458_),
    .B1(_07459_),
    .X(_07460_));
 sky130_fd_sc_hd__xnor2_1 _14290_ (.A(_07401_),
    .B(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__nand2_2 _14291_ (.A(_07456_),
    .B(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__mux2_1 _14292_ (.A0(_07423_),
    .A1(_07144_),
    .S(_07371_),
    .X(_07463_));
 sky130_fd_sc_hd__nor2_1 _14293_ (.A(_07384_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__a2bb2o_1 _14294_ (.A1_N(_07400_),
    .A2_N(_07460_),
    .B1(_07464_),
    .B2(_07459_),
    .X(_07465_));
 sky130_fd_sc_hd__o21ba_2 _14295_ (.A1(_07459_),
    .A2(_07464_),
    .B1_N(_07465_),
    .X(_07466_));
 sky130_fd_sc_hd__xnor2_4 _14296_ (.A(_07462_),
    .B(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__and2b_1 _14297_ (.A_N(_07454_),
    .B(_07453_),
    .X(_07468_));
 sky130_fd_sc_hd__xnor2_1 _14298_ (.A(_07435_),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__and2_1 _14299_ (.A(_07312_),
    .B(_07315_),
    .X(_07470_));
 sky130_fd_sc_hd__or2_2 _14300_ (.A(_07316_),
    .B(_07470_),
    .X(_07471_));
 sky130_fd_sc_hd__clkbuf_4 _14301_ (.A(_07471_),
    .X(_07472_));
 sky130_fd_sc_hd__or2_1 _14302_ (.A(_07143_),
    .B(_07472_),
    .X(_07473_));
 sky130_fd_sc_hd__nor2_1 _14303_ (.A(_07410_),
    .B(_07473_),
    .Y(_07474_));
 sky130_fd_sc_hd__and2_1 _14304_ (.A(_07406_),
    .B(_07410_),
    .X(_07475_));
 sky130_fd_sc_hd__nor2_1 _14305_ (.A(_07411_),
    .B(_07475_),
    .Y(_07476_));
 sky130_fd_sc_hd__xnor2_1 _14306_ (.A(_07411_),
    .B(_07414_),
    .Y(_07477_));
 sky130_fd_sc_hd__or2_1 _14307_ (.A(_07423_),
    .B(_07405_),
    .X(_07478_));
 sky130_fd_sc_hd__o2bb2a_1 _14308_ (.A1_N(_06932_),
    .A2_N(_07373_),
    .B1(_07397_),
    .B2(_07387_),
    .X(_07479_));
 sky130_fd_sc_hd__nor2_1 _14309_ (.A(_07478_),
    .B(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__or3b_1 _14310_ (.A(_07440_),
    .B(_06814_),
    .C_N(_07370_),
    .X(_07481_));
 sky130_fd_sc_hd__and2_1 _14311_ (.A(_06826_),
    .B(_07369_),
    .X(_07482_));
 sky130_fd_sc_hd__xnor2_2 _14312_ (.A(_07415_),
    .B(_07482_),
    .Y(_07483_));
 sky130_fd_sc_hd__or2b_1 _14313_ (.A(_07441_),
    .B_N(_07483_),
    .X(_07484_));
 sky130_fd_sc_hd__xnor2_1 _14314_ (.A(_07424_),
    .B(_07426_),
    .Y(_07485_));
 sky130_fd_sc_hd__a21oi_1 _14315_ (.A1(_07481_),
    .A2(_07484_),
    .B1(_07485_),
    .Y(_07486_));
 sky130_fd_sc_hd__and3_1 _14316_ (.A(_07481_),
    .B(_07484_),
    .C(_07485_),
    .X(_07487_));
 sky130_fd_sc_hd__nor2_1 _14317_ (.A(_07486_),
    .B(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__a21oi_1 _14318_ (.A1(_07480_),
    .A2(_07488_),
    .B1(_07486_),
    .Y(_07489_));
 sky130_fd_sc_hd__nor2_1 _14319_ (.A(_07477_),
    .B(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__and2_1 _14320_ (.A(_07477_),
    .B(_07489_),
    .X(_07491_));
 sky130_fd_sc_hd__nor2_1 _14321_ (.A(_07490_),
    .B(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__a31o_1 _14322_ (.A1(_07474_),
    .A2(_07476_),
    .A3(_07492_),
    .B1(_07490_),
    .X(_07493_));
 sky130_fd_sc_hd__xnor2_1 _14323_ (.A(_07439_),
    .B(_07450_),
    .Y(_07494_));
 sky130_fd_sc_hd__nand2_1 _14324_ (.A(_07474_),
    .B(_07476_),
    .Y(_07495_));
 sky130_fd_sc_hd__xnor2_1 _14325_ (.A(_07495_),
    .B(_07492_),
    .Y(_07496_));
 sky130_fd_sc_hd__and2b_1 _14326_ (.A_N(_07416_),
    .B(_07441_),
    .X(_07497_));
 sky130_fd_sc_hd__nor2_1 _14327_ (.A(_07417_),
    .B(_07497_),
    .Y(_07498_));
 sky130_fd_sc_hd__xor2_2 _14328_ (.A(_07480_),
    .B(_07488_),
    .X(_07499_));
 sky130_fd_sc_hd__xor2_1 _14329_ (.A(_07442_),
    .B(_07443_),
    .X(_07500_));
 sky130_fd_sc_hd__and3_1 _14330_ (.A(_07498_),
    .B(_07499_),
    .C(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__a21oi_1 _14331_ (.A1(_07498_),
    .A2(_07499_),
    .B1(_07500_),
    .Y(_07502_));
 sky130_fd_sc_hd__nor2_1 _14332_ (.A(_07501_),
    .B(_07502_),
    .Y(_07503_));
 sky130_fd_sc_hd__a21oi_1 _14333_ (.A1(_07496_),
    .A2(_07503_),
    .B1(_07501_),
    .Y(_07504_));
 sky130_fd_sc_hd__nand2_1 _14334_ (.A(_07494_),
    .B(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__nor2_1 _14335_ (.A(_07494_),
    .B(_07504_),
    .Y(_07506_));
 sky130_fd_sc_hd__a21oi_1 _14336_ (.A1(_07493_),
    .A2(_07505_),
    .B1(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__nor2_1 _14337_ (.A(_07469_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__and2_1 _14338_ (.A(_07402_),
    .B(_07455_),
    .X(_07509_));
 sky130_fd_sc_hd__nor2_1 _14339_ (.A(_07456_),
    .B(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__and2_1 _14340_ (.A(_07508_),
    .B(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__or2_1 _14341_ (.A(_07456_),
    .B(_07461_),
    .X(_07512_));
 sky130_fd_sc_hd__and2_1 _14342_ (.A(_07462_),
    .B(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__nand2_1 _14343_ (.A(_07511_),
    .B(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__or2_1 _14344_ (.A(_07511_),
    .B(_07513_),
    .X(_07515_));
 sky130_fd_sc_hd__and2_1 _14345_ (.A(_07514_),
    .B(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__inv_2 _14346_ (.A(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__and2b_1 _14347_ (.A_N(_07506_),
    .B(_07505_),
    .X(_07518_));
 sky130_fd_sc_hd__xnor2_1 _14348_ (.A(_07493_),
    .B(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__xnor2_1 _14349_ (.A(_07496_),
    .B(_07503_),
    .Y(_07520_));
 sky130_fd_sc_hd__and2_1 _14350_ (.A(_07313_),
    .B(_07314_),
    .X(_07521_));
 sky130_fd_sc_hd__nor2_1 _14351_ (.A(_07315_),
    .B(_07521_),
    .Y(_07522_));
 sky130_fd_sc_hd__buf_2 _14352_ (.A(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__or2_1 _14353_ (.A(_07330_),
    .B(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__or2_1 _14354_ (.A(_07473_),
    .B(_07524_),
    .X(_07525_));
 sky130_fd_sc_hd__o22a_1 _14355_ (.A1(_07143_),
    .A2(_07409_),
    .B1(_07472_),
    .B2(_07330_),
    .X(_07526_));
 sky130_fd_sc_hd__o21a_1 _14356_ (.A1(_07474_),
    .A2(_07526_),
    .B1(_06632_),
    .X(_07527_));
 sky130_fd_sc_hd__or2_1 _14357_ (.A(_07525_),
    .B(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__xnor2_1 _14358_ (.A(_07474_),
    .B(_07476_),
    .Y(_07529_));
 sky130_fd_sc_hd__and2_1 _14359_ (.A(_06903_),
    .B(_07373_),
    .X(_07530_));
 sky130_fd_sc_hd__nand2_1 _14360_ (.A(_07483_),
    .B(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__and2_1 _14361_ (.A(_07478_),
    .B(_07479_),
    .X(_07532_));
 sky130_fd_sc_hd__or2_1 _14362_ (.A(_07480_),
    .B(_07532_),
    .X(_07533_));
 sky130_fd_sc_hd__a21o_1 _14363_ (.A1(_07481_),
    .A2(_07531_),
    .B1(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__nand3_1 _14364_ (.A(_07481_),
    .B(_07531_),
    .C(_07533_),
    .Y(_07535_));
 sky130_fd_sc_hd__nand2_1 _14365_ (.A(_07534_),
    .B(_07535_),
    .Y(_07536_));
 sky130_fd_sc_hd__or2_1 _14366_ (.A(_07387_),
    .B(_07404_),
    .X(_07537_));
 sky130_fd_sc_hd__nor2_1 _14367_ (.A(_07281_),
    .B(_07396_),
    .Y(_07538_));
 sky130_fd_sc_hd__xnor2_1 _14368_ (.A(_07537_),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__or3b_1 _14369_ (.A(_06803_),
    .B(_07409_),
    .C_N(_07539_),
    .X(_07540_));
 sky130_fd_sc_hd__o31a_1 _14370_ (.A1(_07281_),
    .A2(_07397_),
    .A3(_07537_),
    .B1(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__o21a_1 _14371_ (.A1(_07536_),
    .A2(_07541_),
    .B1(_07534_),
    .X(_07542_));
 sky130_fd_sc_hd__xor2_1 _14372_ (.A(_07529_),
    .B(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__xnor2_1 _14373_ (.A(_07528_),
    .B(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__xnor2_1 _14374_ (.A(_07498_),
    .B(_07499_),
    .Y(_07545_));
 sky130_fd_sc_hd__xor2_1 _14375_ (.A(_07536_),
    .B(_07541_),
    .X(_07546_));
 sky130_fd_sc_hd__xor2_1 _14376_ (.A(_07441_),
    .B(_07483_),
    .X(_07547_));
 sky130_fd_sc_hd__o211a_1 _14377_ (.A1(_07227_),
    .A2(_07388_),
    .B1(_07547_),
    .C1(_06632_),
    .X(_07548_));
 sky130_fd_sc_hd__xnor2_1 _14378_ (.A(_07483_),
    .B(_07530_),
    .Y(_07549_));
 sky130_fd_sc_hd__nand2_1 _14379_ (.A(_06870_),
    .B(_07370_),
    .Y(_07550_));
 sky130_fd_sc_hd__or2_1 _14380_ (.A(_07230_),
    .B(_07388_),
    .X(_07551_));
 sky130_fd_sc_hd__or3b_1 _14381_ (.A(_07227_),
    .B(_07230_),
    .C_N(_07369_),
    .X(_07552_));
 sky130_fd_sc_hd__a21bo_1 _14382_ (.A1(_07550_),
    .A2(_07551_),
    .B1_N(_07552_),
    .X(_07553_));
 sky130_fd_sc_hd__o21a_1 _14383_ (.A1(_07549_),
    .A2(_07553_),
    .B1(_07552_),
    .X(_07554_));
 sky130_fd_sc_hd__nand2_1 _14384_ (.A(_07548_),
    .B(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__nor2_1 _14385_ (.A(_07548_),
    .B(_07554_),
    .Y(_07556_));
 sky130_fd_sc_hd__a21oi_2 _14386_ (.A1(_07546_),
    .A2(_07555_),
    .B1(_07556_),
    .Y(_07557_));
 sky130_fd_sc_hd__xor2_1 _14387_ (.A(_07545_),
    .B(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__nor2_1 _14388_ (.A(_07545_),
    .B(_07557_),
    .Y(_07559_));
 sky130_fd_sc_hd__a21oi_1 _14389_ (.A1(_07544_),
    .A2(_07558_),
    .B1(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__xnor2_1 _14390_ (.A(_07520_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__or2b_1 _14391_ (.A(_07528_),
    .B_N(_07543_),
    .X(_07562_));
 sky130_fd_sc_hd__o21ai_1 _14392_ (.A1(_07529_),
    .A2(_07542_),
    .B1(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__or2b_1 _14393_ (.A(_07561_),
    .B_N(_07563_),
    .X(_07564_));
 sky130_fd_sc_hd__o21a_1 _14394_ (.A1(_07520_),
    .A2(_07560_),
    .B1(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__nor2_1 _14395_ (.A(_07519_),
    .B(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__and2_1 _14396_ (.A(_07469_),
    .B(_07507_),
    .X(_07567_));
 sky130_fd_sc_hd__nor2_1 _14397_ (.A(_07508_),
    .B(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__and2_1 _14398_ (.A(_07566_),
    .B(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__nor2_1 _14399_ (.A(_07566_),
    .B(_07568_),
    .Y(_07570_));
 sky130_fd_sc_hd__or2_1 _14400_ (.A(_07569_),
    .B(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__xor2_1 _14401_ (.A(_07563_),
    .B(_07561_),
    .X(_07572_));
 sky130_fd_sc_hd__buf_2 _14402_ (.A(_07314_),
    .X(_07573_));
 sky130_fd_sc_hd__or2_1 _14403_ (.A(_07143_),
    .B(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__nor2_2 _14404_ (.A(_07524_),
    .B(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__nand2_1 _14405_ (.A(_07473_),
    .B(_07524_),
    .Y(_07576_));
 sky130_fd_sc_hd__and2_1 _14406_ (.A(_07525_),
    .B(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__nand2_1 _14407_ (.A(_07525_),
    .B(_07527_),
    .Y(_07578_));
 sky130_fd_sc_hd__nand2_1 _14408_ (.A(_07528_),
    .B(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__and2b_1 _14409_ (.A_N(_07440_),
    .B(_07372_),
    .X(_07580_));
 sky130_fd_sc_hd__xnor2_1 _14410_ (.A(_07482_),
    .B(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__or2_1 _14411_ (.A(_07223_),
    .B(_07397_),
    .X(_07582_));
 sky130_fd_sc_hd__and2_1 _14412_ (.A(_07482_),
    .B(_07580_),
    .X(_07583_));
 sky130_fd_sc_hd__o21bai_2 _14413_ (.A1(_07581_),
    .A2(_07582_),
    .B1_N(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__o21bai_1 _14414_ (.A1(_07423_),
    .A2(_07409_),
    .B1_N(_07539_),
    .Y(_07585_));
 sky130_fd_sc_hd__and2_1 _14415_ (.A(_07540_),
    .B(_07585_),
    .X(_07586_));
 sky130_fd_sc_hd__xnor2_2 _14416_ (.A(_07584_),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__or2_1 _14417_ (.A(_07423_),
    .B(_07471_),
    .X(_07588_));
 sky130_fd_sc_hd__nor2_1 _14418_ (.A(_07281_),
    .B(_07405_),
    .Y(_07589_));
 sky130_fd_sc_hd__nor2_1 _14419_ (.A(_07387_),
    .B(_07408_),
    .Y(_07590_));
 sky130_fd_sc_hd__xnor2_1 _14420_ (.A(_07589_),
    .B(_07590_),
    .Y(_07591_));
 sky130_fd_sc_hd__nand2_1 _14421_ (.A(_07589_),
    .B(_07590_),
    .Y(_07592_));
 sky130_fd_sc_hd__o21a_1 _14422_ (.A1(_07588_),
    .A2(_07591_),
    .B1(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__nor2_1 _14423_ (.A(_07587_),
    .B(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__a21oi_1 _14424_ (.A1(_07584_),
    .A2(_07586_),
    .B1(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__xor2_1 _14425_ (.A(_07579_),
    .B(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__nor2_1 _14426_ (.A(_07579_),
    .B(_07595_),
    .Y(_07597_));
 sky130_fd_sc_hd__a31o_1 _14427_ (.A1(_07575_),
    .A2(_07577_),
    .A3(_07596_),
    .B1(_07597_),
    .X(_07598_));
 sky130_fd_sc_hd__xnor2_1 _14428_ (.A(_07544_),
    .B(_07558_),
    .Y(_07599_));
 sky130_fd_sc_hd__nand2_1 _14429_ (.A(_07575_),
    .B(_07577_),
    .Y(_07600_));
 sky130_fd_sc_hd__xnor2_1 _14430_ (.A(_07600_),
    .B(_07596_),
    .Y(_07601_));
 sky130_fd_sc_hd__and2b_1 _14431_ (.A_N(_07556_),
    .B(_07555_),
    .X(_07602_));
 sky130_fd_sc_hd__xnor2_1 _14432_ (.A(_07546_),
    .B(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__xor2_2 _14433_ (.A(_07587_),
    .B(_07593_),
    .X(_07604_));
 sky130_fd_sc_hd__xnor2_1 _14434_ (.A(_07549_),
    .B(_07553_),
    .Y(_07605_));
 sky130_fd_sc_hd__xor2_1 _14435_ (.A(_07581_),
    .B(_07582_),
    .X(_07606_));
 sky130_fd_sc_hd__o2bb2a_1 _14436_ (.A1_N(_06872_),
    .A2_N(_07370_),
    .B1(_07388_),
    .B2(_06976_),
    .X(_07607_));
 sky130_fd_sc_hd__nand2_1 _14437_ (.A(_06810_),
    .B(_07369_),
    .Y(_07608_));
 sky130_fd_sc_hd__or3b_1 _14438_ (.A(_06863_),
    .B(_07227_),
    .C_N(_07369_),
    .X(_07609_));
 sky130_fd_sc_hd__a21bo_1 _14439_ (.A1(_07608_),
    .A2(_07609_),
    .B1_N(_07552_),
    .X(_07610_));
 sky130_fd_sc_hd__a21boi_1 _14440_ (.A1(_07550_),
    .A2(_07607_),
    .B1_N(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__a21bo_1 _14441_ (.A1(_07606_),
    .A2(_07611_),
    .B1_N(_07610_),
    .X(_07612_));
 sky130_fd_sc_hd__xnor2_1 _14442_ (.A(_07605_),
    .B(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__and2b_1 _14443_ (.A_N(_07605_),
    .B(_07612_),
    .X(_07614_));
 sky130_fd_sc_hd__a21oi_1 _14444_ (.A1(_07604_),
    .A2(_07613_),
    .B1(_07614_),
    .Y(_07615_));
 sky130_fd_sc_hd__xor2_1 _14445_ (.A(_07603_),
    .B(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__nor2_1 _14446_ (.A(_07603_),
    .B(_07615_),
    .Y(_07617_));
 sky130_fd_sc_hd__a21o_1 _14447_ (.A1(_07601_),
    .A2(_07616_),
    .B1(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__xnor2_1 _14448_ (.A(_07599_),
    .B(_07618_),
    .Y(_07619_));
 sky130_fd_sc_hd__or2b_1 _14449_ (.A(_07599_),
    .B_N(_07618_),
    .X(_07620_));
 sky130_fd_sc_hd__a21boi_1 _14450_ (.A1(_07598_),
    .A2(_07619_),
    .B1_N(_07620_),
    .Y(_07621_));
 sky130_fd_sc_hd__or2_1 _14451_ (.A(_07572_),
    .B(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__and2_1 _14452_ (.A(_07519_),
    .B(_07565_),
    .X(_07623_));
 sky130_fd_sc_hd__or2_1 _14453_ (.A(_07566_),
    .B(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__nor2_1 _14454_ (.A(_07622_),
    .B(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__xnor2_1 _14455_ (.A(_07571_),
    .B(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__inv_2 _14456_ (.A(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__nand2_1 _14457_ (.A(_07572_),
    .B(_07621_),
    .Y(_07628_));
 sky130_fd_sc_hd__and2_1 _14458_ (.A(_07622_),
    .B(_07628_),
    .X(_07629_));
 sky130_fd_sc_hd__or2_1 _14459_ (.A(_06814_),
    .B(_07396_),
    .X(_07630_));
 sky130_fd_sc_hd__or3b_1 _14460_ (.A(_07630_),
    .B(_07440_),
    .C_N(_07372_),
    .X(_07631_));
 sky130_fd_sc_hd__nor2_1 _14461_ (.A(_07440_),
    .B(_07397_),
    .Y(_07632_));
 sky130_fd_sc_hd__a21o_1 _14462_ (.A1(_06826_),
    .A2(_07372_),
    .B1(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__nor2_1 _14463_ (.A(_07223_),
    .B(_07405_),
    .Y(_07634_));
 sky130_fd_sc_hd__nand3_1 _14464_ (.A(_07631_),
    .B(_07633_),
    .C(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__xnor2_1 _14465_ (.A(_07588_),
    .B(_07591_),
    .Y(_07636_));
 sky130_fd_sc_hd__a21o_1 _14466_ (.A1(_07631_),
    .A2(_07635_),
    .B1(_07636_),
    .X(_07637_));
 sky130_fd_sc_hd__nand3_1 _14467_ (.A(_07631_),
    .B(_07635_),
    .C(_07636_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_1 _14468_ (.A(_07637_),
    .B(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__or2_1 _14469_ (.A(_07281_),
    .B(_07471_),
    .X(_07640_));
 sky130_fd_sc_hd__inv_2 _14470_ (.A(_07640_),
    .Y(_07641_));
 sky130_fd_sc_hd__or2_1 _14471_ (.A(_07423_),
    .B(_07522_),
    .X(_07642_));
 sky130_fd_sc_hd__o22a_1 _14472_ (.A1(_07281_),
    .A2(_07408_),
    .B1(_07471_),
    .B2(_07387_),
    .X(_07643_));
 sky130_fd_sc_hd__a21o_1 _14473_ (.A1(_07590_),
    .A2(_07641_),
    .B1(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__o2bb2a_1 _14474_ (.A1_N(_07590_),
    .A2_N(_07641_),
    .B1(_07642_),
    .B2(_07644_),
    .X(_07645_));
 sky130_fd_sc_hd__or2_1 _14475_ (.A(_07639_),
    .B(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__xnor2_1 _14476_ (.A(_07575_),
    .B(_07577_),
    .Y(_07647_));
 sky130_fd_sc_hd__a21oi_2 _14477_ (.A1(_07637_),
    .A2(_07646_),
    .B1(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__xnor2_1 _14478_ (.A(_07601_),
    .B(_07616_),
    .Y(_07649_));
 sky130_fd_sc_hd__and3_1 _14479_ (.A(_07637_),
    .B(_07646_),
    .C(_07647_),
    .X(_07650_));
 sky130_fd_sc_hd__nor2_1 _14480_ (.A(_07648_),
    .B(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__xnor2_2 _14481_ (.A(_07604_),
    .B(_07613_),
    .Y(_07652_));
 sky130_fd_sc_hd__xor2_1 _14482_ (.A(_07639_),
    .B(_07645_),
    .X(_07653_));
 sky130_fd_sc_hd__xnor2_1 _14483_ (.A(_07606_),
    .B(_07611_),
    .Y(_07654_));
 sky130_fd_sc_hd__a21o_1 _14484_ (.A1(_07631_),
    .A2(_07633_),
    .B1(_07634_),
    .X(_07655_));
 sky130_fd_sc_hd__and2_1 _14485_ (.A(_07635_),
    .B(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__o21a_1 _14486_ (.A1(_06864_),
    .A2(_06870_),
    .B1(_07370_),
    .X(_07657_));
 sky130_fd_sc_hd__nand2_1 _14487_ (.A(_07609_),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__nand4_2 _14488_ (.A(_06864_),
    .B(_06870_),
    .C(_07373_),
    .D(_07370_),
    .Y(_07659_));
 sky130_fd_sc_hd__nand2_1 _14489_ (.A(_07608_),
    .B(_07659_),
    .Y(_07660_));
 sky130_fd_sc_hd__xnor2_1 _14490_ (.A(_07658_),
    .B(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__or2b_1 _14491_ (.A(_07658_),
    .B_N(_07660_),
    .X(_07662_));
 sky130_fd_sc_hd__a21bo_1 _14492_ (.A1(_07656_),
    .A2(_07661_),
    .B1_N(_07662_),
    .X(_07663_));
 sky130_fd_sc_hd__xnor2_1 _14493_ (.A(_07654_),
    .B(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__and2b_1 _14494_ (.A_N(_07654_),
    .B(_07663_),
    .X(_07665_));
 sky130_fd_sc_hd__a21oi_2 _14495_ (.A1(_07653_),
    .A2(_07664_),
    .B1(_07665_),
    .Y(_07666_));
 sky130_fd_sc_hd__xor2_2 _14496_ (.A(_07652_),
    .B(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__nor2_1 _14497_ (.A(_07652_),
    .B(_07666_),
    .Y(_07668_));
 sky130_fd_sc_hd__a21oi_1 _14498_ (.A1(_07651_),
    .A2(_07667_),
    .B1(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__xor2_1 _14499_ (.A(_07649_),
    .B(_07669_),
    .X(_07670_));
 sky130_fd_sc_hd__xnor2_1 _14500_ (.A(_07648_),
    .B(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__nor2_1 _14501_ (.A(_06814_),
    .B(_07405_),
    .Y(_07672_));
 sky130_fd_sc_hd__nand2_1 _14502_ (.A(_07632_),
    .B(_07672_),
    .Y(_07673_));
 sky130_fd_sc_hd__nor2_1 _14503_ (.A(_07440_),
    .B(_07404_),
    .Y(_07674_));
 sky130_fd_sc_hd__xnor2_1 _14504_ (.A(_07630_),
    .B(_07674_),
    .Y(_07675_));
 sky130_fd_sc_hd__nor2_1 _14505_ (.A(_07223_),
    .B(_07409_),
    .Y(_07676_));
 sky130_fd_sc_hd__nand2_1 _14506_ (.A(_07675_),
    .B(_07676_),
    .Y(_07677_));
 sky130_fd_sc_hd__xnor2_1 _14507_ (.A(_07642_),
    .B(_07644_),
    .Y(_07678_));
 sky130_fd_sc_hd__a21o_1 _14508_ (.A1(_07673_),
    .A2(_07677_),
    .B1(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__nand3_1 _14509_ (.A(_07673_),
    .B(_07677_),
    .C(_07678_),
    .Y(_07680_));
 sky130_fd_sc_hd__nand2_1 _14510_ (.A(_07679_),
    .B(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__nor2_1 _14511_ (.A(_07387_),
    .B(_07472_),
    .Y(_07682_));
 sky130_fd_sc_hd__nor2_1 _14512_ (.A(_07281_),
    .B(_07522_),
    .Y(_07683_));
 sky130_fd_sc_hd__o21a_1 _14513_ (.A1(_07387_),
    .A2(_07522_),
    .B1(_07640_),
    .X(_07684_));
 sky130_fd_sc_hd__a21oi_1 _14514_ (.A1(_07682_),
    .A2(_07683_),
    .B1(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__or3b_1 _14515_ (.A(_07423_),
    .B(_07573_),
    .C_N(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__o31a_1 _14516_ (.A1(_07387_),
    .A2(_07523_),
    .A3(_07640_),
    .B1(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__or2_1 _14517_ (.A(_07681_),
    .B(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__o22a_1 _14518_ (.A1(_07330_),
    .A2(_07573_),
    .B1(_07523_),
    .B2(_07143_),
    .X(_07689_));
 sky130_fd_sc_hd__or2_1 _14519_ (.A(_07575_),
    .B(_07689_),
    .X(_07690_));
 sky130_fd_sc_hd__a21oi_4 _14520_ (.A1(_07679_),
    .A2(_07688_),
    .B1(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__xnor2_2 _14521_ (.A(_07651_),
    .B(_07667_),
    .Y(_07692_));
 sky130_fd_sc_hd__and3_1 _14522_ (.A(_07679_),
    .B(_07688_),
    .C(_07690_),
    .X(_07693_));
 sky130_fd_sc_hd__nor2_1 _14523_ (.A(_07691_),
    .B(_07693_),
    .Y(_07694_));
 sky130_fd_sc_hd__xor2_1 _14524_ (.A(_07653_),
    .B(_07664_),
    .X(_07695_));
 sky130_fd_sc_hd__xor2_1 _14525_ (.A(_07681_),
    .B(_07687_),
    .X(_07696_));
 sky130_fd_sc_hd__xnor2_1 _14526_ (.A(_07656_),
    .B(_07661_),
    .Y(_07697_));
 sky130_fd_sc_hd__a22o_1 _14527_ (.A1(_06870_),
    .A2(_07373_),
    .B1(_07370_),
    .B2(_06864_),
    .X(_07698_));
 sky130_fd_sc_hd__nor2_1 _14528_ (.A(_07227_),
    .B(_07397_),
    .Y(_07699_));
 sky130_fd_sc_hd__a22o_1 _14529_ (.A1(_06872_),
    .A2(_07372_),
    .B1(_07369_),
    .B2(_06871_),
    .X(_07700_));
 sky130_fd_sc_hd__nand3_1 _14530_ (.A(_06810_),
    .B(_07373_),
    .C(_07370_),
    .Y(_07701_));
 sky130_fd_sc_hd__a21bo_2 _14531_ (.A1(_07699_),
    .A2(_07700_),
    .B1_N(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__or2_1 _14532_ (.A(_07675_),
    .B(_07676_),
    .X(_07703_));
 sky130_fd_sc_hd__and2_1 _14533_ (.A(_07677_),
    .B(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__nand2_1 _14534_ (.A(_07659_),
    .B(_07698_),
    .Y(_07705_));
 sky130_fd_sc_hd__xnor2_2 _14535_ (.A(_07705_),
    .B(_07702_),
    .Y(_07706_));
 sky130_fd_sc_hd__a32oi_4 _14536_ (.A1(_07659_),
    .A2(_07698_),
    .A3(_07702_),
    .B1(_07704_),
    .B2(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__xor2_1 _14537_ (.A(_07697_),
    .B(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__nor2_1 _14538_ (.A(_07697_),
    .B(_07707_),
    .Y(_07709_));
 sky130_fd_sc_hd__a21oi_1 _14539_ (.A1(_07696_),
    .A2(_07708_),
    .B1(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__xnor2_1 _14540_ (.A(_07695_),
    .B(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__or2b_1 _14541_ (.A(_07710_),
    .B_N(_07695_),
    .X(_07712_));
 sky130_fd_sc_hd__a21boi_2 _14542_ (.A1(_07694_),
    .A2(_07711_),
    .B1_N(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__xor2_2 _14543_ (.A(_07692_),
    .B(_07713_),
    .X(_07714_));
 sky130_fd_sc_hd__nor2_1 _14544_ (.A(_07692_),
    .B(_07713_),
    .Y(_07715_));
 sky130_fd_sc_hd__a21oi_2 _14545_ (.A1(_07691_),
    .A2(_07714_),
    .B1(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__nor2_1 _14546_ (.A(_07671_),
    .B(_07716_),
    .Y(_07717_));
 sky130_fd_sc_hd__xnor2_1 _14547_ (.A(_07598_),
    .B(_07619_),
    .Y(_07718_));
 sky130_fd_sc_hd__nor2_1 _14548_ (.A(_07649_),
    .B(_07669_),
    .Y(_07719_));
 sky130_fd_sc_hd__a21oi_1 _14549_ (.A1(_07648_),
    .A2(_07670_),
    .B1(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__nor2_1 _14550_ (.A(_07718_),
    .B(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__and2_1 _14551_ (.A(_07718_),
    .B(_07720_),
    .X(_07722_));
 sky130_fd_sc_hd__nor2_1 _14552_ (.A(_07721_),
    .B(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__and2_1 _14553_ (.A(_07717_),
    .B(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__nor2_1 _14554_ (.A(_07721_),
    .B(_07724_),
    .Y(_07725_));
 sky130_fd_sc_hd__xnor2_1 _14555_ (.A(_07629_),
    .B(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__xnor2_2 _14556_ (.A(_07691_),
    .B(_07714_),
    .Y(_07727_));
 sky130_fd_sc_hd__nor2_1 _14557_ (.A(_06814_),
    .B(_07409_),
    .Y(_07728_));
 sky130_fd_sc_hd__nand2_1 _14558_ (.A(_07674_),
    .B(_07728_),
    .Y(_07729_));
 sky130_fd_sc_hd__nor2_1 _14559_ (.A(_07440_),
    .B(_07409_),
    .Y(_07730_));
 sky130_fd_sc_hd__xnor2_1 _14560_ (.A(_07672_),
    .B(_07730_),
    .Y(_07731_));
 sky130_fd_sc_hd__or3_1 _14561_ (.A(_07223_),
    .B(_07472_),
    .C(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__o21bai_1 _14562_ (.A1(_07423_),
    .A2(_07573_),
    .B1_N(_07685_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand2_1 _14563_ (.A(_07686_),
    .B(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__nand3_1 _14564_ (.A(_07729_),
    .B(_07732_),
    .C(_07734_),
    .Y(_07735_));
 sky130_fd_sc_hd__nor2_1 _14565_ (.A(_07387_),
    .B(_07573_),
    .Y(_07736_));
 sky130_fd_sc_hd__and2_1 _14566_ (.A(_07683_),
    .B(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__a21o_1 _14567_ (.A1(_07729_),
    .A2(_07732_),
    .B1(_07734_),
    .X(_07738_));
 sky130_fd_sc_hd__a21boi_1 _14568_ (.A1(_07735_),
    .A2(_07737_),
    .B1_N(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__nor2_1 _14569_ (.A(_07574_),
    .B(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__xnor2_1 _14570_ (.A(_07694_),
    .B(_07711_),
    .Y(_07741_));
 sky130_fd_sc_hd__and2_1 _14571_ (.A(_07574_),
    .B(_07739_),
    .X(_07742_));
 sky130_fd_sc_hd__nor2_1 _14572_ (.A(_07740_),
    .B(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__xnor2_1 _14573_ (.A(_07696_),
    .B(_07708_),
    .Y(_07744_));
 sky130_fd_sc_hd__nand2_1 _14574_ (.A(_07738_),
    .B(_07735_),
    .Y(_07745_));
 sky130_fd_sc_hd__xnor2_1 _14575_ (.A(_07745_),
    .B(_07737_),
    .Y(_07746_));
 sky130_fd_sc_hd__xnor2_1 _14576_ (.A(_07704_),
    .B(_07706_),
    .Y(_07747_));
 sky130_fd_sc_hd__nor2_1 _14577_ (.A(_07223_),
    .B(_07472_),
    .Y(_07748_));
 sky130_fd_sc_hd__xnor2_1 _14578_ (.A(_07731_),
    .B(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__nand3_1 _14579_ (.A(_07701_),
    .B(_07699_),
    .C(_07700_),
    .Y(_07750_));
 sky130_fd_sc_hd__a21o_1 _14580_ (.A1(_07701_),
    .A2(_07700_),
    .B1(_07699_),
    .X(_07751_));
 sky130_fd_sc_hd__nor2_1 _14581_ (.A(_07227_),
    .B(_07405_),
    .Y(_07752_));
 sky130_fd_sc_hd__nor2_1 _14582_ (.A(_07230_),
    .B(_07397_),
    .Y(_07753_));
 sky130_fd_sc_hd__a21o_1 _14583_ (.A1(_06871_),
    .A2(_07373_),
    .B1(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__or2_1 _14584_ (.A(_06976_),
    .B(_07396_),
    .X(_07755_));
 sky130_fd_sc_hd__or3b_1 _14585_ (.A(_07755_),
    .B(_07230_),
    .C_N(_07372_),
    .X(_07756_));
 sky130_fd_sc_hd__a21bo_1 _14586_ (.A1(_07752_),
    .A2(_07754_),
    .B1_N(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__a21o_1 _14587_ (.A1(_07750_),
    .A2(_07751_),
    .B1(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__nand3_1 _14588_ (.A(_07750_),
    .B(_07751_),
    .C(_07757_),
    .Y(_07759_));
 sky130_fd_sc_hd__a21bo_1 _14589_ (.A1(_07749_),
    .A2(_07758_),
    .B1_N(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__xnor2_1 _14590_ (.A(_07747_),
    .B(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__or2b_1 _14591_ (.A(_07747_),
    .B_N(_07760_),
    .X(_07762_));
 sky130_fd_sc_hd__a21bo_1 _14592_ (.A1(_07746_),
    .A2(_07761_),
    .B1_N(_07762_),
    .X(_07763_));
 sky130_fd_sc_hd__xnor2_1 _14593_ (.A(_07744_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__or2b_1 _14594_ (.A(_07744_),
    .B_N(_07763_),
    .X(_07765_));
 sky130_fd_sc_hd__a21boi_1 _14595_ (.A1(_07743_),
    .A2(_07764_),
    .B1_N(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__xor2_1 _14596_ (.A(_07741_),
    .B(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__nor2_1 _14597_ (.A(_07741_),
    .B(_07766_),
    .Y(_07768_));
 sky130_fd_sc_hd__a21oi_2 _14598_ (.A1(_07740_),
    .A2(_07767_),
    .B1(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__nor2_1 _14599_ (.A(_07727_),
    .B(_07769_),
    .Y(_07770_));
 sky130_fd_sc_hd__xor2_1 _14600_ (.A(_07671_),
    .B(_07716_),
    .X(_07771_));
 sky130_fd_sc_hd__and2_1 _14601_ (.A(_07770_),
    .B(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__nor2_1 _14602_ (.A(_07717_),
    .B(_07772_),
    .Y(_07773_));
 sky130_fd_sc_hd__xnor2_1 _14603_ (.A(_07723_),
    .B(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__xor2_1 _14604_ (.A(_07727_),
    .B(_07769_),
    .X(_07775_));
 sky130_fd_sc_hd__nor2_1 _14605_ (.A(_07440_),
    .B(_07472_),
    .Y(_07776_));
 sky130_fd_sc_hd__nand2_1 _14606_ (.A(_07728_),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__or2_1 _14607_ (.A(_07728_),
    .B(_07776_),
    .X(_07778_));
 sky130_fd_sc_hd__nand2_1 _14608_ (.A(_07777_),
    .B(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__or3_1 _14609_ (.A(_07223_),
    .B(_07523_),
    .C(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__nor2_1 _14610_ (.A(_07683_),
    .B(_07736_),
    .Y(_07781_));
 sky130_fd_sc_hd__or2_1 _14611_ (.A(_07737_),
    .B(_07781_),
    .X(_07782_));
 sky130_fd_sc_hd__a21oi_2 _14612_ (.A1(_07777_),
    .A2(_07780_),
    .B1(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__xnor2_1 _14613_ (.A(_07746_),
    .B(_07761_),
    .Y(_07784_));
 sky130_fd_sc_hd__and3_1 _14614_ (.A(_07759_),
    .B(_07749_),
    .C(_07758_),
    .X(_07785_));
 sky130_fd_sc_hd__a21oi_1 _14615_ (.A1(_07759_),
    .A2(_07758_),
    .B1(_07749_),
    .Y(_07786_));
 sky130_fd_sc_hd__nor2_1 _14616_ (.A(_07223_),
    .B(_07523_),
    .Y(_07787_));
 sky130_fd_sc_hd__xnor2_1 _14617_ (.A(_07779_),
    .B(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__nand3_1 _14618_ (.A(_07756_),
    .B(_07752_),
    .C(_07754_),
    .Y(_07789_));
 sky130_fd_sc_hd__a21o_1 _14619_ (.A1(_07756_),
    .A2(_07754_),
    .B1(_07752_),
    .X(_07790_));
 sky130_fd_sc_hd__nor2_1 _14620_ (.A(_06976_),
    .B(_07405_),
    .Y(_07791_));
 sky130_fd_sc_hd__nor2_1 _14621_ (.A(_07227_),
    .B(_07409_),
    .Y(_07792_));
 sky130_fd_sc_hd__nor2_1 _14622_ (.A(_07230_),
    .B(_07405_),
    .Y(_07793_));
 sky130_fd_sc_hd__xnor2_1 _14623_ (.A(_07755_),
    .B(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__a22o_1 _14624_ (.A1(_07753_),
    .A2(_07791_),
    .B1(_07792_),
    .B2(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__a21o_1 _14625_ (.A1(_07789_),
    .A2(_07790_),
    .B1(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__and3_1 _14626_ (.A(_07789_),
    .B(_07790_),
    .C(_07795_),
    .X(_07797_));
 sky130_fd_sc_hd__a21oi_1 _14627_ (.A1(_07788_),
    .A2(_07796_),
    .B1(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__or3_1 _14628_ (.A(_07785_),
    .B(_07786_),
    .C(_07798_),
    .X(_07799_));
 sky130_fd_sc_hd__and3_1 _14629_ (.A(_07777_),
    .B(_07780_),
    .C(_07782_),
    .X(_07800_));
 sky130_fd_sc_hd__nor2_1 _14630_ (.A(_07783_),
    .B(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__o21ai_1 _14631_ (.A1(_07785_),
    .A2(_07786_),
    .B1(_07798_),
    .Y(_07802_));
 sky130_fd_sc_hd__nand3_1 _14632_ (.A(_07799_),
    .B(_07801_),
    .C(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__and2_1 _14633_ (.A(_07799_),
    .B(_07803_),
    .X(_07804_));
 sky130_fd_sc_hd__nand2_1 _14634_ (.A(_07784_),
    .B(_07804_),
    .Y(_07805_));
 sky130_fd_sc_hd__nor2_1 _14635_ (.A(_07784_),
    .B(_07804_),
    .Y(_07806_));
 sky130_fd_sc_hd__a21oi_2 _14636_ (.A1(_07783_),
    .A2(_07805_),
    .B1(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__xnor2_2 _14637_ (.A(_07743_),
    .B(_07764_),
    .Y(_07808_));
 sky130_fd_sc_hd__xor2_1 _14638_ (.A(_07740_),
    .B(_07767_),
    .X(_07809_));
 sky130_fd_sc_hd__nor3b_4 _14639_ (.A(_07807_),
    .B(_07808_),
    .C_N(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__and2_1 _14640_ (.A(_07775_),
    .B(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__xor2_1 _14641_ (.A(_07775_),
    .B(_07810_),
    .X(_07812_));
 sky130_fd_sc_hd__and2b_1 _14642_ (.A_N(_07806_),
    .B(_07805_),
    .X(_07813_));
 sky130_fd_sc_hd__xor2_1 _14643_ (.A(_07783_),
    .B(_07813_),
    .X(_07814_));
 sky130_fd_sc_hd__or2_1 _14644_ (.A(_07281_),
    .B(_07573_),
    .X(_07815_));
 sky130_fd_sc_hd__nor2_1 _14645_ (.A(_06814_),
    .B(_07523_),
    .Y(_07816_));
 sky130_fd_sc_hd__o22a_1 _14646_ (.A1(_06814_),
    .A2(_07472_),
    .B1(_07523_),
    .B2(_07440_),
    .X(_07817_));
 sky130_fd_sc_hd__a21o_1 _14647_ (.A1(_07776_),
    .A2(_07816_),
    .B1(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__inv_2 _14648_ (.A(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__nor2_1 _14649_ (.A(_07223_),
    .B(_07573_),
    .Y(_07820_));
 sky130_fd_sc_hd__a22oi_1 _14650_ (.A1(_07776_),
    .A2(_07816_),
    .B1(_07819_),
    .B2(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__nor2_1 _14651_ (.A(_07815_),
    .B(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__a21o_1 _14652_ (.A1(_07799_),
    .A2(_07802_),
    .B1(_07801_),
    .X(_07823_));
 sky130_fd_sc_hd__xnor2_1 _14653_ (.A(_07792_),
    .B(_07794_),
    .Y(_07824_));
 sky130_fd_sc_hd__nor2_1 _14654_ (.A(_06976_),
    .B(_07409_),
    .Y(_07825_));
 sky130_fd_sc_hd__or2_1 _14655_ (.A(_07227_),
    .B(_07472_),
    .X(_07826_));
 sky130_fd_sc_hd__o22a_1 _14656_ (.A1(_06976_),
    .A2(_07405_),
    .B1(_07409_),
    .B2(_07230_),
    .X(_07827_));
 sky130_fd_sc_hd__a21o_1 _14657_ (.A1(_07793_),
    .A2(_07825_),
    .B1(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__o2bb2a_1 _14658_ (.A1_N(_07793_),
    .A2_N(_07825_),
    .B1(_07826_),
    .B2(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__or2_1 _14659_ (.A(_07824_),
    .B(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__xnor2_1 _14660_ (.A(_07818_),
    .B(_07820_),
    .Y(_07831_));
 sky130_fd_sc_hd__nand2_1 _14661_ (.A(_07824_),
    .B(_07829_),
    .Y(_07832_));
 sky130_fd_sc_hd__and2_1 _14662_ (.A(_07830_),
    .B(_07832_),
    .X(_07833_));
 sky130_fd_sc_hd__nand2_1 _14663_ (.A(_07831_),
    .B(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__and2b_1 _14664_ (.A_N(_07797_),
    .B(_07796_),
    .X(_07835_));
 sky130_fd_sc_hd__xnor2_1 _14665_ (.A(_07788_),
    .B(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__a21o_1 _14666_ (.A1(_07830_),
    .A2(_07834_),
    .B1(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__inv_2 _14667_ (.A(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__and2_1 _14668_ (.A(_07815_),
    .B(_07821_),
    .X(_07839_));
 sky130_fd_sc_hd__nor2_1 _14669_ (.A(_07822_),
    .B(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__nand3_1 _14670_ (.A(_07836_),
    .B(_07830_),
    .C(_07834_),
    .Y(_07841_));
 sky130_fd_sc_hd__and3_1 _14671_ (.A(_07837_),
    .B(_07840_),
    .C(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__a211o_1 _14672_ (.A1(_07803_),
    .A2(_07823_),
    .B1(_07838_),
    .C1(_07842_),
    .X(_07843_));
 sky130_fd_sc_hd__o211ai_1 _14673_ (.A1(_07838_),
    .A2(_07842_),
    .B1(_07803_),
    .C1(_07823_),
    .Y(_07844_));
 sky130_fd_sc_hd__a21bo_1 _14674_ (.A1(_07822_),
    .A2(_07843_),
    .B1_N(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__xor2_1 _14675_ (.A(_07808_),
    .B(_07807_),
    .X(_07846_));
 sky130_fd_sc_hd__and4_2 _14676_ (.A(_07809_),
    .B(_07814_),
    .C(_07845_),
    .D(_07846_),
    .X(_07847_));
 sky130_fd_sc_hd__xor2_1 _14677_ (.A(_07812_),
    .B(_07847_),
    .X(_07848_));
 sky130_fd_sc_hd__nor2_1 _14678_ (.A(_07814_),
    .B(_07845_),
    .Y(_07849_));
 sky130_fd_sc_hd__and3_1 _14679_ (.A(_07822_),
    .B(_07844_),
    .C(_07843_),
    .X(_07850_));
 sky130_fd_sc_hd__a21oi_1 _14680_ (.A1(_07844_),
    .A2(_07843_),
    .B1(_07822_),
    .Y(_07851_));
 sky130_fd_sc_hd__nor2_1 _14681_ (.A(_07440_),
    .B(_07573_),
    .Y(_07852_));
 sky130_fd_sc_hd__and2_1 _14682_ (.A(_07816_),
    .B(_07852_),
    .X(_07853_));
 sky130_fd_sc_hd__or2_1 _14683_ (.A(_07227_),
    .B(_07523_),
    .X(_07854_));
 sky130_fd_sc_hd__nor2_1 _14684_ (.A(_07230_),
    .B(_07472_),
    .Y(_07855_));
 sky130_fd_sc_hd__xnor2_1 _14685_ (.A(_07825_),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__or2_1 _14686_ (.A(_07854_),
    .B(_07856_),
    .X(_07857_));
 sky130_fd_sc_hd__nand2_1 _14687_ (.A(_07854_),
    .B(_07856_),
    .Y(_07858_));
 sky130_fd_sc_hd__nand2_1 _14688_ (.A(_07857_),
    .B(_07858_),
    .Y(_07859_));
 sky130_fd_sc_hd__or2_1 _14689_ (.A(_06976_),
    .B(_07472_),
    .X(_07860_));
 sky130_fd_sc_hd__nor2_1 _14690_ (.A(_07227_),
    .B(_07573_),
    .Y(_07861_));
 sky130_fd_sc_hd__nor2_1 _14691_ (.A(_07230_),
    .B(_07523_),
    .Y(_07862_));
 sky130_fd_sc_hd__xnor2_1 _14692_ (.A(_07860_),
    .B(_07862_),
    .Y(_07863_));
 sky130_fd_sc_hd__nand2_1 _14693_ (.A(_07861_),
    .B(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__o31a_1 _14694_ (.A1(_07230_),
    .A2(_07523_),
    .A3(_07860_),
    .B1(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__or2_1 _14695_ (.A(_07859_),
    .B(_07865_),
    .X(_07866_));
 sky130_fd_sc_hd__or2_1 _14696_ (.A(_06814_),
    .B(_07573_),
    .X(_07867_));
 sky130_fd_sc_hd__nand2_1 _14697_ (.A(_07859_),
    .B(_07865_),
    .Y(_07868_));
 sky130_fd_sc_hd__nand2_1 _14698_ (.A(_07866_),
    .B(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__or2_1 _14699_ (.A(_07867_),
    .B(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__and3_1 _14700_ (.A(_06810_),
    .B(_07315_),
    .C(_07864_),
    .X(_07871_));
 sky130_fd_sc_hd__o21ai_1 _14701_ (.A1(_07861_),
    .A2(_07863_),
    .B1(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__a21o_1 _14702_ (.A1(_07867_),
    .A2(_07869_),
    .B1(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__xor2_1 _14703_ (.A(_07816_),
    .B(_07852_),
    .X(_07874_));
 sky130_fd_sc_hd__xnor2_1 _14704_ (.A(_07826_),
    .B(_07828_),
    .Y(_07875_));
 sky130_fd_sc_hd__a21bo_1 _14705_ (.A1(_07825_),
    .A2(_07855_),
    .B1_N(_07857_),
    .X(_07876_));
 sky130_fd_sc_hd__xnor2_1 _14706_ (.A(_07875_),
    .B(_07876_),
    .Y(_07877_));
 sky130_fd_sc_hd__nand2_1 _14707_ (.A(_07874_),
    .B(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__or2_1 _14708_ (.A(_07874_),
    .B(_07877_),
    .X(_07879_));
 sky130_fd_sc_hd__o2bb2a_1 _14709_ (.A1_N(_07878_),
    .A2_N(_07879_),
    .B1(_07866_),
    .B2(_07873_),
    .X(_07880_));
 sky130_fd_sc_hd__a31oi_1 _14710_ (.A1(_07866_),
    .A2(_07870_),
    .A3(_07873_),
    .B1(_07880_),
    .Y(_07881_));
 sky130_fd_sc_hd__or2b_1 _14711_ (.A(_07875_),
    .B_N(_07876_),
    .X(_07882_));
 sky130_fd_sc_hd__and2_1 _14712_ (.A(_07882_),
    .B(_07878_),
    .X(_07883_));
 sky130_fd_sc_hd__or2_1 _14713_ (.A(_07831_),
    .B(_07833_),
    .X(_07884_));
 sky130_fd_sc_hd__nand2_1 _14714_ (.A(_07834_),
    .B(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__a2bb2o_1 _14715_ (.A1_N(_07853_),
    .A2_N(_07881_),
    .B1(_07883_),
    .B2(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__a21o_1 _14716_ (.A1(_07882_),
    .A2(_07878_),
    .B1(_07885_),
    .X(_07887_));
 sky130_fd_sc_hd__nand2_1 _14717_ (.A(_07853_),
    .B(_07881_),
    .Y(_07888_));
 sky130_fd_sc_hd__a21oi_1 _14718_ (.A1(_07837_),
    .A2(_07841_),
    .B1(_07840_),
    .Y(_07889_));
 sky130_fd_sc_hd__a311o_1 _14719_ (.A1(_07886_),
    .A2(_07887_),
    .A3(_07888_),
    .B1(_07889_),
    .C1(_07842_),
    .X(_07890_));
 sky130_fd_sc_hd__or3_1 _14720_ (.A(_07850_),
    .B(_07851_),
    .C(_07890_),
    .X(_07891_));
 sky130_fd_sc_hd__and4bb_2 _14721_ (.A_N(_07849_),
    .B_N(_07891_),
    .C(_07809_),
    .D(_07846_),
    .X(_07892_));
 sky130_fd_sc_hd__and2_1 _14722_ (.A(_07812_),
    .B(_07847_),
    .X(_07893_));
 sky130_fd_sc_hd__a21o_1 _14723_ (.A1(_07848_),
    .A2(_07892_),
    .B1(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__nor2_1 _14724_ (.A(_07770_),
    .B(_07811_),
    .Y(_07895_));
 sky130_fd_sc_hd__xnor2_1 _14725_ (.A(_07771_),
    .B(_07895_),
    .Y(_07896_));
 sky130_fd_sc_hd__a22o_1 _14726_ (.A1(_07811_),
    .A2(_07771_),
    .B1(_07894_),
    .B2(_07896_),
    .X(_07897_));
 sky130_fd_sc_hd__a22o_1 _14727_ (.A1(_07772_),
    .A2(_07723_),
    .B1(_07774_),
    .B2(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__a22o_1 _14728_ (.A1(_07629_),
    .A2(_07724_),
    .B1(_07726_),
    .B2(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__nand2_1 _14729_ (.A(_07721_),
    .B(_07629_),
    .Y(_07900_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(_07622_),
    .B(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__xnor2_1 _14731_ (.A(_07624_),
    .B(_07901_),
    .Y(_07902_));
 sky130_fd_sc_hd__o2bb2a_1 _14732_ (.A1_N(_07899_),
    .A2_N(_07902_),
    .B1(_07624_),
    .B2(_07900_),
    .X(_07903_));
 sky130_fd_sc_hd__nor2_1 _14733_ (.A(_07508_),
    .B(_07510_),
    .Y(_07904_));
 sky130_fd_sc_hd__nor2_1 _14734_ (.A(_07511_),
    .B(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__xnor2_1 _14735_ (.A(_07569_),
    .B(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__and2b_1 _14736_ (.A_N(_07571_),
    .B(_07625_),
    .X(_07907_));
 sky130_fd_sc_hd__o21ai_1 _14737_ (.A1(_07569_),
    .A2(_07907_),
    .B1(_07905_),
    .Y(_07908_));
 sky130_fd_sc_hd__o31a_1 _14738_ (.A1(_07627_),
    .A2(_07903_),
    .A3(_07906_),
    .B1(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__o21ai_2 _14739_ (.A1(_07517_),
    .A2(_07909_),
    .B1(_07514_),
    .Y(_07910_));
 sky130_fd_sc_hd__xor2_4 _14740_ (.A(_07467_),
    .B(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__nand2_1 _14741_ (.A(_07462_),
    .B(_07514_),
    .Y(_07912_));
 sky130_fd_sc_hd__nand2_1 _14742_ (.A(_07516_),
    .B(_07467_),
    .Y(_07913_));
 sky130_fd_sc_hd__o2bb2a_1 _14743_ (.A1_N(_07466_),
    .A2_N(_07912_),
    .B1(_07908_),
    .B2(_07913_),
    .X(_07914_));
 sky130_fd_sc_hd__or4_1 _14744_ (.A(_07627_),
    .B(_07903_),
    .C(_07906_),
    .D(_07913_),
    .X(_07915_));
 sky130_fd_sc_hd__o21bai_1 _14745_ (.A1(_07330_),
    .A2(_07388_),
    .B1_N(_07375_),
    .Y(_07916_));
 sky130_fd_sc_hd__nor4_1 _14746_ (.A(_06567_),
    .B(_07384_),
    .C(_07465_),
    .D(_07916_),
    .Y(_07917_));
 sky130_fd_sc_hd__a21o_1 _14747_ (.A1(_07914_),
    .A2(_07915_),
    .B1(_07917_),
    .X(_07918_));
 sky130_fd_sc_hd__nand3_1 _14748_ (.A(_07914_),
    .B(_07915_),
    .C(_07917_),
    .Y(_07919_));
 sky130_fd_sc_hd__and3_2 _14749_ (.A(_06845_),
    .B(_07918_),
    .C(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__a211o_1 _14750_ (.A1(_06626_),
    .A2(_07911_),
    .B1(_07920_),
    .C1(_06792_),
    .X(_07921_));
 sky130_fd_sc_hd__xnor2_1 _14751_ (.A(_07516_),
    .B(_07909_),
    .Y(_07922_));
 sky130_fd_sc_hd__o21bai_1 _14752_ (.A1(_07627_),
    .A2(_07903_),
    .B1_N(_07907_),
    .Y(_07923_));
 sky130_fd_sc_hd__xnor2_1 _14753_ (.A(_07906_),
    .B(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__mux2_1 _14754_ (.A0(_07922_),
    .A1(_07924_),
    .S(_06626_),
    .X(_07925_));
 sky130_fd_sc_hd__or2_1 _14755_ (.A(_06642_),
    .B(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__o21ai_1 _14756_ (.A1(_06845_),
    .A2(_07918_),
    .B1(_06632_),
    .Y(_07927_));
 sky130_fd_sc_hd__and3_1 _14757_ (.A(_06751_),
    .B(_06792_),
    .C(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__a31oi_1 _14758_ (.A1(_06606_),
    .A2(_07921_),
    .A3(_07926_),
    .B1(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__nand2_1 _14759_ (.A(_06602_),
    .B(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__buf_2 _14760_ (.A(_06845_),
    .X(_07931_));
 sky130_fd_sc_hd__xnor2_1 _14761_ (.A(_07626_),
    .B(_07903_),
    .Y(_07932_));
 sky130_fd_sc_hd__xnor2_1 _14762_ (.A(_07899_),
    .B(_07902_),
    .Y(_07933_));
 sky130_fd_sc_hd__nor2_1 _14763_ (.A(_07931_),
    .B(_07933_),
    .Y(_07934_));
 sky130_fd_sc_hd__a21oi_1 _14764_ (.A1(_07931_),
    .A2(_07932_),
    .B1(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__xnor2_1 _14765_ (.A(_07897_),
    .B(_07774_),
    .Y(_07936_));
 sky130_fd_sc_hd__or2_1 _14766_ (.A(_06845_),
    .B(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__xnor2_1 _14767_ (.A(_07898_),
    .B(_07726_),
    .Y(_07938_));
 sky130_fd_sc_hd__or2_1 _14768_ (.A(_06625_),
    .B(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__nand2_1 _14769_ (.A(_07937_),
    .B(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__nand2_1 _14770_ (.A(_06792_),
    .B(_07940_),
    .Y(_07941_));
 sky130_fd_sc_hd__o21ai_1 _14771_ (.A1(_06792_),
    .A2(_07935_),
    .B1(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__xnor2_1 _14772_ (.A(_07894_),
    .B(_07896_),
    .Y(_07943_));
 sky130_fd_sc_hd__or2_1 _14773_ (.A(_06625_),
    .B(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__xnor2_1 _14774_ (.A(_07848_),
    .B(_07892_),
    .Y(_07945_));
 sky130_fd_sc_hd__or2_1 _14775_ (.A(_07931_),
    .B(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__nand2_1 _14776_ (.A(_07944_),
    .B(_07946_),
    .Y(_07947_));
 sky130_fd_sc_hd__a221o_1 _14777_ (.A1(_06751_),
    .A2(_07942_),
    .B1(_07947_),
    .B2(_06729_),
    .C1(_06602_),
    .X(_07948_));
 sky130_fd_sc_hd__or2_2 _14778_ (.A(_06567_),
    .B(_06578_),
    .X(_07949_));
 sky130_fd_sc_hd__clkbuf_4 _14779_ (.A(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__a31o_1 _14780_ (.A1(_06545_),
    .A2(_07930_),
    .A3(_07948_),
    .B1(_07950_),
    .X(_07951_));
 sky130_fd_sc_hd__and4b_1 _14781_ (.A_N(_04493_),
    .B(_04495_),
    .C(_04490_),
    .D(_06335_),
    .X(_07952_));
 sky130_fd_sc_hd__clkbuf_4 _14782_ (.A(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__clkbuf_4 _14783_ (.A(_07953_),
    .X(_07954_));
 sky130_fd_sc_hd__mux2_1 _14784_ (.A0(\rbzero.wall_tracer.stepDistY[-11] ),
    .A1(_07951_),
    .S(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__clkbuf_1 _14785_ (.A(_07955_),
    .X(_00391_));
 sky130_fd_sc_hd__buf_2 _14786_ (.A(_06698_),
    .X(_07956_));
 sky130_fd_sc_hd__and3_1 _14787_ (.A(_06625_),
    .B(_07918_),
    .C(_07919_),
    .X(_07957_));
 sky130_fd_sc_hd__a211o_1 _14788_ (.A1(_07931_),
    .A2(_07911_),
    .B1(_07957_),
    .C1(_06739_),
    .X(_07958_));
 sky130_fd_sc_hd__clkbuf_4 _14789_ (.A(_06682_),
    .X(_07959_));
 sky130_fd_sc_hd__nor2_1 _14790_ (.A(_06626_),
    .B(_07918_),
    .Y(_07960_));
 sky130_fd_sc_hd__or2_1 _14791_ (.A(_07959_),
    .B(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__a21o_1 _14792_ (.A1(_06606_),
    .A2(_06672_),
    .B1(_06661_),
    .X(_07962_));
 sky130_fd_sc_hd__and2_1 _14793_ (.A(_06588_),
    .B(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__a31o_1 _14794_ (.A1(_07956_),
    .A2(_07958_),
    .A3(_07961_),
    .B1(_07963_),
    .X(_07964_));
 sky130_fd_sc_hd__nand2_2 _14795_ (.A(_06588_),
    .B(_07962_),
    .Y(_07965_));
 sky130_fd_sc_hd__nor2_1 _14796_ (.A(_06845_),
    .B(_07938_),
    .Y(_07966_));
 sky130_fd_sc_hd__nor2_1 _14797_ (.A(_06625_),
    .B(_07936_),
    .Y(_07967_));
 sky130_fd_sc_hd__or2_1 _14798_ (.A(_07966_),
    .B(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__nor2_1 _14799_ (.A(_06845_),
    .B(_07943_),
    .Y(_07969_));
 sky130_fd_sc_hd__o21bai_1 _14800_ (.A1(_06626_),
    .A2(_07945_),
    .B1_N(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__mux2_1 _14801_ (.A0(_07922_),
    .A1(_07924_),
    .S(_06845_),
    .X(_07971_));
 sky130_fd_sc_hd__nor2_1 _14802_ (.A(_06625_),
    .B(_07933_),
    .Y(_07972_));
 sky130_fd_sc_hd__and2_1 _14803_ (.A(_06625_),
    .B(_07932_),
    .X(_07973_));
 sky130_fd_sc_hd__or2_1 _14804_ (.A(_07972_),
    .B(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__mux4_2 _14805_ (.A0(_07968_),
    .A1(_07970_),
    .A2(_07971_),
    .A3(_07974_),
    .S0(_06682_),
    .S1(_06673_),
    .X(_07975_));
 sky130_fd_sc_hd__or2_1 _14806_ (.A(_07965_),
    .B(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__a31o_1 _14807_ (.A1(_06545_),
    .A2(_07964_),
    .A3(_07976_),
    .B1(_07950_),
    .X(_07977_));
 sky130_fd_sc_hd__mux2_1 _14808_ (.A0(\rbzero.wall_tracer.stepDistY[-10] ),
    .A1(_07977_),
    .S(_07954_),
    .X(_07978_));
 sky130_fd_sc_hd__clkbuf_1 _14809_ (.A(_07978_),
    .X(_00392_));
 sky130_fd_sc_hd__inv_2 _14810_ (.A(_06583_),
    .Y(_07979_));
 sky130_fd_sc_hd__or2_1 _14811_ (.A(_06792_),
    .B(_07927_),
    .X(_07980_));
 sky130_fd_sc_hd__a211o_1 _14812_ (.A1(_06626_),
    .A2(_07911_),
    .B1(_07920_),
    .C1(_06642_),
    .X(_07981_));
 sky130_fd_sc_hd__and3_1 _14813_ (.A(_06606_),
    .B(_07980_),
    .C(_07981_),
    .X(_07982_));
 sky130_fd_sc_hd__nor2_1 _14814_ (.A(_06642_),
    .B(_07935_),
    .Y(_07983_));
 sky130_fd_sc_hd__a211o_1 _14815_ (.A1(_06642_),
    .A2(_07925_),
    .B1(_07983_),
    .C1(_06606_),
    .X(_07984_));
 sky130_fd_sc_hd__nor2_1 _14816_ (.A(_06695_),
    .B(_06602_),
    .Y(_07985_));
 sky130_fd_sc_hd__o221a_1 _14817_ (.A1(_06692_),
    .A2(_07940_),
    .B1(_07947_),
    .B2(_06754_),
    .C1(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__a21o_1 _14818_ (.A1(_07984_),
    .A2(_07986_),
    .B1(_07950_),
    .X(_07987_));
 sky130_fd_sc_hd__a21o_1 _14819_ (.A1(_07979_),
    .A2(_07982_),
    .B1(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__mux2_1 _14820_ (.A0(\rbzero.wall_tracer.stepDistY[-9] ),
    .A1(_07988_),
    .S(_07954_),
    .X(_07989_));
 sky130_fd_sc_hd__clkbuf_1 _14821_ (.A(_07989_),
    .X(_00393_));
 sky130_fd_sc_hd__nor2_1 _14822_ (.A(_07972_),
    .B(_07966_),
    .Y(_07990_));
 sky130_fd_sc_hd__nor2_1 _14823_ (.A(_07969_),
    .B(_07967_),
    .Y(_07991_));
 sky130_fd_sc_hd__o22ai_1 _14824_ (.A1(_06692_),
    .A2(_07990_),
    .B1(_07991_),
    .B2(_06754_),
    .Y(_07992_));
 sky130_fd_sc_hd__xnor2_1 _14825_ (.A(_07517_),
    .B(_07909_),
    .Y(_07993_));
 sky130_fd_sc_hd__nor2_1 _14826_ (.A(_07931_),
    .B(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__a211o_1 _14827_ (.A1(_07931_),
    .A2(_07911_),
    .B1(_07994_),
    .C1(_06792_),
    .X(_07995_));
 sky130_fd_sc_hd__a21oi_1 _14828_ (.A1(_07931_),
    .A2(_07924_),
    .B1(_07973_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_1 _14829_ (.A(_06792_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__a31o_1 _14830_ (.A1(_06751_),
    .A2(_07995_),
    .A3(_07997_),
    .B1(_06602_),
    .X(_07998_));
 sky130_fd_sc_hd__or2_1 _14831_ (.A(_07957_),
    .B(_07960_),
    .X(_07999_));
 sky130_fd_sc_hd__a21o_1 _14832_ (.A1(_06708_),
    .A2(_07999_),
    .B1(_06661_),
    .X(_08000_));
 sky130_fd_sc_hd__o211ai_2 _14833_ (.A1(_07992_),
    .A2(_07998_),
    .B1(_08000_),
    .C1(_06545_),
    .Y(_08001_));
 sky130_fd_sc_hd__nand2_1 _14834_ (.A(_06739_),
    .B(_07970_),
    .Y(_08002_));
 sky130_fd_sc_hd__nor2_1 _14835_ (.A(_06698_),
    .B(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__a21oi_1 _14836_ (.A1(_06675_),
    .A2(_08003_),
    .B1(_07950_),
    .Y(_08004_));
 sky130_fd_sc_hd__nand2_2 _14837_ (.A(_08001_),
    .B(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__mux2_1 _14838_ (.A0(\rbzero.wall_tracer.stepDistY[-8] ),
    .A1(_08005_),
    .S(_07954_),
    .X(_08006_));
 sky130_fd_sc_hd__clkbuf_1 _14839_ (.A(_08006_),
    .X(_00394_));
 sky130_fd_sc_hd__nand3_1 _14840_ (.A(_06751_),
    .B(_07921_),
    .C(_07926_),
    .Y(_08007_));
 sky130_fd_sc_hd__a21oi_1 _14841_ (.A1(_06606_),
    .A2(_07942_),
    .B1(_06602_),
    .Y(_08008_));
 sky130_fd_sc_hd__nand2_1 _14842_ (.A(_06708_),
    .B(_07927_),
    .Y(_08009_));
 sky130_fd_sc_hd__a21o_1 _14843_ (.A1(_06602_),
    .A2(_08009_),
    .B1(_06695_),
    .X(_08010_));
 sky130_fd_sc_hd__a21o_1 _14844_ (.A1(_08007_),
    .A2(_08008_),
    .B1(_08010_),
    .X(_08011_));
 sky130_fd_sc_hd__buf_2 _14845_ (.A(_06673_),
    .X(_08012_));
 sky130_fd_sc_hd__clkinv_2 _14846_ (.A(_07946_),
    .Y(_08013_));
 sky130_fd_sc_hd__nand2_1 _14847_ (.A(_07937_),
    .B(_07944_),
    .Y(_08014_));
 sky130_fd_sc_hd__mux2_1 _14848_ (.A0(_08013_),
    .A1(_08014_),
    .S(_06739_),
    .X(_08015_));
 sky130_fd_sc_hd__a31oi_2 _14849_ (.A1(_06695_),
    .A2(_08012_),
    .A3(_08015_),
    .B1(_07950_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand2_2 _14850_ (.A(_08011_),
    .B(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__mux2_1 _14851_ (.A0(\rbzero.wall_tracer.stepDistY[-7] ),
    .A1(_08017_),
    .S(_07954_),
    .X(_08018_));
 sky130_fd_sc_hd__clkbuf_1 _14852_ (.A(_08018_),
    .X(_00395_));
 sky130_fd_sc_hd__nor2_1 _14853_ (.A(_06567_),
    .B(_06578_),
    .Y(_08019_));
 sky130_fd_sc_hd__clkbuf_4 _14854_ (.A(_08019_),
    .X(_08020_));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(_07990_),
    .A1(_07996_),
    .S(_06642_),
    .X(_08021_));
 sky130_fd_sc_hd__or3_1 _14856_ (.A(_06792_),
    .B(_07957_),
    .C(_07960_),
    .X(_08022_));
 sky130_fd_sc_hd__a211o_1 _14857_ (.A1(_07931_),
    .A2(_07911_),
    .B1(_07994_),
    .C1(_06642_),
    .X(_08023_));
 sky130_fd_sc_hd__a21oi_1 _14858_ (.A1(_08022_),
    .A2(_08023_),
    .B1(_06606_),
    .Y(_08024_));
 sky130_fd_sc_hd__nand2_1 _14859_ (.A(_06545_),
    .B(_06661_),
    .Y(_08025_));
 sky130_fd_sc_hd__a211o_1 _14860_ (.A1(_06606_),
    .A2(_08021_),
    .B1(_08024_),
    .C1(_08025_),
    .X(_08026_));
 sky130_fd_sc_hd__mux2_1 _14861_ (.A0(_07968_),
    .A1(_07970_),
    .S(_07959_),
    .X(_08027_));
 sky130_fd_sc_hd__nand2_1 _14862_ (.A(_08012_),
    .B(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__or2_1 _14863_ (.A(_06697_),
    .B(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__nand3_2 _14864_ (.A(_08020_),
    .B(_08026_),
    .C(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__mux2_1 _14865_ (.A0(\rbzero.wall_tracer.stepDistY[-6] ),
    .A1(_08030_),
    .S(_07954_),
    .X(_08031_));
 sky130_fd_sc_hd__clkbuf_1 _14866_ (.A(_08031_),
    .X(_00396_));
 sky130_fd_sc_hd__a21o_1 _14867_ (.A1(_07980_),
    .A2(_07981_),
    .B1(_06606_),
    .X(_08032_));
 sky130_fd_sc_hd__a211o_1 _14868_ (.A1(_06642_),
    .A2(_07925_),
    .B1(_07983_),
    .C1(_06751_),
    .X(_08033_));
 sky130_fd_sc_hd__and2_1 _14869_ (.A(_07985_),
    .B(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__clkinv_2 _14870_ (.A(_08014_),
    .Y(_08035_));
 sky130_fd_sc_hd__o21a_1 _14871_ (.A1(_06845_),
    .A2(_07933_),
    .B1(_07939_),
    .X(_08036_));
 sky130_fd_sc_hd__mux2_1 _14872_ (.A0(_08035_),
    .A1(_08036_),
    .S(_06739_),
    .X(_08037_));
 sky130_fd_sc_hd__o32a_1 _14873_ (.A1(_06606_),
    .A2(_06642_),
    .A3(_07946_),
    .B1(_08037_),
    .B2(_07956_),
    .X(_08038_));
 sky130_fd_sc_hd__o21ai_1 _14874_ (.A1(_06697_),
    .A2(_08038_),
    .B1(_08020_),
    .Y(_08039_));
 sky130_fd_sc_hd__a21oi_4 _14875_ (.A1(_08032_),
    .A2(_08034_),
    .B1(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__nor2_1 _14876_ (.A(\rbzero.wall_tracer.stepDistY[-5] ),
    .B(_07954_),
    .Y(_08041_));
 sky130_fd_sc_hd__a21oi_1 _14877_ (.A1(_07954_),
    .A2(_08040_),
    .B1(_08041_),
    .Y(_00397_));
 sky130_fd_sc_hd__a21o_1 _14878_ (.A1(_07995_),
    .A2(_07997_),
    .B1(_06751_),
    .X(_08042_));
 sky130_fd_sc_hd__o21ai_1 _14879_ (.A1(_07957_),
    .A2(_07960_),
    .B1(_06792_),
    .Y(_08043_));
 sky130_fd_sc_hd__a21oi_1 _14880_ (.A1(_06751_),
    .A2(_08043_),
    .B1(_08025_),
    .Y(_08044_));
 sky130_fd_sc_hd__a211o_1 _14881_ (.A1(_06626_),
    .A2(_07932_),
    .B1(_07972_),
    .C1(_07959_),
    .X(_08045_));
 sky130_fd_sc_hd__o21ai_1 _14882_ (.A1(_06739_),
    .A2(_07968_),
    .B1(_08045_),
    .Y(_08046_));
 sky130_fd_sc_hd__mux2_1 _14883_ (.A0(_08002_),
    .A1(_08046_),
    .S(_08012_),
    .X(_08047_));
 sky130_fd_sc_hd__o21ai_1 _14884_ (.A1(_06697_),
    .A2(_08047_),
    .B1(_08020_),
    .Y(_08048_));
 sky130_fd_sc_hd__a21o_2 _14885_ (.A1(_08042_),
    .A2(_08044_),
    .B1(_08048_),
    .X(_08049_));
 sky130_fd_sc_hd__buf_4 _14886_ (.A(_07953_),
    .X(_08050_));
 sky130_fd_sc_hd__mux2_1 _14887_ (.A0(\rbzero.wall_tracer.stepDistY[-4] ),
    .A1(_08049_),
    .S(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__clkbuf_1 _14888_ (.A(_08051_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _14889_ (.A0(_07924_),
    .A1(_07932_),
    .S(_06845_),
    .X(_08052_));
 sky130_fd_sc_hd__nand2_1 _14890_ (.A(_07959_),
    .B(_08036_),
    .Y(_08053_));
 sky130_fd_sc_hd__o21ai_1 _14891_ (.A1(_07959_),
    .A2(_08052_),
    .B1(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__nand2_1 _14892_ (.A(_07956_),
    .B(_08015_),
    .Y(_08055_));
 sky130_fd_sc_hd__o21a_1 _14893_ (.A1(_07956_),
    .A2(_08054_),
    .B1(_08055_),
    .X(_08056_));
 sky130_fd_sc_hd__o221a_2 _14894_ (.A1(_08025_),
    .A2(_07929_),
    .B1(_08056_),
    .B2(_06697_),
    .C1(_08020_),
    .X(_08057_));
 sky130_fd_sc_hd__nor2_1 _14895_ (.A(\rbzero.wall_tracer.stepDistY[-3] ),
    .B(_07954_),
    .Y(_08058_));
 sky130_fd_sc_hd__a21oi_1 _14896_ (.A1(_07954_),
    .A2(_08057_),
    .B1(_08058_),
    .Y(_00399_));
 sky130_fd_sc_hd__and3_1 _14897_ (.A(_06606_),
    .B(_08022_),
    .C(_08023_),
    .X(_08059_));
 sky130_fd_sc_hd__a21o_1 _14898_ (.A1(_06675_),
    .A2(_07975_),
    .B1(_07949_),
    .X(_08060_));
 sky130_fd_sc_hd__a21o_4 _14899_ (.A1(_07985_),
    .A2(_08059_),
    .B1(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__mux2_1 _14900_ (.A0(\rbzero.wall_tracer.stepDistY[-2] ),
    .A1(_08061_),
    .S(_08050_),
    .X(_08062_));
 sky130_fd_sc_hd__clkbuf_1 _14901_ (.A(_08062_),
    .X(_00400_));
 sky130_fd_sc_hd__nor2_1 _14902_ (.A(_06626_),
    .B(_07993_),
    .Y(_08063_));
 sky130_fd_sc_hd__a211o_1 _14903_ (.A1(_06626_),
    .A2(_07911_),
    .B1(_08063_),
    .C1(_07959_),
    .X(_08064_));
 sky130_fd_sc_hd__or2_1 _14904_ (.A(_06739_),
    .B(_08052_),
    .X(_08065_));
 sky130_fd_sc_hd__nor2_1 _14905_ (.A(_08012_),
    .B(_08037_),
    .Y(_08066_));
 sky130_fd_sc_hd__a311o_1 _14906_ (.A1(_08012_),
    .A2(_08064_),
    .A3(_08065_),
    .B1(_08066_),
    .C1(_07963_),
    .X(_08067_));
 sky130_fd_sc_hd__a22o_1 _14907_ (.A1(_06661_),
    .A2(_07982_),
    .B1(_08067_),
    .B2(_06675_),
    .X(_08068_));
 sky130_fd_sc_hd__or2_4 _14908_ (.A(_07950_),
    .B(_08068_),
    .X(_08069_));
 sky130_fd_sc_hd__mux2_1 _14909_ (.A0(\rbzero.wall_tracer.stepDistY[-1] ),
    .A1(_08069_),
    .S(_08050_),
    .X(_08070_));
 sky130_fd_sc_hd__clkbuf_1 _14910_ (.A(_08070_),
    .X(_00401_));
 sky130_fd_sc_hd__a211o_1 _14911_ (.A1(_07931_),
    .A2(_07911_),
    .B1(_07957_),
    .C1(_07959_),
    .X(_08071_));
 sky130_fd_sc_hd__or2_1 _14912_ (.A(_06739_),
    .B(_07971_),
    .X(_08072_));
 sky130_fd_sc_hd__nor2_1 _14913_ (.A(_08012_),
    .B(_08046_),
    .Y(_08073_));
 sky130_fd_sc_hd__a31o_1 _14914_ (.A1(_08012_),
    .A2(_08071_),
    .A3(_08072_),
    .B1(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__nor2_2 _14915_ (.A(_06545_),
    .B(_07965_),
    .Y(_08075_));
 sky130_fd_sc_hd__a21o_1 _14916_ (.A1(_08075_),
    .A2(_08003_),
    .B1(_07949_),
    .X(_08076_));
 sky130_fd_sc_hd__a31o_1 _14917_ (.A1(_06661_),
    .A2(_06708_),
    .A3(_07999_),
    .B1(_08076_),
    .X(_08077_));
 sky130_fd_sc_hd__a21o_2 _14918_ (.A1(_06675_),
    .A2(_08074_),
    .B1(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__mux2_1 _14919_ (.A0(\rbzero.wall_tracer.stepDistY[0] ),
    .A1(_08078_),
    .S(_08050_),
    .X(_08079_));
 sky130_fd_sc_hd__clkbuf_1 _14920_ (.A(_08079_),
    .X(_00402_));
 sky130_fd_sc_hd__nor2_1 _14921_ (.A(_07931_),
    .B(_07918_),
    .Y(_08080_));
 sky130_fd_sc_hd__a211o_1 _14922_ (.A1(_06626_),
    .A2(_07911_),
    .B1(_08063_),
    .C1(_06739_),
    .X(_08081_));
 sky130_fd_sc_hd__o31ai_4 _14923_ (.A1(_07959_),
    .A2(_08080_),
    .A3(_07920_),
    .B1(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__mux2_2 _14924_ (.A0(_08082_),
    .A1(_08054_),
    .S(_07956_),
    .X(_08083_));
 sky130_fd_sc_hd__o221ai_4 _14925_ (.A1(_06602_),
    .A2(_08009_),
    .B1(_08083_),
    .B2(_06697_),
    .C1(_08019_),
    .Y(_08084_));
 sky130_fd_sc_hd__mux2_1 _14926_ (.A0(\rbzero.wall_tracer.stepDistY[1] ),
    .A1(_08084_),
    .S(_08050_),
    .X(_08085_));
 sky130_fd_sc_hd__clkbuf_1 _14927_ (.A(_08085_),
    .X(_00403_));
 sky130_fd_sc_hd__inv_2 _14928_ (.A(_08028_),
    .Y(_08086_));
 sky130_fd_sc_hd__and2_1 _14929_ (.A(_07958_),
    .B(_07961_),
    .X(_08087_));
 sky130_fd_sc_hd__mux2_1 _14930_ (.A0(_07971_),
    .A1(_07974_),
    .S(_07959_),
    .X(_08088_));
 sky130_fd_sc_hd__mux2_1 _14931_ (.A0(_08087_),
    .A1(_08088_),
    .S(_07956_),
    .X(_08089_));
 sky130_fd_sc_hd__a221o_4 _14932_ (.A1(_08075_),
    .A2(_08086_),
    .B1(_08089_),
    .B2(_06675_),
    .C1(_07949_),
    .X(_08090_));
 sky130_fd_sc_hd__mux2_1 _14933_ (.A0(\rbzero.wall_tracer.stepDistY[2] ),
    .A1(_08090_),
    .S(_08050_),
    .X(_08091_));
 sky130_fd_sc_hd__clkbuf_1 _14934_ (.A(_08091_),
    .X(_00404_));
 sky130_fd_sc_hd__nand2_1 _14935_ (.A(_07963_),
    .B(_08038_),
    .Y(_08092_));
 sky130_fd_sc_hd__and2_1 _14936_ (.A(_08064_),
    .B(_08065_),
    .X(_08093_));
 sky130_fd_sc_hd__o21a_1 _14937_ (.A1(_08080_),
    .A2(_07920_),
    .B1(_07959_),
    .X(_08094_));
 sky130_fd_sc_hd__a21o_1 _14938_ (.A1(_08012_),
    .A2(_08094_),
    .B1(_07963_),
    .X(_08095_));
 sky130_fd_sc_hd__a21o_1 _14939_ (.A1(_07956_),
    .A2(_08093_),
    .B1(_08095_),
    .X(_08096_));
 sky130_fd_sc_hd__a31o_2 _14940_ (.A1(_06695_),
    .A2(_08092_),
    .A3(_08096_),
    .B1(_07950_),
    .X(_08097_));
 sky130_fd_sc_hd__mux2_1 _14941_ (.A0(\rbzero.wall_tracer.stepDistY[3] ),
    .A1(_08097_),
    .S(_08050_),
    .X(_08098_));
 sky130_fd_sc_hd__clkbuf_1 _14942_ (.A(_08098_),
    .X(_00405_));
 sky130_fd_sc_hd__nand3_1 _14943_ (.A(_07956_),
    .B(_08071_),
    .C(_08072_),
    .Y(_08099_));
 sky130_fd_sc_hd__o41a_1 _14944_ (.A1(_06648_),
    .A2(_06626_),
    .A3(_07956_),
    .A4(_07918_),
    .B1(_07965_),
    .X(_08100_));
 sky130_fd_sc_hd__a22o_1 _14945_ (.A1(_07963_),
    .A2(_08047_),
    .B1(_08099_),
    .B2(_08100_),
    .X(_08101_));
 sky130_fd_sc_hd__o21ai_1 _14946_ (.A1(_06545_),
    .A2(_08101_),
    .B1(_08020_),
    .Y(_08102_));
 sky130_fd_sc_hd__buf_2 _14947_ (.A(_08102_),
    .X(_08103_));
 sky130_fd_sc_hd__mux2_1 _14948_ (.A0(\rbzero.wall_tracer.stepDistY[4] ),
    .A1(_08103_),
    .S(_08050_),
    .X(_08104_));
 sky130_fd_sc_hd__clkbuf_1 _14949_ (.A(_08104_),
    .X(_00406_));
 sky130_fd_sc_hd__nand2_1 _14950_ (.A(_06695_),
    .B(_07956_),
    .Y(_08105_));
 sky130_fd_sc_hd__o221ai_4 _14951_ (.A1(_08105_),
    .A2(_08082_),
    .B1(_08056_),
    .B2(_06795_),
    .C1(_08020_),
    .Y(_08106_));
 sky130_fd_sc_hd__mux2_1 _14952_ (.A0(\rbzero.wall_tracer.stepDistY[5] ),
    .A1(_08106_),
    .S(_08050_),
    .X(_08107_));
 sky130_fd_sc_hd__clkbuf_1 _14953_ (.A(_08107_),
    .X(_00407_));
 sky130_fd_sc_hd__nor2_1 _14954_ (.A(_06545_),
    .B(_08012_),
    .Y(_08108_));
 sky130_fd_sc_hd__a21o_1 _14955_ (.A1(_08075_),
    .A2(_07975_),
    .B1(_07950_),
    .X(_08109_));
 sky130_fd_sc_hd__a21o_1 _14956_ (.A1(_08108_),
    .A2(_08087_),
    .B1(_08109_),
    .X(_08110_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(\rbzero.wall_tracer.stepDistY[6] ),
    .A1(_08110_),
    .S(_08050_),
    .X(_08111_));
 sky130_fd_sc_hd__clkbuf_1 _14958_ (.A(_08111_),
    .X(_00408_));
 sky130_fd_sc_hd__a211o_1 _14959_ (.A1(_08012_),
    .A2(_08093_),
    .B1(_08066_),
    .C1(_07965_),
    .X(_08112_));
 sky130_fd_sc_hd__a21o_1 _14960_ (.A1(_08108_),
    .A2(_08094_),
    .B1(_08075_),
    .X(_08113_));
 sky130_fd_sc_hd__a21o_1 _14961_ (.A1(_08112_),
    .A2(_08113_),
    .B1(_07950_),
    .X(_08114_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(\rbzero.wall_tracer.stepDistY[7] ),
    .A1(_08114_),
    .S(_07953_),
    .X(_08115_));
 sky130_fd_sc_hd__clkbuf_1 _14963_ (.A(_08115_),
    .X(_00409_));
 sky130_fd_sc_hd__a31o_1 _14964_ (.A1(_06639_),
    .A2(_08108_),
    .A3(_07960_),
    .B1(_08075_),
    .X(_08116_));
 sky130_fd_sc_hd__o21ai_1 _14965_ (.A1(_07965_),
    .A2(_08074_),
    .B1(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__nand2_1 _14966_ (.A(_08020_),
    .B(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__mux2_1 _14967_ (.A0(\rbzero.wall_tracer.stepDistY[8] ),
    .A1(_08118_),
    .S(_07953_),
    .X(_08119_));
 sky130_fd_sc_hd__clkbuf_1 _14968_ (.A(_08119_),
    .X(_00410_));
 sky130_fd_sc_hd__o21ai_2 _14969_ (.A1(_06795_),
    .A2(_08083_),
    .B1(_08020_),
    .Y(_08120_));
 sky130_fd_sc_hd__mux2_1 _14970_ (.A0(\rbzero.wall_tracer.stepDistY[9] ),
    .A1(_08120_),
    .S(_07953_),
    .X(_08121_));
 sky130_fd_sc_hd__clkbuf_1 _14971_ (.A(_08121_),
    .X(_00411_));
 sky130_fd_sc_hd__and3_1 _14972_ (.A(_08020_),
    .B(_08075_),
    .C(_08089_),
    .X(_08122_));
 sky130_fd_sc_hd__mux2_1 _14973_ (.A0(\rbzero.wall_tracer.stepDistY[10] ),
    .A1(_08122_),
    .S(_07953_),
    .X(_08123_));
 sky130_fd_sc_hd__clkbuf_1 _14974_ (.A(_08123_),
    .X(_00412_));
 sky130_fd_sc_hd__clkbuf_4 _14975_ (.A(_06332_),
    .X(_08124_));
 sky130_fd_sc_hd__or3_2 _14976_ (.A(_06162_),
    .B(_06237_),
    .C(_06330_),
    .X(_08125_));
 sky130_fd_sc_hd__clkbuf_4 _14977_ (.A(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__clkbuf_4 _14978_ (.A(_06331_),
    .X(_08127_));
 sky130_fd_sc_hd__buf_4 _14979_ (.A(_04491_),
    .X(_08128_));
 sky130_fd_sc_hd__o21a_1 _14980_ (.A1(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A2(_08127_),
    .B1(_08128_),
    .X(_08129_));
 sky130_fd_sc_hd__o221a_1 _14981_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(_08124_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[-11] ),
    .C1(_08129_),
    .X(_00413_));
 sky130_fd_sc_hd__clkbuf_4 _14982_ (.A(_06332_),
    .X(_08130_));
 sky130_fd_sc_hd__buf_4 _14983_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_08131_));
 sky130_fd_sc_hd__clkbuf_4 _14984_ (.A(_06331_),
    .X(_08132_));
 sky130_fd_sc_hd__clkbuf_4 _14985_ (.A(_08125_),
    .X(_08133_));
 sky130_fd_sc_hd__o221a_1 _14986_ (.A1(_08131_),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[-10] ),
    .C1(_08128_),
    .X(_08134_));
 sky130_fd_sc_hd__o21a_1 _14987_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(_08130_),
    .B1(_08134_),
    .X(_00414_));
 sky130_fd_sc_hd__o22a_1 _14988_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08127_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(_08135_));
 sky130_fd_sc_hd__buf_6 _14989_ (.A(_04491_),
    .X(_08136_));
 sky130_fd_sc_hd__buf_4 _14990_ (.A(_08136_),
    .X(_01633_));
 sky130_fd_sc_hd__o211a_1 _14991_ (.A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .A2(_08130_),
    .B1(_08135_),
    .C1(_01633_),
    .X(_00415_));
 sky130_fd_sc_hd__o221a_1 _14992_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[-8] ),
    .C1(_08128_),
    .X(_08137_));
 sky130_fd_sc_hd__o21a_1 _14993_ (.A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .A2(_08130_),
    .B1(_08137_),
    .X(_00416_));
 sky130_fd_sc_hd__o21a_1 _14994_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_08127_),
    .B1(_08128_),
    .X(_08138_));
 sky130_fd_sc_hd__o221a_1 _14995_ (.A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .A2(_08124_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[-7] ),
    .C1(_08138_),
    .X(_00417_));
 sky130_fd_sc_hd__o22a_1 _14996_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_08127_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(_08139_));
 sky130_fd_sc_hd__o211a_1 _14997_ (.A1(\rbzero.wall_tracer.trackDistX[-6] ),
    .A2(_08124_),
    .B1(_08139_),
    .C1(_01633_),
    .X(_00418_));
 sky130_fd_sc_hd__o22a_1 _14998_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_08127_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[-5] ),
    .X(_08140_));
 sky130_fd_sc_hd__o211a_1 _14999_ (.A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .A2(_08124_),
    .B1(_08140_),
    .C1(_01633_),
    .X(_00419_));
 sky130_fd_sc_hd__o221a_1 _15000_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[-4] ),
    .C1(_08128_),
    .X(_08141_));
 sky130_fd_sc_hd__o21a_1 _15001_ (.A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .A2(_08130_),
    .B1(_08141_),
    .X(_00420_));
 sky130_fd_sc_hd__o21a_1 _15002_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_08127_),
    .B1(_08128_),
    .X(_08142_));
 sky130_fd_sc_hd__o221a_1 _15003_ (.A1(\rbzero.wall_tracer.trackDistX[-3] ),
    .A2(_08124_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[-3] ),
    .C1(_08142_),
    .X(_00421_));
 sky130_fd_sc_hd__o22a_1 _15004_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_08132_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_08143_));
 sky130_fd_sc_hd__o211a_1 _15005_ (.A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .A2(_08124_),
    .B1(_08143_),
    .C1(_01633_),
    .X(_00422_));
 sky130_fd_sc_hd__o221a_1 _15006_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[-1] ),
    .C1(_08136_),
    .X(_08144_));
 sky130_fd_sc_hd__o21a_1 _15007_ (.A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .A2(_08130_),
    .B1(_08144_),
    .X(_00423_));
 sky130_fd_sc_hd__o22a_1 _15008_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_08132_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[0] ),
    .X(_08145_));
 sky130_fd_sc_hd__o211a_1 _15009_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(_08124_),
    .B1(_08145_),
    .C1(_01633_),
    .X(_00424_));
 sky130_fd_sc_hd__o22a_1 _15010_ (.A1(\rbzero.wall_tracer.visualWallDist[1] ),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[1] ),
    .X(_08146_));
 sky130_fd_sc_hd__o211a_1 _15011_ (.A1(\rbzero.wall_tracer.trackDistX[1] ),
    .A2(_08124_),
    .B1(_08146_),
    .C1(_01633_),
    .X(_00425_));
 sky130_fd_sc_hd__o221a_1 _15012_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[2] ),
    .C1(_08136_),
    .X(_08147_));
 sky130_fd_sc_hd__o21a_1 _15013_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_08130_),
    .B1(_08147_),
    .X(_00426_));
 sky130_fd_sc_hd__o221a_1 _15014_ (.A1(\rbzero.wall_tracer.visualWallDist[3] ),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[3] ),
    .C1(_08136_),
    .X(_08148_));
 sky130_fd_sc_hd__o21a_1 _15015_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_08130_),
    .B1(_08148_),
    .X(_00427_));
 sky130_fd_sc_hd__o221a_1 _15016_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_06331_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[4] ),
    .C1(_08136_),
    .X(_08149_));
 sky130_fd_sc_hd__o21a_1 _15017_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(_08130_),
    .B1(_08149_),
    .X(_00428_));
 sky130_fd_sc_hd__o221a_1 _15018_ (.A1(\rbzero.wall_tracer.visualWallDist[5] ),
    .A2(_06331_),
    .B1(_08125_),
    .B2(\rbzero.wall_tracer.trackDistY[5] ),
    .C1(_08136_),
    .X(_08150_));
 sky130_fd_sc_hd__o21a_1 _15019_ (.A1(\rbzero.wall_tracer.trackDistX[5] ),
    .A2(_08130_),
    .B1(_08150_),
    .X(_00429_));
 sky130_fd_sc_hd__o21a_1 _15020_ (.A1(\rbzero.wall_tracer.visualWallDist[6] ),
    .A2(_08127_),
    .B1(_08128_),
    .X(_08151_));
 sky130_fd_sc_hd__o221a_1 _15021_ (.A1(\rbzero.wall_tracer.trackDistX[6] ),
    .A2(_08124_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[6] ),
    .C1(_08151_),
    .X(_00430_));
 sky130_fd_sc_hd__o22a_1 _15022_ (.A1(\rbzero.wall_tracer.visualWallDist[7] ),
    .A2(_08132_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[7] ),
    .X(_08152_));
 sky130_fd_sc_hd__o211a_1 _15023_ (.A1(\rbzero.wall_tracer.trackDistX[7] ),
    .A2(_08124_),
    .B1(_08152_),
    .C1(_01633_),
    .X(_00431_));
 sky130_fd_sc_hd__o22a_1 _15024_ (.A1(\rbzero.wall_tracer.trackDistX[8] ),
    .A2(_06332_),
    .B1(_08133_),
    .B2(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_08153_));
 sky130_fd_sc_hd__o211a_1 _15025_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_08127_),
    .B1(_08153_),
    .C1(_01633_),
    .X(_00432_));
 sky130_fd_sc_hd__o21a_1 _15026_ (.A1(\rbzero.wall_tracer.visualWallDist[9] ),
    .A2(_08127_),
    .B1(_08128_),
    .X(_08154_));
 sky130_fd_sc_hd__o221a_1 _15027_ (.A1(\rbzero.wall_tracer.trackDistX[9] ),
    .A2(_06332_),
    .B1(_08126_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .C1(_08154_),
    .X(_00433_));
 sky130_fd_sc_hd__buf_6 _15028_ (.A(_06162_),
    .X(_08155_));
 sky130_fd_sc_hd__clkbuf_8 _15029_ (.A(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__o21a_1 _15030_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(_06236_),
    .B1(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_08157_));
 sky130_fd_sc_hd__or2_1 _15031_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_06331_),
    .X(_08158_));
 sky130_fd_sc_hd__o311a_1 _15032_ (.A1(_08156_),
    .A2(_06330_),
    .A3(_08157_),
    .B1(_08158_),
    .C1(_04500_),
    .X(_00434_));
 sky130_fd_sc_hd__and4b_1 _15033_ (.A_N(_04495_),
    .B(_04490_),
    .C(_04496_),
    .D(_04493_),
    .X(_08159_));
 sky130_fd_sc_hd__clkbuf_4 _15034_ (.A(_08159_),
    .X(_08160_));
 sky130_fd_sc_hd__clkbuf_4 _15035_ (.A(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__mux2_1 _15036_ (.A0(\rbzero.wall_tracer.stepDistX[-11] ),
    .A1(_07951_),
    .S(_08161_),
    .X(_08162_));
 sky130_fd_sc_hd__clkbuf_1 _15037_ (.A(_08162_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _15038_ (.A0(\rbzero.wall_tracer.stepDistX[-10] ),
    .A1(_07977_),
    .S(_08161_),
    .X(_08163_));
 sky130_fd_sc_hd__clkbuf_1 _15039_ (.A(_08163_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _15040_ (.A0(\rbzero.wall_tracer.stepDistX[-9] ),
    .A1(_07988_),
    .S(_08161_),
    .X(_08164_));
 sky130_fd_sc_hd__clkbuf_1 _15041_ (.A(_08164_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _15042_ (.A0(\rbzero.wall_tracer.stepDistX[-8] ),
    .A1(_08005_),
    .S(_08161_),
    .X(_08165_));
 sky130_fd_sc_hd__clkbuf_1 _15043_ (.A(_08165_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _15044_ (.A0(\rbzero.wall_tracer.stepDistX[-7] ),
    .A1(_08017_),
    .S(_08161_),
    .X(_08166_));
 sky130_fd_sc_hd__clkbuf_1 _15045_ (.A(_08166_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _15046_ (.A0(\rbzero.wall_tracer.stepDistX[-6] ),
    .A1(_08030_),
    .S(_08161_),
    .X(_08167_));
 sky130_fd_sc_hd__clkbuf_1 _15047_ (.A(_08167_),
    .X(_00440_));
 sky130_fd_sc_hd__nor2_1 _15048_ (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(_08161_),
    .Y(_08168_));
 sky130_fd_sc_hd__a21oi_1 _15049_ (.A1(_08040_),
    .A2(_08161_),
    .B1(_08168_),
    .Y(_00441_));
 sky130_fd_sc_hd__buf_4 _15050_ (.A(_08160_),
    .X(_08169_));
 sky130_fd_sc_hd__mux2_1 _15051_ (.A0(\rbzero.wall_tracer.stepDistX[-4] ),
    .A1(_08049_),
    .S(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__clkbuf_1 _15052_ (.A(_08170_),
    .X(_00442_));
 sky130_fd_sc_hd__nor2_1 _15053_ (.A(\rbzero.wall_tracer.stepDistX[-3] ),
    .B(_08161_),
    .Y(_08171_));
 sky130_fd_sc_hd__a21oi_1 _15054_ (.A1(_08057_),
    .A2(_08161_),
    .B1(_08171_),
    .Y(_00443_));
 sky130_fd_sc_hd__mux2_1 _15055_ (.A0(\rbzero.wall_tracer.stepDistX[-2] ),
    .A1(_08061_),
    .S(_08169_),
    .X(_08172_));
 sky130_fd_sc_hd__clkbuf_1 _15056_ (.A(_08172_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _15057_ (.A0(\rbzero.wall_tracer.stepDistX[-1] ),
    .A1(_08069_),
    .S(_08169_),
    .X(_08173_));
 sky130_fd_sc_hd__clkbuf_1 _15058_ (.A(_08173_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _15059_ (.A0(\rbzero.wall_tracer.stepDistX[0] ),
    .A1(_08078_),
    .S(_08169_),
    .X(_08174_));
 sky130_fd_sc_hd__clkbuf_1 _15060_ (.A(_08174_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _15061_ (.A0(\rbzero.wall_tracer.stepDistX[1] ),
    .A1(_08084_),
    .S(_08169_),
    .X(_08175_));
 sky130_fd_sc_hd__clkbuf_1 _15062_ (.A(_08175_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _15063_ (.A0(\rbzero.wall_tracer.stepDistX[2] ),
    .A1(_08090_),
    .S(_08169_),
    .X(_08176_));
 sky130_fd_sc_hd__clkbuf_1 _15064_ (.A(_08176_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _15065_ (.A0(\rbzero.wall_tracer.stepDistX[3] ),
    .A1(_08097_),
    .S(_08169_),
    .X(_08177_));
 sky130_fd_sc_hd__clkbuf_1 _15066_ (.A(_08177_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _15067_ (.A0(\rbzero.wall_tracer.stepDistX[4] ),
    .A1(_08103_),
    .S(_08169_),
    .X(_08178_));
 sky130_fd_sc_hd__clkbuf_1 _15068_ (.A(_08178_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _15069_ (.A0(\rbzero.wall_tracer.stepDistX[5] ),
    .A1(_08106_),
    .S(_08169_),
    .X(_08179_));
 sky130_fd_sc_hd__clkbuf_1 _15070_ (.A(_08179_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _15071_ (.A0(\rbzero.wall_tracer.stepDistX[6] ),
    .A1(_08110_),
    .S(_08169_),
    .X(_08180_));
 sky130_fd_sc_hd__clkbuf_1 _15072_ (.A(_08180_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _15073_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_08114_),
    .S(_08160_),
    .X(_08181_));
 sky130_fd_sc_hd__clkbuf_1 _15074_ (.A(_08181_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _15075_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_08118_),
    .S(_08160_),
    .X(_08182_));
 sky130_fd_sc_hd__clkbuf_1 _15076_ (.A(_08182_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _15077_ (.A0(\rbzero.wall_tracer.stepDistX[9] ),
    .A1(_08120_),
    .S(_08160_),
    .X(_08183_));
 sky130_fd_sc_hd__clkbuf_1 _15078_ (.A(_08183_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _15079_ (.A0(\rbzero.wall_tracer.stepDistX[10] ),
    .A1(_08122_),
    .S(_08160_),
    .X(_08184_));
 sky130_fd_sc_hd__clkbuf_1 _15080_ (.A(_08184_),
    .X(_00456_));
 sky130_fd_sc_hd__nor2_1 _15081_ (.A(net64),
    .B(_05779_),
    .Y(_00457_));
 sky130_fd_sc_hd__nor2_1 _15082_ (.A(net64),
    .B(_05363_),
    .Y(_00458_));
 sky130_fd_sc_hd__buf_4 _15083_ (.A(_04112_),
    .X(_08185_));
 sky130_fd_sc_hd__clkbuf_4 _15084_ (.A(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__and2_1 _15085_ (.A(_08186_),
    .B(_05450_),
    .X(_08187_));
 sky130_fd_sc_hd__clkbuf_1 _15086_ (.A(_08187_),
    .X(_00459_));
 sky130_fd_sc_hd__and2_1 _15087_ (.A(_08186_),
    .B(_05539_),
    .X(_08188_));
 sky130_fd_sc_hd__clkbuf_1 _15088_ (.A(_08188_),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _15089_ (.A(_08186_),
    .B(_05629_),
    .X(_08189_));
 sky130_fd_sc_hd__clkbuf_1 _15090_ (.A(_08189_),
    .X(_00461_));
 sky130_fd_sc_hd__buf_2 _15091_ (.A(_04112_),
    .X(_08190_));
 sky130_fd_sc_hd__and2_1 _15092_ (.A(_08190_),
    .B(_05710_),
    .X(_08191_));
 sky130_fd_sc_hd__clkbuf_1 _15093_ (.A(_08191_),
    .X(_00462_));
 sky130_fd_sc_hd__nor3b_4 _15094_ (.A(_04486_),
    .B(_04487_),
    .C_N(\rbzero.trace_state[3] ),
    .Y(_08192_));
 sky130_fd_sc_hd__buf_6 _15095_ (.A(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__buf_8 _15096_ (.A(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__buf_8 _15097_ (.A(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__nand2_4 _15098_ (.A(_08195_),
    .B(_06330_),
    .Y(_08196_));
 sky130_fd_sc_hd__o21bai_1 _15099_ (.A1(_06272_),
    .A2(_06321_),
    .B1_N(_06280_),
    .Y(_08197_));
 sky130_fd_sc_hd__a2bb2o_1 _15100_ (.A1_N(_06305_),
    .A2_N(_08197_),
    .B1(\rbzero.mapdyw[0] ),
    .B2(_06280_),
    .X(_08198_));
 sky130_fd_sc_hd__mux2_1 _15101_ (.A0(_08198_),
    .A1(\rbzero.mapdxw[0] ),
    .S(_06291_),
    .X(_08199_));
 sky130_fd_sc_hd__buf_4 _15102_ (.A(_04489_),
    .X(_08200_));
 sky130_fd_sc_hd__buf_6 _15103_ (.A(_08200_),
    .X(_08201_));
 sky130_fd_sc_hd__a21oi_1 _15104_ (.A1(_04519_),
    .A2(_08196_),
    .B1(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__o21a_1 _15105_ (.A1(_08196_),
    .A2(_08199_),
    .B1(_08202_),
    .X(_00463_));
 sky130_fd_sc_hd__a2bb2o_1 _15106_ (.A1_N(_06328_),
    .A2_N(_08197_),
    .B1(\rbzero.mapdyw[1] ),
    .B2(_06280_),
    .X(_08203_));
 sky130_fd_sc_hd__mux2_1 _15107_ (.A0(_08203_),
    .A1(\rbzero.mapdxw[1] ),
    .S(_06291_),
    .X(_08204_));
 sky130_fd_sc_hd__a21oi_1 _15108_ (.A1(_04604_),
    .A2(_08196_),
    .B1(_08201_),
    .Y(_08205_));
 sky130_fd_sc_hd__o21a_1 _15109_ (.A1(_08196_),
    .A2(_08204_),
    .B1(_08205_),
    .X(_00464_));
 sky130_fd_sc_hd__buf_4 _15110_ (.A(_04536_),
    .X(_08206_));
 sky130_fd_sc_hd__o211a_1 _15111_ (.A1(_08206_),
    .A2(_08127_),
    .B1(_08130_),
    .C1(_04500_),
    .X(_00465_));
 sky130_fd_sc_hd__nand2_1 _15112_ (.A(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .Y(_08207_));
 sky130_fd_sc_hd__nor2_2 _15113_ (.A(_04487_),
    .B(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__buf_4 _15114_ (.A(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__buf_4 _15115_ (.A(_08209_),
    .X(_08210_));
 sky130_fd_sc_hd__clkbuf_4 _15116_ (.A(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__or2_1 _15117_ (.A(_04487_),
    .B(_08207_),
    .X(_08212_));
 sky130_fd_sc_hd__clkbuf_4 _15118_ (.A(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__buf_4 _15119_ (.A(_08213_),
    .X(_08214_));
 sky130_fd_sc_hd__and3_2 _15120_ (.A(_04493_),
    .B(\rbzero.trace_state[0] ),
    .C(_06335_),
    .X(_08215_));
 sky130_fd_sc_hd__buf_6 _15121_ (.A(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__o31a_2 _15122_ (.A1(_07949_),
    .A2(_08061_),
    .A3(_08068_),
    .B1(_08078_),
    .X(_08217_));
 sky130_fd_sc_hd__nor4_1 _15123_ (.A(_07950_),
    .B(_08061_),
    .C(_08068_),
    .D(_08078_),
    .Y(_08218_));
 sky130_fd_sc_hd__o21ai_1 _15124_ (.A1(_08217_),
    .A2(_08218_),
    .B1(_08214_),
    .Y(_08219_));
 sky130_fd_sc_hd__clkinv_2 _15125_ (.A(_06477_),
    .Y(_08220_));
 sky130_fd_sc_hd__mux2_1 _15126_ (.A0(_06106_),
    .A1(_08220_),
    .S(_04535_),
    .X(_08221_));
 sky130_fd_sc_hd__and2_1 _15127_ (.A(\rbzero.trace_state[1] ),
    .B(_06335_),
    .X(_08222_));
 sky130_fd_sc_hd__clkbuf_8 _15128_ (.A(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__nand2_1 _15129_ (.A(_04494_),
    .B(_08223_),
    .Y(_08224_));
 sky130_fd_sc_hd__buf_4 _15130_ (.A(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__o21a_1 _15131_ (.A1(_08213_),
    .A2(_08221_),
    .B1(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__a22o_1 _15132_ (.A1(\rbzero.wall_tracer.stepDistY[0] ),
    .A2(_08216_),
    .B1(_08219_),
    .B2(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__clkbuf_4 _15133_ (.A(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__nor2_1 _15134_ (.A(_04494_),
    .B(_06336_),
    .Y(_08229_));
 sky130_fd_sc_hd__buf_6 _15135_ (.A(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__buf_4 _15136_ (.A(_08230_),
    .X(_08231_));
 sky130_fd_sc_hd__and2_1 _15137_ (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .B(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__a21oi_4 _15138_ (.A1(_06340_),
    .A2(_08228_),
    .B1(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__buf_6 _15139_ (.A(_06336_),
    .X(_08234_));
 sky130_fd_sc_hd__xor2_1 _15140_ (.A(_08061_),
    .B(_08069_),
    .X(_08235_));
 sky130_fd_sc_hd__nor2_1 _15141_ (.A(_04535_),
    .B(_06114_),
    .Y(_08236_));
 sky130_fd_sc_hd__a211o_1 _15142_ (.A1(_04535_),
    .A2(_06484_),
    .B1(_08213_),
    .C1(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__o21ai_4 _15143_ (.A1(_08209_),
    .A2(_08235_),
    .B1(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__clkbuf_8 _15144_ (.A(_08223_),
    .X(_08239_));
 sky130_fd_sc_hd__and3_2 _15145_ (.A(_04494_),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .C(_08239_),
    .X(_08240_));
 sky130_fd_sc_hd__nand2_1 _15146_ (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .B(_08230_),
    .Y(_08241_));
 sky130_fd_sc_hd__inv_2 _15147_ (.A(_08241_),
    .Y(_08242_));
 sky130_fd_sc_hd__a211oi_4 _15148_ (.A1(_08234_),
    .A2(_08238_),
    .B1(_08240_),
    .C1(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__clkbuf_4 _15149_ (.A(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__or3_1 _15150_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(\rbzero.debug_overlay.playerX[-8] ),
    .C(\rbzero.debug_overlay.playerX[-9] ),
    .X(_08245_));
 sky130_fd_sc_hd__o21ai_1 _15151_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(\rbzero.debug_overlay.playerX[-9] ),
    .B1(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_08246_));
 sky130_fd_sc_hd__and2_1 _15152_ (.A(_08245_),
    .B(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__nor4_1 _15153_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .C(_06463_),
    .D(_06454_),
    .Y(_08248_));
 sky130_fd_sc_hd__and4b_1 _15154_ (.A_N(_06470_),
    .B(_06440_),
    .C(_06449_),
    .D(_08248_),
    .X(_08249_));
 sky130_fd_sc_hd__and4_1 _15155_ (.A(_06484_),
    .B(_06431_),
    .C(_06436_),
    .D(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__and4_1 _15156_ (.A(_06419_),
    .B(_06477_),
    .C(_06427_),
    .D(_08250_),
    .X(_08251_));
 sky130_fd_sc_hd__a21bo_2 _15157_ (.A1(_06414_),
    .A2(_08251_),
    .B1_N(_06403_),
    .X(_08252_));
 sky130_fd_sc_hd__mux2_1 _15158_ (.A0(_08247_),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__or3_1 _15159_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(\rbzero.debug_overlay.playerY[-8] ),
    .C(\rbzero.debug_overlay.playerY[-9] ),
    .X(_08254_));
 sky130_fd_sc_hd__o21ai_1 _15160_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(\rbzero.debug_overlay.playerY[-9] ),
    .B1(\rbzero.debug_overlay.playerY[-7] ),
    .Y(_08255_));
 sky130_fd_sc_hd__a21o_1 _15161_ (.A1(_08254_),
    .A2(_08255_),
    .B1(_06146_),
    .X(_08256_));
 sky130_fd_sc_hd__o211a_1 _15162_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_06135_),
    .B1(_08215_),
    .C1(_08256_),
    .X(_08257_));
 sky130_fd_sc_hd__a211o_1 _15163_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_08225_),
    .B1(_08257_),
    .C1(_08229_),
    .X(_08258_));
 sky130_fd_sc_hd__o21ai_4 _15164_ (.A1(_06338_),
    .A2(_08253_),
    .B1(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__inv_2 _15165_ (.A(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__xor2_1 _15166_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(\rbzero.debug_overlay.playerX[-9] ),
    .X(_08261_));
 sky130_fd_sc_hd__mux2_2 _15167_ (.A0(_08261_),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_08252_),
    .X(_08262_));
 sky130_fd_sc_hd__xor2_1 _15168_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(\rbzero.debug_overlay.playerY[-9] ),
    .X(_08263_));
 sky130_fd_sc_hd__mux2_1 _15169_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(_08263_),
    .S(_06135_),
    .X(_08264_));
 sky130_fd_sc_hd__or2_1 _15170_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_08222_),
    .X(_08265_));
 sky130_fd_sc_hd__mux2_1 _15171_ (.A0(_08264_),
    .A1(_08265_),
    .S(_08224_),
    .X(_08266_));
 sky130_fd_sc_hd__o21ai_4 _15172_ (.A1(_06338_),
    .A2(_08262_),
    .B1(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__buf_2 _15173_ (.A(_08267_),
    .X(_08268_));
 sky130_fd_sc_hd__clkinv_2 _15174_ (.A(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__and4bb_1 _15175_ (.A_N(_08233_),
    .B_N(_08244_),
    .C(_08260_),
    .D(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__clkbuf_4 _15176_ (.A(_08268_),
    .X(_08271_));
 sky130_fd_sc_hd__clkbuf_4 _15177_ (.A(_08259_),
    .X(_08272_));
 sky130_fd_sc_hd__o22a_1 _15178_ (.A1(_08271_),
    .A2(_08233_),
    .B1(_08244_),
    .B2(_08272_),
    .X(_08273_));
 sky130_fd_sc_hd__or2_1 _15179_ (.A(_08270_),
    .B(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__inv_2 _15180_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .Y(_08275_));
 sky130_fd_sc_hd__or2_1 _15181_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08254_),
    .X(_08276_));
 sky130_fd_sc_hd__nand2_1 _15182_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08254_),
    .Y(_08277_));
 sky130_fd_sc_hd__nand2_1 _15183_ (.A(_08276_),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__mux2_1 _15184_ (.A0(_08275_),
    .A1(_08278_),
    .S(_06136_),
    .X(_08279_));
 sky130_fd_sc_hd__mux2_1 _15185_ (.A0(_06445_),
    .A1(_08279_),
    .S(_08216_),
    .X(_08280_));
 sky130_fd_sc_hd__or2_1 _15186_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08245_),
    .X(_08281_));
 sky130_fd_sc_hd__nand2_1 _15187_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08245_),
    .Y(_08282_));
 sky130_fd_sc_hd__nand2_1 _15188_ (.A(_08281_),
    .B(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__inv_2 _15189_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .Y(_08284_));
 sky130_fd_sc_hd__buf_4 _15190_ (.A(_08252_),
    .X(_08285_));
 sky130_fd_sc_hd__mux2_1 _15191_ (.A0(_08283_),
    .A1(_08284_),
    .S(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__mux2_4 _15192_ (.A0(_08280_),
    .A1(_08286_),
    .S(_08230_),
    .X(_08287_));
 sky130_fd_sc_hd__buf_2 _15193_ (.A(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__clkinv_2 _15194_ (.A(_06133_),
    .Y(_08289_));
 sky130_fd_sc_hd__mux2_1 _15195_ (.A0(_08289_),
    .A1(_06427_),
    .S(\rbzero.side_hot ),
    .X(_08290_));
 sky130_fd_sc_hd__a21o_1 _15196_ (.A1(_08208_),
    .A2(_08290_),
    .B1(_08223_),
    .X(_08291_));
 sky130_fd_sc_hd__a21oi_4 _15197_ (.A1(_08061_),
    .A2(_08213_),
    .B1(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__a21oi_4 _15198_ (.A1(\rbzero.wall_tracer.stepDistY[-2] ),
    .A2(_08216_),
    .B1(_08292_),
    .Y(_08293_));
 sky130_fd_sc_hd__a21boi_2 _15199_ (.A1(\rbzero.wall_tracer.stepDistX[-2] ),
    .A2(_08230_),
    .B1_N(_08293_),
    .Y(_08294_));
 sky130_fd_sc_hd__clkbuf_4 _15200_ (.A(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__nor2_1 _15201_ (.A(_08288_),
    .B(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__xnor2_2 _15202_ (.A(_08274_),
    .B(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__clkbuf_4 _15203_ (.A(_08239_),
    .X(_08298_));
 sky130_fd_sc_hd__xnor2_1 _15204_ (.A(_08084_),
    .B(_08217_),
    .Y(_08299_));
 sky130_fd_sc_hd__nand2_1 _15205_ (.A(_04536_),
    .B(_06419_),
    .Y(_08300_));
 sky130_fd_sc_hd__o211a_1 _15206_ (.A1(_04536_),
    .A2(_06103_),
    .B1(_08210_),
    .C1(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__a21oi_2 _15207_ (.A1(_08214_),
    .A2(_08299_),
    .B1(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__clkbuf_4 _15208_ (.A(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__buf_6 _15209_ (.A(_08216_),
    .X(_08304_));
 sky130_fd_sc_hd__a22o_1 _15210_ (.A1(\rbzero.wall_tracer.stepDistX[1] ),
    .A2(_08231_),
    .B1(_08304_),
    .B2(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_08305_));
 sky130_fd_sc_hd__o21ba_1 _15211_ (.A1(_08298_),
    .A2(_08303_),
    .B1_N(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__buf_2 _15212_ (.A(_08306_),
    .X(_08307_));
 sky130_fd_sc_hd__inv_2 _15213_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_08308_));
 sky130_fd_sc_hd__buf_6 _15214_ (.A(_08225_),
    .X(_08309_));
 sky130_fd_sc_hd__nor2_2 _15215_ (.A(_08308_),
    .B(_08309_),
    .Y(_08310_));
 sky130_fd_sc_hd__a221oi_4 _15216_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08234_),
    .B1(_08230_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__buf_2 _15217_ (.A(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__nor2_1 _15218_ (.A(_08307_),
    .B(_08312_),
    .Y(_08313_));
 sky130_fd_sc_hd__clkinv_2 _15219_ (.A(_08131_),
    .Y(_08314_));
 sky130_fd_sc_hd__nor2_1 _15220_ (.A(_04536_),
    .B(_06098_),
    .Y(_08315_));
 sky130_fd_sc_hd__a211o_2 _15221_ (.A1(_04536_),
    .A2(_06414_),
    .B1(_08214_),
    .C1(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__or3_1 _15222_ (.A(_08084_),
    .B(_08090_),
    .C(_08217_),
    .X(_08317_));
 sky130_fd_sc_hd__o21ai_1 _15223_ (.A1(_08084_),
    .A2(_08217_),
    .B1(_08090_),
    .Y(_08318_));
 sky130_fd_sc_hd__a21o_1 _15224_ (.A1(_08317_),
    .A2(_08318_),
    .B1(_08210_),
    .X(_08319_));
 sky130_fd_sc_hd__a21o_1 _15225_ (.A1(_08316_),
    .A2(_08319_),
    .B1(_08239_),
    .X(_08320_));
 sky130_fd_sc_hd__buf_4 _15226_ (.A(_08309_),
    .X(_08321_));
 sky130_fd_sc_hd__nand2_1 _15227_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__or4_1 _15228_ (.A(_08084_),
    .B(_08090_),
    .C(_08097_),
    .D(_08217_),
    .X(_08323_));
 sky130_fd_sc_hd__clkbuf_2 _15229_ (.A(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__o31ai_1 _15230_ (.A1(_08084_),
    .A2(_08090_),
    .A3(_08217_),
    .B1(_08097_),
    .Y(_08325_));
 sky130_fd_sc_hd__mux2_2 _15231_ (.A0(_06091_),
    .A1(_06403_),
    .S(_04535_),
    .X(_08326_));
 sky130_fd_sc_hd__a21o_1 _15232_ (.A1(_08210_),
    .A2(_08326_),
    .B1(_08216_),
    .X(_08327_));
 sky130_fd_sc_hd__a31o_1 _15233_ (.A1(_08214_),
    .A2(_08324_),
    .A3(_08325_),
    .B1(_08327_),
    .X(_08328_));
 sky130_fd_sc_hd__nand2_1 _15234_ (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .B(_08239_),
    .Y(_08329_));
 sky130_fd_sc_hd__a21o_2 _15235_ (.A1(_08328_),
    .A2(_08329_),
    .B1(_08231_),
    .X(_08330_));
 sky130_fd_sc_hd__nor4_1 _15236_ (.A(_08314_),
    .B(_08320_),
    .C(_08322_),
    .D(_08330_),
    .Y(_08331_));
 sky130_fd_sc_hd__o22ai_1 _15237_ (.A1(_08314_),
    .A2(_08320_),
    .B1(_08322_),
    .B2(_08330_),
    .Y(_08332_));
 sky130_fd_sc_hd__and2b_1 _15238_ (.A_N(_08331_),
    .B(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__xor2_2 _15239_ (.A(_08313_),
    .B(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__or2_1 _15240_ (.A(_08239_),
    .B(_08303_),
    .X(_08335_));
 sky130_fd_sc_hd__clkbuf_4 _15241_ (.A(_08320_),
    .X(_08336_));
 sky130_fd_sc_hd__or4_1 _15242_ (.A(_08314_),
    .B(_08335_),
    .C(_08336_),
    .D(_08322_),
    .X(_08337_));
 sky130_fd_sc_hd__nor2_1 _15243_ (.A(_08233_),
    .B(_08312_),
    .Y(_08338_));
 sky130_fd_sc_hd__nor2_2 _15244_ (.A(_08298_),
    .B(_08303_),
    .Y(_08339_));
 sky130_fd_sc_hd__a21oi_2 _15245_ (.A1(_08316_),
    .A2(_08319_),
    .B1(_08298_),
    .Y(_08340_));
 sky130_fd_sc_hd__inv_2 _15246_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .Y(_08341_));
 sky130_fd_sc_hd__nor2_1 _15247_ (.A(_08341_),
    .B(_08215_),
    .Y(_08342_));
 sky130_fd_sc_hd__a22o_1 _15248_ (.A1(_08131_),
    .A2(_08339_),
    .B1(_08340_),
    .B2(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__nand3_1 _15249_ (.A(_08337_),
    .B(_08338_),
    .C(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__nand2_1 _15250_ (.A(_08337_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__xor2_2 _15251_ (.A(_08334_),
    .B(_08345_),
    .X(_08346_));
 sky130_fd_sc_hd__xnor2_2 _15252_ (.A(_08297_),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__a21o_1 _15253_ (.A1(_08337_),
    .A2(_08343_),
    .B1(_08338_),
    .X(_08348_));
 sky130_fd_sc_hd__nor2_2 _15254_ (.A(_08341_),
    .B(_08223_),
    .Y(_08349_));
 sky130_fd_sc_hd__a221o_4 _15255_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08234_),
    .B1(_08231_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08310_),
    .X(_08350_));
 sky130_fd_sc_hd__nand2_2 _15256_ (.A(_08131_),
    .B(_08234_),
    .Y(_08351_));
 sky130_fd_sc_hd__or4bb_1 _15257_ (.A(_08351_),
    .B(_08302_),
    .C_N(_08228_),
    .D_N(_08349_),
    .X(_08352_));
 sky130_fd_sc_hd__nand2_1 _15258_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08234_),
    .Y(_08353_));
 sky130_fd_sc_hd__buf_2 _15259_ (.A(_08353_),
    .X(_08354_));
 sky130_fd_sc_hd__nor2_2 _15260_ (.A(_08314_),
    .B(_08239_),
    .Y(_08355_));
 sky130_fd_sc_hd__a2bb2o_1 _15261_ (.A1_N(_08303_),
    .A2_N(_08354_),
    .B1(_08355_),
    .B2(_08228_),
    .X(_08356_));
 sky130_fd_sc_hd__and4b_1 _15262_ (.A_N(_08243_),
    .B(_08350_),
    .C(_08352_),
    .D(_08356_),
    .X(_08357_));
 sky130_fd_sc_hd__a41o_1 _15263_ (.A1(_08131_),
    .A2(_08228_),
    .A3(_08339_),
    .A4(_08349_),
    .B1(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__a21o_1 _15264_ (.A1(_08344_),
    .A2(_08348_),
    .B1(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__or4_1 _15265_ (.A(_08272_),
    .B(_08268_),
    .C(_08243_),
    .D(_08295_),
    .X(_08360_));
 sky130_fd_sc_hd__inv_2 _15266_ (.A(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__clkbuf_4 _15267_ (.A(_08272_),
    .X(_08362_));
 sky130_fd_sc_hd__o22a_1 _15268_ (.A1(_08271_),
    .A2(_08244_),
    .B1(_08295_),
    .B2(_08362_),
    .X(_08363_));
 sky130_fd_sc_hd__nor2_1 _15269_ (.A(_08361_),
    .B(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__nor2_1 _15270_ (.A(\rbzero.side_hot ),
    .B(_06112_),
    .Y(_08365_));
 sky130_fd_sc_hd__a211o_1 _15271_ (.A1(\rbzero.side_hot ),
    .A2(_06431_),
    .B1(_08213_),
    .C1(_08365_),
    .X(_08366_));
 sky130_fd_sc_hd__o211ai_4 _15272_ (.A1(_08057_),
    .A2(_08209_),
    .B1(_08366_),
    .C1(_06336_),
    .Y(_08367_));
 sky130_fd_sc_hd__o21ai_1 _15273_ (.A1(\rbzero.wall_tracer.stepDistY[-3] ),
    .A2(_08225_),
    .B1(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__o21bai_2 _15274_ (.A1(\rbzero.wall_tracer.stepDistX[-3] ),
    .A2(_06339_),
    .B1_N(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__clkbuf_4 _15275_ (.A(_08369_),
    .X(_08370_));
 sky130_fd_sc_hd__clkbuf_4 _15276_ (.A(_08288_),
    .X(_08371_));
 sky130_fd_sc_hd__nor2_1 _15277_ (.A(_08370_),
    .B(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__xor2_2 _15278_ (.A(_08364_),
    .B(_08372_),
    .X(_08373_));
 sky130_fd_sc_hd__nand3_1 _15279_ (.A(_08344_),
    .B(_08348_),
    .C(_08358_),
    .Y(_08374_));
 sky130_fd_sc_hd__a21boi_2 _15280_ (.A1(_08359_),
    .A2(_08373_),
    .B1_N(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__xor2_1 _15281_ (.A(_08347_),
    .B(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__nand2_1 _15282_ (.A(\rbzero.side_hot ),
    .B(_06436_),
    .Y(_08377_));
 sky130_fd_sc_hd__o211a_1 _15283_ (.A1(_04535_),
    .A2(_06115_),
    .B1(_08208_),
    .C1(_08377_),
    .X(_08378_));
 sky130_fd_sc_hd__a211o_2 _15284_ (.A1(_08049_),
    .A2(_08213_),
    .B1(_08378_),
    .C1(_08223_),
    .X(_08379_));
 sky130_fd_sc_hd__o221ai_4 _15285_ (.A1(\rbzero.wall_tracer.stepDistX[-4] ),
    .A2(_06338_),
    .B1(_08309_),
    .B2(\rbzero.wall_tracer.stepDistY[-4] ),
    .C1(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__nor2_1 _15286_ (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(_06338_),
    .Y(_08381_));
 sky130_fd_sc_hd__nor2_1 _15287_ (.A(\rbzero.side_hot ),
    .B(_06117_),
    .Y(_08382_));
 sky130_fd_sc_hd__a211o_1 _15288_ (.A1(\rbzero.side_hot ),
    .A2(_06440_),
    .B1(_08213_),
    .C1(_08382_),
    .X(_08383_));
 sky130_fd_sc_hd__o21a_1 _15289_ (.A1(_08040_),
    .A2(_08208_),
    .B1(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__a2bb2o_2 _15290_ (.A1_N(\rbzero.wall_tracer.stepDistY[-5] ),
    .A2_N(_08225_),
    .B1(_08384_),
    .B2(_06336_),
    .X(_08385_));
 sky130_fd_sc_hd__or2_1 _15291_ (.A(_08381_),
    .B(_08385_),
    .X(_08386_));
 sky130_fd_sc_hd__buf_2 _15292_ (.A(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__inv_2 _15293_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .Y(_08388_));
 sky130_fd_sc_hd__xnor2_1 _15294_ (.A(_08388_),
    .B(_08281_),
    .Y(_08389_));
 sky130_fd_sc_hd__mux2_1 _15295_ (.A0(_08389_),
    .A1(\rbzero.debug_overlay.playerX[-5] ),
    .S(_08285_),
    .X(_08390_));
 sky130_fd_sc_hd__xnor2_1 _15296_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_08276_),
    .Y(_08391_));
 sky130_fd_sc_hd__nand2_1 _15297_ (.A(_06135_),
    .B(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__o211a_1 _15298_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_06135_),
    .B1(_08215_),
    .C1(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__a211o_1 _15299_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_08225_),
    .B1(_08393_),
    .C1(_08230_),
    .X(_08394_));
 sky130_fd_sc_hd__o21ai_4 _15300_ (.A1(_06339_),
    .A2(_08390_),
    .B1(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__buf_2 _15301_ (.A(_08395_),
    .X(_08396_));
 sky130_fd_sc_hd__or3_1 _15302_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .C(_08276_),
    .X(_08397_));
 sky130_fd_sc_hd__o21ai_1 _15303_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_08276_),
    .B1(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_08398_));
 sky130_fd_sc_hd__nand2_1 _15304_ (.A(_08397_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__nor2_1 _15305_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(_06136_),
    .Y(_08400_));
 sky130_fd_sc_hd__a211o_1 _15306_ (.A1(_06136_),
    .A2(_08399_),
    .B1(_08400_),
    .C1(_08225_),
    .X(_08401_));
 sky130_fd_sc_hd__a21oi_1 _15307_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_06336_),
    .B1(_08230_),
    .Y(_08402_));
 sky130_fd_sc_hd__or3_1 _15308_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(\rbzero.debug_overlay.playerX[-5] ),
    .C(_08281_),
    .X(_08403_));
 sky130_fd_sc_hd__o21ai_1 _15309_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_08281_),
    .B1(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_08404_));
 sky130_fd_sc_hd__nand2_1 _15310_ (.A(_08403_),
    .B(_08404_),
    .Y(_08405_));
 sky130_fd_sc_hd__inv_2 _15311_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_08406_));
 sky130_fd_sc_hd__mux2_1 _15312_ (.A0(_08405_),
    .A1(_08406_),
    .S(_08252_),
    .X(_08407_));
 sky130_fd_sc_hd__a22o_4 _15313_ (.A1(_08401_),
    .A2(_08402_),
    .B1(_08407_),
    .B2(_08230_),
    .X(_08408_));
 sky130_fd_sc_hd__clkbuf_4 _15314_ (.A(_08408_),
    .X(_08409_));
 sky130_fd_sc_hd__or4_1 _15315_ (.A(_08380_),
    .B(_08387_),
    .C(_08396_),
    .D(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__nor2_1 _15316_ (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .B(_06339_),
    .Y(_08411_));
 sky130_fd_sc_hd__a31o_1 _15317_ (.A1(_08020_),
    .A2(_08026_),
    .A3(_08029_),
    .B1(_08209_),
    .X(_08412_));
 sky130_fd_sc_hd__mux2_1 _15318_ (.A0(_06121_),
    .A1(_06470_),
    .S(\rbzero.side_hot ),
    .X(_08413_));
 sky130_fd_sc_hd__a21oi_1 _15319_ (.A1(_08209_),
    .A2(_08413_),
    .B1(_08223_),
    .Y(_08414_));
 sky130_fd_sc_hd__a2bb2o_2 _15320_ (.A1_N(\rbzero.wall_tracer.stepDistY[-6] ),
    .A2_N(_08225_),
    .B1(_08412_),
    .B2(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__or2_1 _15321_ (.A(_08411_),
    .B(_08415_),
    .X(_08416_));
 sky130_fd_sc_hd__clkbuf_2 _15322_ (.A(_08416_),
    .X(_08417_));
 sky130_fd_sc_hd__or2_1 _15323_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08403_),
    .X(_08418_));
 sky130_fd_sc_hd__nand2_1 _15324_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08403_),
    .Y(_08419_));
 sky130_fd_sc_hd__and2_1 _15325_ (.A(_08418_),
    .B(_08419_),
    .X(_08420_));
 sky130_fd_sc_hd__mux2_1 _15326_ (.A0(_08420_),
    .A1(\rbzero.debug_overlay.playerX[-3] ),
    .S(_08285_),
    .X(_08421_));
 sky130_fd_sc_hd__or2_1 _15327_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08397_),
    .X(_08422_));
 sky130_fd_sc_hd__nand2_1 _15328_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08397_),
    .Y(_08423_));
 sky130_fd_sc_hd__nand2_1 _15329_ (.A(_08422_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__nand2_1 _15330_ (.A(_06136_),
    .B(_08424_),
    .Y(_08425_));
 sky130_fd_sc_hd__o211a_1 _15331_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_06136_),
    .B1(_08216_),
    .C1(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__a211o_1 _15332_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_08309_),
    .B1(_08426_),
    .C1(_08230_),
    .X(_08427_));
 sky130_fd_sc_hd__o21ai_4 _15333_ (.A1(_06339_),
    .A2(_08421_),
    .B1(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__clkbuf_4 _15334_ (.A(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__buf_2 _15335_ (.A(_08380_),
    .X(_08430_));
 sky130_fd_sc_hd__o22ai_1 _15336_ (.A1(_08430_),
    .A2(_08396_),
    .B1(_08409_),
    .B2(_08387_),
    .Y(_08431_));
 sky130_fd_sc_hd__nand2_1 _15337_ (.A(_08410_),
    .B(_08431_),
    .Y(_08432_));
 sky130_fd_sc_hd__or3_1 _15338_ (.A(_08417_),
    .B(_08429_),
    .C(_08432_),
    .X(_08433_));
 sky130_fd_sc_hd__nand2_1 _15339_ (.A(_08410_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__a21oi_2 _15340_ (.A1(_08364_),
    .A2(_08372_),
    .B1(_08361_),
    .Y(_08435_));
 sky130_fd_sc_hd__or2_1 _15341_ (.A(_08370_),
    .B(_08409_),
    .X(_08436_));
 sky130_fd_sc_hd__or3_1 _15342_ (.A(_08430_),
    .B(_08396_),
    .C(_08436_),
    .X(_08437_));
 sky130_fd_sc_hd__clkbuf_4 _15343_ (.A(_08396_),
    .X(_08438_));
 sky130_fd_sc_hd__o22ai_1 _15344_ (.A1(_08370_),
    .A2(_08438_),
    .B1(_08409_),
    .B2(_08430_),
    .Y(_08439_));
 sky130_fd_sc_hd__nand2_1 _15345_ (.A(_08437_),
    .B(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__or3_1 _15346_ (.A(_08387_),
    .B(_08429_),
    .C(_08440_),
    .X(_08441_));
 sky130_fd_sc_hd__clkbuf_4 _15347_ (.A(_08429_),
    .X(_08442_));
 sky130_fd_sc_hd__o21ai_1 _15348_ (.A1(_08387_),
    .A2(_08442_),
    .B1(_08440_),
    .Y(_08443_));
 sky130_fd_sc_hd__nand2_1 _15349_ (.A(_08441_),
    .B(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__xnor2_1 _15350_ (.A(_08435_),
    .B(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__xnor2_1 _15351_ (.A(_08434_),
    .B(_08445_),
    .Y(_08446_));
 sky130_fd_sc_hd__xnor2_1 _15352_ (.A(_08376_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__nand2_1 _15353_ (.A(_08374_),
    .B(_08359_),
    .Y(_08448_));
 sky130_fd_sc_hd__xor2_2 _15354_ (.A(_08448_),
    .B(_08373_),
    .X(_08449_));
 sky130_fd_sc_hd__a2bb2oi_1 _15355_ (.A1_N(_08244_),
    .A2_N(_08312_),
    .B1(_08352_),
    .B2(_08356_),
    .Y(_08450_));
 sky130_fd_sc_hd__nand2_1 _15356_ (.A(_08227_),
    .B(_08349_),
    .Y(_08451_));
 sky130_fd_sc_hd__nand2_1 _15357_ (.A(_08238_),
    .B(_08355_),
    .Y(_08452_));
 sky130_fd_sc_hd__xnor2_2 _15358_ (.A(_08451_),
    .B(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__or2_1 _15359_ (.A(_08294_),
    .B(_08311_),
    .X(_08454_));
 sky130_fd_sc_hd__nor2_1 _15360_ (.A(_08451_),
    .B(_08452_),
    .Y(_08455_));
 sky130_fd_sc_hd__o21ba_1 _15361_ (.A1(_08453_),
    .A2(_08454_),
    .B1_N(_08455_),
    .X(_08456_));
 sky130_fd_sc_hd__nor2_1 _15362_ (.A(_08357_),
    .B(_08450_),
    .Y(_08457_));
 sky130_fd_sc_hd__xnor2_2 _15363_ (.A(_08457_),
    .B(_08456_),
    .Y(_08458_));
 sky130_fd_sc_hd__or4_1 _15364_ (.A(_08369_),
    .B(_08259_),
    .C(_08268_),
    .D(_08294_),
    .X(_08459_));
 sky130_fd_sc_hd__o22ai_1 _15365_ (.A1(_08370_),
    .A2(_08272_),
    .B1(_08268_),
    .B2(_08295_),
    .Y(_08460_));
 sky130_fd_sc_hd__nand2_1 _15366_ (.A(_08459_),
    .B(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__or3_1 _15367_ (.A(_08380_),
    .B(_08288_),
    .C(_08461_),
    .X(_08462_));
 sky130_fd_sc_hd__o21ai_1 _15368_ (.A1(_08430_),
    .A2(_08288_),
    .B1(_08461_),
    .Y(_08463_));
 sky130_fd_sc_hd__and2_1 _15369_ (.A(_08462_),
    .B(_08463_),
    .X(_08464_));
 sky130_fd_sc_hd__nand2_1 _15370_ (.A(_08458_),
    .B(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__o31a_1 _15371_ (.A1(_08357_),
    .A2(_08450_),
    .A3(_08456_),
    .B1(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__xor2_1 _15372_ (.A(_08449_),
    .B(_08466_),
    .X(_08467_));
 sky130_fd_sc_hd__nor2_2 _15373_ (.A(_08411_),
    .B(_08415_),
    .Y(_08468_));
 sky130_fd_sc_hd__clkinv_2 _15374_ (.A(_08408_),
    .Y(_08469_));
 sky130_fd_sc_hd__a2bb2o_1 _15375_ (.A1_N(_08386_),
    .A2_N(_08396_),
    .B1(_08468_),
    .B2(_08469_),
    .X(_08470_));
 sky130_fd_sc_hd__nor2_1 _15376_ (.A(\rbzero.wall_tracer.stepDistX[-7] ),
    .B(_06338_),
    .Y(_08471_));
 sky130_fd_sc_hd__a21o_1 _15377_ (.A1(_08011_),
    .A2(_08016_),
    .B1(_08209_),
    .X(_08472_));
 sky130_fd_sc_hd__nand2_1 _15378_ (.A(_04535_),
    .B(_06449_),
    .Y(_08473_));
 sky130_fd_sc_hd__o211a_1 _15379_ (.A1(_04535_),
    .A2(_06123_),
    .B1(_08208_),
    .C1(_08473_),
    .X(_08474_));
 sky130_fd_sc_hd__nor2_1 _15380_ (.A(_08223_),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__a2bb2o_4 _15381_ (.A1_N(\rbzero.wall_tracer.stepDistY[-7] ),
    .A2_N(_08225_),
    .B1(_08472_),
    .B2(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__or2_1 _15382_ (.A(_08471_),
    .B(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__clkbuf_4 _15383_ (.A(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__nor2_1 _15384_ (.A(_08478_),
    .B(_08429_),
    .Y(_08479_));
 sky130_fd_sc_hd__or4_1 _15385_ (.A(_08386_),
    .B(_08396_),
    .C(_08417_),
    .D(_08408_),
    .X(_08480_));
 sky130_fd_sc_hd__a21bo_1 _15386_ (.A1(_08470_),
    .A2(_08479_),
    .B1_N(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__o21ai_1 _15387_ (.A1(_08417_),
    .A2(_08442_),
    .B1(_08432_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand2_1 _15388_ (.A(_08433_),
    .B(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__a21o_1 _15389_ (.A1(_08459_),
    .A2(_08462_),
    .B1(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__nand3_1 _15390_ (.A(_08459_),
    .B(_08462_),
    .C(_08483_),
    .Y(_08485_));
 sky130_fd_sc_hd__nand2_1 _15391_ (.A(_08484_),
    .B(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__xnor2_1 _15392_ (.A(_08481_),
    .B(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__nor2_1 _15393_ (.A(_08449_),
    .B(_08466_),
    .Y(_08488_));
 sky130_fd_sc_hd__a21oi_1 _15394_ (.A1(_08467_),
    .A2(_08487_),
    .B1(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__nor2_1 _15395_ (.A(_08447_),
    .B(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__and2_1 _15396_ (.A(_08447_),
    .B(_08489_),
    .X(_08491_));
 sky130_fd_sc_hd__nor2_1 _15397_ (.A(_08490_),
    .B(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__buf_4 _15398_ (.A(_08234_),
    .X(_08493_));
 sky130_fd_sc_hd__nand2_4 _15399_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__buf_4 _15400_ (.A(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__buf_6 _15401_ (.A(_08493_),
    .X(_08496_));
 sky130_fd_sc_hd__mux2_1 _15402_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(_04535_),
    .X(_08497_));
 sky130_fd_sc_hd__a21o_1 _15403_ (.A1(_08210_),
    .A2(_08497_),
    .B1(_08216_),
    .X(_08498_));
 sky130_fd_sc_hd__a21o_2 _15404_ (.A1(_07951_),
    .A2(_08214_),
    .B1(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__o211ai_4 _15405_ (.A1(\rbzero.wall_tracer.stepDistY[-11] ),
    .A2(_08496_),
    .B1(_06340_),
    .C1(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__nor2_2 _15406_ (.A(_08495_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__mux2_1 _15407_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(\rbzero.side_hot ),
    .X(_08502_));
 sky130_fd_sc_hd__or2_1 _15408_ (.A(_08213_),
    .B(_08502_),
    .X(_08503_));
 sky130_fd_sc_hd__o211a_2 _15409_ (.A1(_07977_),
    .A2(_08209_),
    .B1(_08503_),
    .C1(_08309_),
    .X(_08504_));
 sky130_fd_sc_hd__a211oi_4 _15410_ (.A1(\rbzero.wall_tracer.stepDistY[-10] ),
    .A2(_08239_),
    .B1(_08230_),
    .C1(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__nand2_4 _15411_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08234_),
    .Y(_08506_));
 sky130_fd_sc_hd__nor2_2 _15412_ (.A(_08505_),
    .B(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__nand2_2 _15413_ (.A(_08501_),
    .B(_08507_),
    .Y(_08508_));
 sky130_fd_sc_hd__clkbuf_4 _15414_ (.A(_08505_),
    .X(_08509_));
 sky130_fd_sc_hd__clkbuf_4 _15415_ (.A(_08506_),
    .X(_08510_));
 sky130_fd_sc_hd__clkbuf_4 _15416_ (.A(_08500_),
    .X(_08511_));
 sky130_fd_sc_hd__o22ai_4 _15417_ (.A1(_08495_),
    .A2(_08509_),
    .B1(_08510_),
    .B2(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__or3_2 _15418_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .B(\rbzero.debug_overlay.playerX[-2] ),
    .C(_08418_),
    .X(_08513_));
 sky130_fd_sc_hd__or3_2 _15419_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .C(_08422_),
    .X(_08514_));
 sky130_fd_sc_hd__inv_2 _15420_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .Y(_08515_));
 sky130_fd_sc_hd__o32a_1 _15421_ (.A1(_06146_),
    .A2(_08309_),
    .A3(_08514_),
    .B1(_08239_),
    .B2(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__o31a_4 _15422_ (.A1(_06339_),
    .A2(_08285_),
    .A3(_08513_),
    .B1(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__mux2_1 _15423_ (.A0(_06126_),
    .A1(_06463_),
    .S(_04535_),
    .X(_08518_));
 sky130_fd_sc_hd__mux2_1 _15424_ (.A0(_07988_),
    .A1(_08518_),
    .S(_08209_),
    .X(_08519_));
 sky130_fd_sc_hd__o22ai_4 _15425_ (.A1(\rbzero.wall_tracer.stepDistY[-9] ),
    .A2(_08309_),
    .B1(_08519_),
    .B2(_08223_),
    .Y(_08520_));
 sky130_fd_sc_hd__o21bai_4 _15426_ (.A1(\rbzero.wall_tracer.stepDistX[-9] ),
    .A2(_06339_),
    .B1_N(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__buf_2 _15427_ (.A(_08521_),
    .X(_08522_));
 sky130_fd_sc_hd__nor2_2 _15428_ (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .B(_06338_),
    .Y(_08523_));
 sky130_fd_sc_hd__a21o_1 _15429_ (.A1(_08001_),
    .A2(_08004_),
    .B1(_08209_),
    .X(_08524_));
 sky130_fd_sc_hd__mux2_1 _15430_ (.A0(_06125_),
    .A1(_06454_),
    .S(\rbzero.side_hot ),
    .X(_08525_));
 sky130_fd_sc_hd__a21oi_1 _15431_ (.A1(_08209_),
    .A2(_08525_),
    .B1(_08223_),
    .Y(_08526_));
 sky130_fd_sc_hd__a2bb2o_2 _15432_ (.A1_N(\rbzero.wall_tracer.stepDistY[-8] ),
    .A2_N(_08225_),
    .B1(_08524_),
    .B2(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__or2_1 _15433_ (.A(_08523_),
    .B(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__clkbuf_4 _15434_ (.A(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__xor2_1 _15435_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_08418_),
    .X(_08530_));
 sky130_fd_sc_hd__mux2_1 _15436_ (.A0(_08530_),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_08285_),
    .X(_08531_));
 sky130_fd_sc_hd__xnor2_1 _15437_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_08422_),
    .Y(_08532_));
 sky130_fd_sc_hd__nand2_1 _15438_ (.A(_06136_),
    .B(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__o211a_1 _15439_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_06136_),
    .B1(_08216_),
    .C1(_08533_),
    .X(_08534_));
 sky130_fd_sc_hd__a211o_1 _15440_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_08309_),
    .B1(_08534_),
    .C1(_08231_),
    .X(_08535_));
 sky130_fd_sc_hd__o21ai_4 _15441_ (.A1(_06339_),
    .A2(_08531_),
    .B1(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__or2_1 _15442_ (.A(_08529_),
    .B(_08536_),
    .X(_08537_));
 sky130_fd_sc_hd__o21ai_1 _15443_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_08418_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_08538_));
 sky130_fd_sc_hd__and2_1 _15444_ (.A(_08513_),
    .B(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__mux2_1 _15445_ (.A0(_08539_),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_08285_),
    .X(_08540_));
 sky130_fd_sc_hd__o21ai_1 _15446_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_08422_),
    .B1(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_08541_));
 sky130_fd_sc_hd__and2_1 _15447_ (.A(_08514_),
    .B(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__mux2_1 _15448_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(_08542_),
    .S(_06136_),
    .X(_08543_));
 sky130_fd_sc_hd__or2_1 _15449_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(_08223_),
    .X(_08544_));
 sky130_fd_sc_hd__mux2_1 _15450_ (.A0(_08543_),
    .A1(_08544_),
    .S(_08309_),
    .X(_08545_));
 sky130_fd_sc_hd__o21ai_4 _15451_ (.A1(_06339_),
    .A2(_08540_),
    .B1(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__clkbuf_4 _15452_ (.A(_08536_),
    .X(_08547_));
 sky130_fd_sc_hd__o22ai_1 _15453_ (.A1(_08478_),
    .A2(_08547_),
    .B1(_08546_),
    .B2(_08529_),
    .Y(_08548_));
 sky130_fd_sc_hd__o31a_1 _15454_ (.A1(_08478_),
    .A2(_08537_),
    .A3(_08546_),
    .B1(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__or3b_1 _15455_ (.A(_08517_),
    .B(_08522_),
    .C_N(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__clkbuf_4 _15456_ (.A(_08517_),
    .X(_08551_));
 sky130_fd_sc_hd__o21bai_1 _15457_ (.A1(_08522_),
    .A2(_08551_),
    .B1_N(_08549_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_1 _15458_ (.A(_08550_),
    .B(_08552_),
    .Y(_08553_));
 sky130_fd_sc_hd__inv_2 _15459_ (.A(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_08554_));
 sky130_fd_sc_hd__a21o_4 _15460_ (.A1(_08554_),
    .A2(_08231_),
    .B1(_08505_),
    .X(_08555_));
 sky130_fd_sc_hd__nor2_1 _15461_ (.A(_08517_),
    .B(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__nor2_1 _15462_ (.A(_08546_),
    .B(_08522_),
    .Y(_08557_));
 sky130_fd_sc_hd__xnor2_1 _15463_ (.A(_08537_),
    .B(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__buf_4 _15464_ (.A(_08546_),
    .X(_08559_));
 sky130_fd_sc_hd__or3_1 _15465_ (.A(_08537_),
    .B(_08559_),
    .C(_08522_),
    .X(_08560_));
 sky130_fd_sc_hd__a21boi_1 _15466_ (.A1(_08556_),
    .A2(_08558_),
    .B1_N(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__nor2_1 _15467_ (.A(_08553_),
    .B(_08561_),
    .Y(_08562_));
 sky130_fd_sc_hd__and2_1 _15468_ (.A(_08553_),
    .B(_08561_),
    .X(_08563_));
 sky130_fd_sc_hd__nor2_1 _15469_ (.A(_08562_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__a31o_1 _15470_ (.A1(_08508_),
    .A2(_08512_),
    .A3(_08564_),
    .B1(_08562_),
    .X(_08565_));
 sky130_fd_sc_hd__or2b_1 _15471_ (.A(_08486_),
    .B_N(_08481_),
    .X(_08566_));
 sky130_fd_sc_hd__clkbuf_4 _15472_ (.A(_08520_),
    .X(_08567_));
 sky130_fd_sc_hd__nor2_1 _15473_ (.A(_08494_),
    .B(_08567_),
    .Y(_08568_));
 sky130_fd_sc_hd__or2_1 _15474_ (.A(_08507_),
    .B(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__nand2_1 _15475_ (.A(_08507_),
    .B(_08568_),
    .Y(_08570_));
 sky130_fd_sc_hd__nand2_1 _15476_ (.A(_08569_),
    .B(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__nand2_1 _15477_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08493_),
    .Y(_08572_));
 sky130_fd_sc_hd__buf_2 _15478_ (.A(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__nor2_1 _15479_ (.A(_08511_),
    .B(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__xnor2_1 _15480_ (.A(_08571_),
    .B(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__or2_1 _15481_ (.A(_08478_),
    .B(_08536_),
    .X(_08576_));
 sky130_fd_sc_hd__or2_1 _15482_ (.A(_08417_),
    .B(_08546_),
    .X(_08577_));
 sky130_fd_sc_hd__or2_1 _15483_ (.A(_08576_),
    .B(_08577_),
    .X(_08578_));
 sky130_fd_sc_hd__o22ai_1 _15484_ (.A1(_08417_),
    .A2(_08547_),
    .B1(_08546_),
    .B2(_08478_),
    .Y(_08579_));
 sky130_fd_sc_hd__nand2_1 _15485_ (.A(_08578_),
    .B(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__nor2_1 _15486_ (.A(_08529_),
    .B(_08517_),
    .Y(_08581_));
 sky130_fd_sc_hd__xnor2_1 _15487_ (.A(_08580_),
    .B(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__buf_4 _15488_ (.A(_08559_),
    .X(_08583_));
 sky130_fd_sc_hd__o31a_1 _15489_ (.A1(_08529_),
    .A2(_08583_),
    .A3(_08576_),
    .B1(_08550_),
    .X(_08584_));
 sky130_fd_sc_hd__xnor2_1 _15490_ (.A(_08582_),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__nand2_1 _15491_ (.A(_08575_),
    .B(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__or2_1 _15492_ (.A(_08575_),
    .B(_08585_),
    .X(_08587_));
 sky130_fd_sc_hd__nand2_1 _15493_ (.A(_08586_),
    .B(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__a21o_1 _15494_ (.A1(_08484_),
    .A2(_08566_),
    .B1(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__nand3_1 _15495_ (.A(_08484_),
    .B(_08566_),
    .C(_08588_),
    .Y(_08590_));
 sky130_fd_sc_hd__nand2_1 _15496_ (.A(_08589_),
    .B(_08590_),
    .Y(_08591_));
 sky130_fd_sc_hd__xnor2_1 _15497_ (.A(_08565_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__xnor2_1 _15498_ (.A(_08492_),
    .B(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__xnor2_1 _15499_ (.A(_08467_),
    .B(_08487_),
    .Y(_08594_));
 sky130_fd_sc_hd__xnor2_2 _15500_ (.A(_08458_),
    .B(_08464_),
    .Y(_08595_));
 sky130_fd_sc_hd__xnor2_2 _15501_ (.A(_08453_),
    .B(_08454_),
    .Y(_08596_));
 sky130_fd_sc_hd__nand2_1 _15502_ (.A(_08292_),
    .B(_08342_),
    .Y(_08597_));
 sky130_fd_sc_hd__or3b_1 _15503_ (.A(_08351_),
    .B(_08597_),
    .C_N(_08238_),
    .X(_08598_));
 sky130_fd_sc_hd__nor2_1 _15504_ (.A(_08314_),
    .B(_08216_),
    .Y(_08599_));
 sky130_fd_sc_hd__a22o_1 _15505_ (.A1(_08238_),
    .A2(_08349_),
    .B1(_08599_),
    .B2(_08292_),
    .X(_08600_));
 sky130_fd_sc_hd__or4bb_1 _15506_ (.A(_08369_),
    .B(_08311_),
    .C_N(_08598_),
    .D_N(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__and2_1 _15507_ (.A(_08598_),
    .B(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__xor2_2 _15508_ (.A(_08596_),
    .B(_08602_),
    .X(_08603_));
 sky130_fd_sc_hd__or4_1 _15509_ (.A(_08369_),
    .B(_08259_),
    .C(_08268_),
    .D(_08380_),
    .X(_08604_));
 sky130_fd_sc_hd__o22ai_1 _15510_ (.A1(_08369_),
    .A2(_08268_),
    .B1(_08380_),
    .B2(_08259_),
    .Y(_08605_));
 sky130_fd_sc_hd__nand2_1 _15511_ (.A(_08604_),
    .B(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__or3_1 _15512_ (.A(_08606_),
    .B(_08287_),
    .C(_08386_),
    .X(_08607_));
 sky130_fd_sc_hd__o21ai_1 _15513_ (.A1(_08287_),
    .A2(_08387_),
    .B1(_08606_),
    .Y(_08608_));
 sky130_fd_sc_hd__and2_1 _15514_ (.A(_08607_),
    .B(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__nor2_1 _15515_ (.A(_08596_),
    .B(_08602_),
    .Y(_08610_));
 sky130_fd_sc_hd__a21o_1 _15516_ (.A1(_08603_),
    .A2(_08609_),
    .B1(_08610_),
    .X(_08611_));
 sky130_fd_sc_hd__xnor2_1 _15517_ (.A(_08595_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__nor2_1 _15518_ (.A(_08395_),
    .B(_08417_),
    .Y(_08613_));
 sky130_fd_sc_hd__nor2_1 _15519_ (.A(_08408_),
    .B(_08478_),
    .Y(_08614_));
 sky130_fd_sc_hd__xor2_1 _15520_ (.A(_08613_),
    .B(_08614_),
    .X(_08615_));
 sky130_fd_sc_hd__nor2_1 _15521_ (.A(_08428_),
    .B(_08529_),
    .Y(_08616_));
 sky130_fd_sc_hd__a22o_1 _15522_ (.A1(_08613_),
    .A2(_08614_),
    .B1(_08615_),
    .B2(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__nand2_1 _15523_ (.A(_08480_),
    .B(_08470_),
    .Y(_08618_));
 sky130_fd_sc_hd__xor2_1 _15524_ (.A(_08618_),
    .B(_08479_),
    .X(_08619_));
 sky130_fd_sc_hd__a21o_1 _15525_ (.A1(_08604_),
    .A2(_08607_),
    .B1(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__nand3_1 _15526_ (.A(_08604_),
    .B(_08607_),
    .C(_08619_),
    .Y(_08621_));
 sky130_fd_sc_hd__and2_1 _15527_ (.A(_08620_),
    .B(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__xor2_1 _15528_ (.A(_08617_),
    .B(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__and2b_1 _15529_ (.A_N(_08595_),
    .B(_08611_),
    .X(_08624_));
 sky130_fd_sc_hd__a21oi_1 _15530_ (.A1(_08612_),
    .A2(_08623_),
    .B1(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__nand2_1 _15531_ (.A(_08594_),
    .B(_08625_),
    .Y(_08626_));
 sky130_fd_sc_hd__xnor2_1 _15532_ (.A(_08556_),
    .B(_08558_),
    .Y(_08627_));
 sky130_fd_sc_hd__nor2_1 _15533_ (.A(_08547_),
    .B(_08555_),
    .Y(_08628_));
 sky130_fd_sc_hd__buf_4 _15534_ (.A(_08231_),
    .X(_08629_));
 sky130_fd_sc_hd__o211a_2 _15535_ (.A1(\rbzero.wall_tracer.stepDistY[-11] ),
    .A2(_08234_),
    .B1(_06339_),
    .C1(_08499_),
    .X(_08630_));
 sky130_fd_sc_hd__a21oi_2 _15536_ (.A1(\rbzero.wall_tracer.stepDistX[-11] ),
    .A2(_08629_),
    .B1(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__or2_1 _15537_ (.A(_08517_),
    .B(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__o22a_1 _15538_ (.A1(_08547_),
    .A2(_08522_),
    .B1(_08555_),
    .B2(_08546_),
    .X(_08633_));
 sky130_fd_sc_hd__o2bb2a_1 _15539_ (.A1_N(_08557_),
    .A2_N(_08628_),
    .B1(_08632_),
    .B2(_08633_),
    .X(_08634_));
 sky130_fd_sc_hd__xor2_1 _15540_ (.A(_08627_),
    .B(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__nand2_2 _15541_ (.A(_08501_),
    .B(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__o21ai_2 _15542_ (.A1(_08627_),
    .A2(_08634_),
    .B1(_08636_),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_1 _15543_ (.A(_08617_),
    .B(_08622_),
    .Y(_08638_));
 sky130_fd_sc_hd__nand2_1 _15544_ (.A(_08508_),
    .B(_08512_),
    .Y(_08639_));
 sky130_fd_sc_hd__xor2_1 _15545_ (.A(_08639_),
    .B(_08564_),
    .X(_08640_));
 sky130_fd_sc_hd__a21o_1 _15546_ (.A1(_08620_),
    .A2(_08638_),
    .B1(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__nand3_1 _15547_ (.A(_08620_),
    .B(_08638_),
    .C(_08640_),
    .Y(_08642_));
 sky130_fd_sc_hd__nand2_1 _15548_ (.A(_08641_),
    .B(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__xnor2_2 _15549_ (.A(_08637_),
    .B(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__nor2_1 _15550_ (.A(_08594_),
    .B(_08625_),
    .Y(_08645_));
 sky130_fd_sc_hd__a21oi_1 _15551_ (.A1(_08626_),
    .A2(_08644_),
    .B1(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__xor2_1 _15552_ (.A(_08593_),
    .B(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__or2b_1 _15553_ (.A(_08643_),
    .B_N(_08637_),
    .X(_08648_));
 sky130_fd_sc_hd__a21oi_4 _15554_ (.A1(_08641_),
    .A2(_08648_),
    .B1(_08508_),
    .Y(_08649_));
 sky130_fd_sc_hd__and3_1 _15555_ (.A(_08508_),
    .B(_08641_),
    .C(_08648_),
    .X(_08650_));
 sky130_fd_sc_hd__nor2_1 _15556_ (.A(_08649_),
    .B(_08650_),
    .Y(_08651_));
 sky130_fd_sc_hd__xnor2_1 _15557_ (.A(_08647_),
    .B(_08651_),
    .Y(_08652_));
 sky130_fd_sc_hd__and2b_1 _15558_ (.A_N(_08645_),
    .B(_08626_),
    .X(_08653_));
 sky130_fd_sc_hd__xnor2_2 _15559_ (.A(_08653_),
    .B(_08644_),
    .Y(_08654_));
 sky130_fd_sc_hd__xnor2_1 _15560_ (.A(_08612_),
    .B(_08623_),
    .Y(_08655_));
 sky130_fd_sc_hd__xnor2_2 _15561_ (.A(_08603_),
    .B(_08609_),
    .Y(_08656_));
 sky130_fd_sc_hd__a2bb2o_1 _15562_ (.A1_N(_08370_),
    .A2_N(_08311_),
    .B1(_08598_),
    .B2(_08600_),
    .X(_08657_));
 sky130_fd_sc_hd__or2_1 _15563_ (.A(_08380_),
    .B(_08311_),
    .X(_08658_));
 sky130_fd_sc_hd__and3_1 _15564_ (.A(_08131_),
    .B(_08234_),
    .C(_08367_),
    .X(_08659_));
 sky130_fd_sc_hd__xor2_1 _15565_ (.A(_08597_),
    .B(_08659_),
    .X(_08660_));
 sky130_fd_sc_hd__clkbuf_4 _15566_ (.A(_08368_),
    .X(_08661_));
 sky130_fd_sc_hd__or3_1 _15567_ (.A(_08661_),
    .B(_08351_),
    .C(_08597_),
    .X(_08662_));
 sky130_fd_sc_hd__o21ai_1 _15568_ (.A1(_08658_),
    .A2(_08660_),
    .B1(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__nand3_1 _15569_ (.A(_08601_),
    .B(_08657_),
    .C(_08663_),
    .Y(_08664_));
 sky130_fd_sc_hd__or2_1 _15570_ (.A(_08287_),
    .B(_08417_),
    .X(_08665_));
 sky130_fd_sc_hd__or3_1 _15571_ (.A(_08267_),
    .B(_08381_),
    .C(_08385_),
    .X(_08666_));
 sky130_fd_sc_hd__or3_1 _15572_ (.A(_08259_),
    .B(_08380_),
    .C(_08666_),
    .X(_08667_));
 sky130_fd_sc_hd__o22ai_1 _15573_ (.A1(_08268_),
    .A2(_08380_),
    .B1(_08386_),
    .B2(_08259_),
    .Y(_08668_));
 sky130_fd_sc_hd__and2_1 _15574_ (.A(_08667_),
    .B(_08668_),
    .X(_08669_));
 sky130_fd_sc_hd__xnor2_1 _15575_ (.A(_08665_),
    .B(_08669_),
    .Y(_08670_));
 sky130_fd_sc_hd__a21o_1 _15576_ (.A1(_08601_),
    .A2(_08657_),
    .B1(_08663_),
    .X(_08671_));
 sky130_fd_sc_hd__nand3_1 _15577_ (.A(_08664_),
    .B(_08670_),
    .C(_08671_),
    .Y(_08672_));
 sky130_fd_sc_hd__and2_1 _15578_ (.A(_08664_),
    .B(_08672_),
    .X(_08673_));
 sky130_fd_sc_hd__xor2_1 _15579_ (.A(_08656_),
    .B(_08673_),
    .X(_08674_));
 sky130_fd_sc_hd__nor2_1 _15580_ (.A(_08428_),
    .B(_08522_),
    .Y(_08675_));
 sky130_fd_sc_hd__clkinv_2 _15581_ (.A(_08395_),
    .Y(_08676_));
 sky130_fd_sc_hd__nor2_1 _15582_ (.A(_08471_),
    .B(_08476_),
    .Y(_08677_));
 sky130_fd_sc_hd__clkbuf_4 _15583_ (.A(_08527_),
    .X(_08678_));
 sky130_fd_sc_hd__nor2_1 _15584_ (.A(_08523_),
    .B(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__a22o_1 _15585_ (.A1(_08676_),
    .A2(_08677_),
    .B1(_08679_),
    .B2(_08469_),
    .X(_08680_));
 sky130_fd_sc_hd__or4_1 _15586_ (.A(_08395_),
    .B(_08408_),
    .C(_08477_),
    .D(_08528_),
    .X(_08681_));
 sky130_fd_sc_hd__a21bo_1 _15587_ (.A1(_08675_),
    .A2(_08680_),
    .B1_N(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__or2b_1 _15588_ (.A(_08665_),
    .B_N(_08669_),
    .X(_08683_));
 sky130_fd_sc_hd__xnor2_1 _15589_ (.A(_08615_),
    .B(_08616_),
    .Y(_08684_));
 sky130_fd_sc_hd__a21o_1 _15590_ (.A1(_08667_),
    .A2(_08683_),
    .B1(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__nand3_1 _15591_ (.A(_08667_),
    .B(_08683_),
    .C(_08684_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand2_1 _15592_ (.A(_08685_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__xnor2_1 _15593_ (.A(_08682_),
    .B(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__nor2_1 _15594_ (.A(_08656_),
    .B(_08673_),
    .Y(_08689_));
 sky130_fd_sc_hd__a21oi_1 _15595_ (.A1(_08674_),
    .A2(_08688_),
    .B1(_08689_),
    .Y(_08690_));
 sky130_fd_sc_hd__nor2_1 _15596_ (.A(_08655_),
    .B(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__and2_1 _15597_ (.A(_08655_),
    .B(_08690_),
    .X(_08692_));
 sky130_fd_sc_hd__nor2_1 _15598_ (.A(_08691_),
    .B(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__clkbuf_4 _15599_ (.A(_08631_),
    .X(_08694_));
 sky130_fd_sc_hd__nor2_1 _15600_ (.A(_08559_),
    .B(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__nand2_1 _15601_ (.A(_08628_),
    .B(_08695_),
    .Y(_08696_));
 sky130_fd_sc_hd__a21oi_1 _15602_ (.A1(_08557_),
    .A2(_08628_),
    .B1(_08633_),
    .Y(_08697_));
 sky130_fd_sc_hd__xnor2_1 _15603_ (.A(_08632_),
    .B(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__or2b_1 _15604_ (.A(_08696_),
    .B_N(_08698_),
    .X(_08699_));
 sky130_fd_sc_hd__a21bo_1 _15605_ (.A1(_08682_),
    .A2(_08686_),
    .B1_N(_08685_),
    .X(_08700_));
 sky130_fd_sc_hd__or2_1 _15606_ (.A(_08501_),
    .B(_08635_),
    .X(_08701_));
 sky130_fd_sc_hd__nand2_1 _15607_ (.A(_08636_),
    .B(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__xnor2_2 _15608_ (.A(_08700_),
    .B(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__xnor2_1 _15609_ (.A(_08699_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__a21oi_1 _15610_ (.A1(_08693_),
    .A2(_08704_),
    .B1(_08691_),
    .Y(_08705_));
 sky130_fd_sc_hd__xnor2_2 _15611_ (.A(_08654_),
    .B(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__and3_1 _15612_ (.A(_08628_),
    .B(_08695_),
    .C(_08698_),
    .X(_08707_));
 sky130_fd_sc_hd__a32oi_4 _15613_ (.A1(_08636_),
    .A2(_08700_),
    .A3(_08701_),
    .B1(_08703_),
    .B2(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__or2_1 _15614_ (.A(_08654_),
    .B(_08705_),
    .X(_08709_));
 sky130_fd_sc_hd__o21a_1 _15615_ (.A1(_08706_),
    .A2(_08708_),
    .B1(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__nor2_1 _15616_ (.A(_08652_),
    .B(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__and2_1 _15617_ (.A(_08652_),
    .B(_08710_),
    .X(_08712_));
 sky130_fd_sc_hd__or2_1 _15618_ (.A(_08711_),
    .B(_08712_),
    .X(_08713_));
 sky130_fd_sc_hd__and2_1 _15619_ (.A(_08681_),
    .B(_08680_),
    .X(_08714_));
 sky130_fd_sc_hd__xnor2_1 _15620_ (.A(_08675_),
    .B(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__nand2_1 _15621_ (.A(_08260_),
    .B(_08468_),
    .Y(_08716_));
 sky130_fd_sc_hd__xor2_1 _15622_ (.A(_08666_),
    .B(_08716_),
    .X(_08717_));
 sky130_fd_sc_hd__nor2_1 _15623_ (.A(_08287_),
    .B(_08478_),
    .Y(_08718_));
 sky130_fd_sc_hd__a2bb2o_1 _15624_ (.A1_N(_08666_),
    .A2_N(_08716_),
    .B1(_08717_),
    .B2(_08718_),
    .X(_08719_));
 sky130_fd_sc_hd__or2b_1 _15625_ (.A(_08715_),
    .B_N(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__xor2_1 _15626_ (.A(_08719_),
    .B(_08715_),
    .X(_08721_));
 sky130_fd_sc_hd__nand2_1 _15627_ (.A(_08676_),
    .B(_08679_),
    .Y(_08722_));
 sky130_fd_sc_hd__or2_1 _15628_ (.A(_08408_),
    .B(_08521_),
    .X(_08723_));
 sky130_fd_sc_hd__nor2_1 _15629_ (.A(_08429_),
    .B(_08555_),
    .Y(_08724_));
 sky130_fd_sc_hd__xor2_1 _15630_ (.A(_08722_),
    .B(_08723_),
    .X(_08725_));
 sky130_fd_sc_hd__a2bb2o_1 _15631_ (.A1_N(_08722_),
    .A2_N(_08723_),
    .B1(_08724_),
    .B2(_08725_),
    .X(_08726_));
 sky130_fd_sc_hd__or2b_1 _15632_ (.A(_08721_),
    .B_N(_08726_),
    .X(_08727_));
 sky130_fd_sc_hd__a21o_1 _15633_ (.A1(_08628_),
    .A2(_08695_),
    .B1(_08698_),
    .X(_08728_));
 sky130_fd_sc_hd__nand2_1 _15634_ (.A(_08699_),
    .B(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__a21oi_2 _15635_ (.A1(_08720_),
    .A2(_08727_),
    .B1(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__xnor2_1 _15636_ (.A(_08693_),
    .B(_08704_),
    .Y(_08731_));
 sky130_fd_sc_hd__xnor2_1 _15637_ (.A(_08674_),
    .B(_08688_),
    .Y(_08732_));
 sky130_fd_sc_hd__a21o_1 _15638_ (.A1(_08664_),
    .A2(_08671_),
    .B1(_08670_),
    .X(_08733_));
 sky130_fd_sc_hd__xor2_1 _15639_ (.A(_08718_),
    .B(_08717_),
    .X(_08734_));
 sky130_fd_sc_hd__xnor2_1 _15640_ (.A(_08658_),
    .B(_08660_),
    .Y(_08735_));
 sky130_fd_sc_hd__or3_1 _15641_ (.A(_08381_),
    .B(_08385_),
    .C(_08311_),
    .X(_08736_));
 sky130_fd_sc_hd__o21ai_4 _15642_ (.A1(\rbzero.wall_tracer.stepDistY[-4] ),
    .A2(_08309_),
    .B1(_08379_),
    .Y(_08737_));
 sky130_fd_sc_hd__o22a_1 _15643_ (.A1(_08661_),
    .A2(_08354_),
    .B1(_08351_),
    .B2(_08737_),
    .X(_08738_));
 sky130_fd_sc_hd__or3b_1 _15644_ (.A(_08737_),
    .B(_08354_),
    .C_N(_08659_),
    .X(_08739_));
 sky130_fd_sc_hd__o21a_1 _15645_ (.A1(_08736_),
    .A2(_08738_),
    .B1(_08739_),
    .X(_08740_));
 sky130_fd_sc_hd__nand2_1 _15646_ (.A(_08735_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__nor2_1 _15647_ (.A(_08735_),
    .B(_08740_),
    .Y(_08742_));
 sky130_fd_sc_hd__a21o_1 _15648_ (.A1(_08734_),
    .A2(_08741_),
    .B1(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__nand3_1 _15649_ (.A(_08672_),
    .B(_08733_),
    .C(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__xnor2_1 _15650_ (.A(_08726_),
    .B(_08721_),
    .Y(_08745_));
 sky130_fd_sc_hd__a21o_1 _15651_ (.A1(_08672_),
    .A2(_08733_),
    .B1(_08743_),
    .X(_08746_));
 sky130_fd_sc_hd__nand3_1 _15652_ (.A(_08744_),
    .B(_08745_),
    .C(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__and2_1 _15653_ (.A(_08744_),
    .B(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__xor2_1 _15654_ (.A(_08732_),
    .B(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__and3_1 _15655_ (.A(_08720_),
    .B(_08727_),
    .C(_08729_),
    .X(_08750_));
 sky130_fd_sc_hd__nor2_1 _15656_ (.A(_08730_),
    .B(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__nor2_1 _15657_ (.A(_08732_),
    .B(_08748_),
    .Y(_08752_));
 sky130_fd_sc_hd__a21oi_1 _15658_ (.A1(_08749_),
    .A2(_08751_),
    .B1(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__xor2_1 _15659_ (.A(_08731_),
    .B(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__xnor2_1 _15660_ (.A(_08730_),
    .B(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__nand2_1 _15661_ (.A(_08269_),
    .B(_08468_),
    .Y(_08756_));
 sky130_fd_sc_hd__nand2_1 _15662_ (.A(_08260_),
    .B(_08677_),
    .Y(_08757_));
 sky130_fd_sc_hd__xor2_1 _15663_ (.A(_08756_),
    .B(_08757_),
    .X(_08758_));
 sky130_fd_sc_hd__nor2_1 _15664_ (.A(_08288_),
    .B(_08529_),
    .Y(_08759_));
 sky130_fd_sc_hd__a2bb2oi_1 _15665_ (.A1_N(_08756_),
    .A2_N(_08757_),
    .B1(_08758_),
    .B2(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__xnor2_1 _15666_ (.A(_08724_),
    .B(_08725_),
    .Y(_08761_));
 sky130_fd_sc_hd__or2_1 _15667_ (.A(_08760_),
    .B(_08761_),
    .X(_08762_));
 sky130_fd_sc_hd__xnor2_1 _15668_ (.A(_08760_),
    .B(_08761_),
    .Y(_08763_));
 sky130_fd_sc_hd__nor2_1 _15669_ (.A(_08429_),
    .B(_08694_),
    .Y(_08764_));
 sky130_fd_sc_hd__a211o_1 _15670_ (.A1(_08554_),
    .A2(_08231_),
    .B1(_08505_),
    .C1(_08408_),
    .X(_08765_));
 sky130_fd_sc_hd__o21ai_1 _15671_ (.A1(_08396_),
    .A2(_08522_),
    .B1(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__or3_1 _15672_ (.A(_08396_),
    .B(_08521_),
    .C(_08765_),
    .X(_08767_));
 sky130_fd_sc_hd__a21bo_1 _15673_ (.A1(_08764_),
    .A2(_08766_),
    .B1_N(_08767_),
    .X(_08768_));
 sky130_fd_sc_hd__or2b_1 _15674_ (.A(_08763_),
    .B_N(_08768_),
    .X(_08769_));
 sky130_fd_sc_hd__or2_1 _15675_ (.A(_08628_),
    .B(_08695_),
    .X(_08770_));
 sky130_fd_sc_hd__nand2_1 _15676_ (.A(_08696_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__a21oi_1 _15677_ (.A1(_08762_),
    .A2(_08769_),
    .B1(_08771_),
    .Y(_08772_));
 sky130_fd_sc_hd__xnor2_1 _15678_ (.A(_08749_),
    .B(_08751_),
    .Y(_08773_));
 sky130_fd_sc_hd__a21o_1 _15679_ (.A1(_08744_),
    .A2(_08746_),
    .B1(_08745_),
    .X(_08774_));
 sky130_fd_sc_hd__xnor2_1 _15680_ (.A(_08768_),
    .B(_08763_),
    .Y(_08775_));
 sky130_fd_sc_hd__and2b_1 _15681_ (.A_N(_08742_),
    .B(_08741_),
    .X(_08776_));
 sky130_fd_sc_hd__xnor2_1 _15682_ (.A(_08734_),
    .B(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__xor2_1 _15683_ (.A(_08759_),
    .B(_08758_),
    .X(_08778_));
 sky130_fd_sc_hd__inv_2 _15684_ (.A(_08737_),
    .Y(_08779_));
 sky130_fd_sc_hd__a31o_1 _15685_ (.A1(_08779_),
    .A2(_08349_),
    .A3(_08659_),
    .B1(_08738_),
    .X(_08780_));
 sky130_fd_sc_hd__xnor2_1 _15686_ (.A(_08736_),
    .B(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__or4_1 _15687_ (.A(_08737_),
    .B(_08385_),
    .C(_08353_),
    .D(_08351_),
    .X(_08782_));
 sky130_fd_sc_hd__clkbuf_4 _15688_ (.A(_08385_),
    .X(_08783_));
 sky130_fd_sc_hd__o22ai_1 _15689_ (.A1(_08737_),
    .A2(_08354_),
    .B1(_08351_),
    .B2(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__nand4_1 _15690_ (.A(_08468_),
    .B(_08350_),
    .C(_08782_),
    .D(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__and2_1 _15691_ (.A(_08782_),
    .B(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__xor2_1 _15692_ (.A(_08781_),
    .B(_08786_),
    .X(_08787_));
 sky130_fd_sc_hd__nor2_1 _15693_ (.A(_08781_),
    .B(_08786_),
    .Y(_08788_));
 sky130_fd_sc_hd__a21oi_1 _15694_ (.A1(_08778_),
    .A2(_08787_),
    .B1(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__xor2_1 _15695_ (.A(_08777_),
    .B(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__nor2_1 _15696_ (.A(_08777_),
    .B(_08789_),
    .Y(_08791_));
 sky130_fd_sc_hd__a21o_1 _15697_ (.A1(_08775_),
    .A2(_08790_),
    .B1(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__a21o_1 _15698_ (.A1(_08747_),
    .A2(_08774_),
    .B1(_08792_),
    .X(_08793_));
 sky130_fd_sc_hd__and3_1 _15699_ (.A(_08762_),
    .B(_08769_),
    .C(_08771_),
    .X(_08794_));
 sky130_fd_sc_hd__nor2_1 _15700_ (.A(_08772_),
    .B(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand3_1 _15701_ (.A(_08747_),
    .B(_08774_),
    .C(_08792_),
    .Y(_08796_));
 sky130_fd_sc_hd__a21boi_1 _15702_ (.A1(_08793_),
    .A2(_08795_),
    .B1_N(_08796_),
    .Y(_08797_));
 sky130_fd_sc_hd__xor2_1 _15703_ (.A(_08773_),
    .B(_08797_),
    .X(_08798_));
 sky130_fd_sc_hd__nor2_1 _15704_ (.A(_08773_),
    .B(_08797_),
    .Y(_08799_));
 sky130_fd_sc_hd__a21oi_1 _15705_ (.A1(_08772_),
    .A2(_08798_),
    .B1(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__nor2_1 _15706_ (.A(_08755_),
    .B(_08800_),
    .Y(_08801_));
 sky130_fd_sc_hd__xnor2_2 _15707_ (.A(_08706_),
    .B(_08708_),
    .Y(_08802_));
 sky130_fd_sc_hd__nor2_1 _15708_ (.A(_08731_),
    .B(_08753_),
    .Y(_08803_));
 sky130_fd_sc_hd__a21oi_2 _15709_ (.A1(_08730_),
    .A2(_08754_),
    .B1(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__xor2_2 _15710_ (.A(_08802_),
    .B(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__nand2_1 _15711_ (.A(_08801_),
    .B(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__xnor2_1 _15712_ (.A(_08772_),
    .B(_08798_),
    .Y(_08807_));
 sky130_fd_sc_hd__clkbuf_4 _15713_ (.A(_08547_),
    .X(_08808_));
 sky130_fd_sc_hd__buf_4 _15714_ (.A(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__or2_1 _15715_ (.A(_08809_),
    .B(_08694_),
    .X(_08810_));
 sky130_fd_sc_hd__or2_1 _15716_ (.A(_08288_),
    .B(_08522_),
    .X(_08811_));
 sky130_fd_sc_hd__o22a_1 _15717_ (.A1(_08268_),
    .A2(_08478_),
    .B1(_08529_),
    .B2(_08272_),
    .X(_08812_));
 sky130_fd_sc_hd__or4_1 _15718_ (.A(_08259_),
    .B(_08268_),
    .C(_08477_),
    .D(_08528_),
    .X(_08813_));
 sky130_fd_sc_hd__o21ai_1 _15719_ (.A1(_08811_),
    .A2(_08812_),
    .B1(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__and2_1 _15720_ (.A(_08767_),
    .B(_08766_),
    .X(_08815_));
 sky130_fd_sc_hd__xor2_1 _15721_ (.A(_08764_),
    .B(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__xnor2_1 _15722_ (.A(_08814_),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__or2_2 _15723_ (.A(_08438_),
    .B(_08694_),
    .X(_08818_));
 sky130_fd_sc_hd__nand2_1 _15724_ (.A(_08814_),
    .B(_08816_),
    .Y(_08819_));
 sky130_fd_sc_hd__o31a_1 _15725_ (.A1(_08765_),
    .A2(_08817_),
    .A3(_08818_),
    .B1(_08819_),
    .X(_08820_));
 sky130_fd_sc_hd__nor2_1 _15726_ (.A(_08810_),
    .B(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__and3_1 _15727_ (.A(_08796_),
    .B(_08793_),
    .C(_08795_),
    .X(_08822_));
 sky130_fd_sc_hd__a21oi_1 _15728_ (.A1(_08796_),
    .A2(_08793_),
    .B1(_08795_),
    .Y(_08823_));
 sky130_fd_sc_hd__or2_1 _15729_ (.A(_08822_),
    .B(_08823_),
    .X(_08824_));
 sky130_fd_sc_hd__xnor2_1 _15730_ (.A(_08775_),
    .B(_08790_),
    .Y(_08825_));
 sky130_fd_sc_hd__nor2_1 _15731_ (.A(_08765_),
    .B(_08818_),
    .Y(_08826_));
 sky130_fd_sc_hd__xnor2_1 _15732_ (.A(_08817_),
    .B(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__xnor2_1 _15733_ (.A(_08778_),
    .B(_08787_),
    .Y(_08828_));
 sky130_fd_sc_hd__a22o_1 _15734_ (.A1(_08468_),
    .A2(_08350_),
    .B1(_08782_),
    .B2(_08784_),
    .X(_08829_));
 sky130_fd_sc_hd__clkbuf_4 _15735_ (.A(_08351_),
    .X(_08830_));
 sky130_fd_sc_hd__clkbuf_4 _15736_ (.A(_08415_),
    .X(_08831_));
 sky130_fd_sc_hd__or2_1 _15737_ (.A(_08831_),
    .B(_08354_),
    .X(_08832_));
 sky130_fd_sc_hd__nor3_1 _15738_ (.A(_08783_),
    .B(_08830_),
    .C(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__or4_1 _15739_ (.A(_08385_),
    .B(_08415_),
    .C(_08354_),
    .D(_08351_),
    .X(_08834_));
 sky130_fd_sc_hd__o22ai_1 _15740_ (.A1(_08783_),
    .A2(_08354_),
    .B1(_08351_),
    .B2(_08415_),
    .Y(_08835_));
 sky130_fd_sc_hd__and4_1 _15741_ (.A(_08677_),
    .B(_08350_),
    .C(_08834_),
    .D(_08835_),
    .X(_08836_));
 sky130_fd_sc_hd__or2_1 _15742_ (.A(_08833_),
    .B(_08836_),
    .X(_08837_));
 sky130_fd_sc_hd__and2b_1 _15743_ (.A_N(_08812_),
    .B(_08813_),
    .X(_08838_));
 sky130_fd_sc_hd__xnor2_1 _15744_ (.A(_08811_),
    .B(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__nand2_1 _15745_ (.A(_08785_),
    .B(_08829_),
    .Y(_08840_));
 sky130_fd_sc_hd__xnor2_1 _15746_ (.A(_08840_),
    .B(_08837_),
    .Y(_08841_));
 sky130_fd_sc_hd__a32o_1 _15747_ (.A1(_08785_),
    .A2(_08829_),
    .A3(_08837_),
    .B1(_08839_),
    .B2(_08841_),
    .X(_08842_));
 sky130_fd_sc_hd__xnor2_1 _15748_ (.A(_08828_),
    .B(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__and2b_1 _15749_ (.A_N(_08828_),
    .B(_08842_),
    .X(_08844_));
 sky130_fd_sc_hd__a21oi_1 _15750_ (.A1(_08827_),
    .A2(_08843_),
    .B1(_08844_),
    .Y(_08845_));
 sky130_fd_sc_hd__and2_1 _15751_ (.A(_08810_),
    .B(_08820_),
    .X(_08846_));
 sky130_fd_sc_hd__nor2_1 _15752_ (.A(_08821_),
    .B(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__xor2_1 _15753_ (.A(_08825_),
    .B(_08845_),
    .X(_08848_));
 sky130_fd_sc_hd__nand2_1 _15754_ (.A(_08847_),
    .B(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__o21a_1 _15755_ (.A1(_08825_),
    .A2(_08845_),
    .B1(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__xor2_1 _15756_ (.A(_08824_),
    .B(_08850_),
    .X(_08851_));
 sky130_fd_sc_hd__nor2_1 _15757_ (.A(_08824_),
    .B(_08850_),
    .Y(_08852_));
 sky130_fd_sc_hd__a21oi_1 _15758_ (.A1(_08821_),
    .A2(_08851_),
    .B1(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__nor2_1 _15759_ (.A(_08807_),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__xor2_1 _15760_ (.A(_08755_),
    .B(_08800_),
    .X(_08855_));
 sky130_fd_sc_hd__and2_1 _15761_ (.A(_08854_),
    .B(_08855_),
    .X(_08856_));
 sky130_fd_sc_hd__xor2_1 _15762_ (.A(_08807_),
    .B(_08853_),
    .X(_08857_));
 sky130_fd_sc_hd__xor2_1 _15763_ (.A(_08821_),
    .B(_08851_),
    .X(_08858_));
 sky130_fd_sc_hd__xnor2_1 _15764_ (.A(_08827_),
    .B(_08843_),
    .Y(_08859_));
 sky130_fd_sc_hd__nand2_1 _15765_ (.A(_08839_),
    .B(_08841_),
    .Y(_08860_));
 sky130_fd_sc_hd__or2_1 _15766_ (.A(_08839_),
    .B(_08841_),
    .X(_08861_));
 sky130_fd_sc_hd__o2bb2a_1 _15767_ (.A1_N(_08834_),
    .A2_N(_08835_),
    .B1(_08478_),
    .B2(_08311_),
    .X(_08862_));
 sky130_fd_sc_hd__or2_1 _15768_ (.A(_08836_),
    .B(_08862_),
    .X(_08863_));
 sky130_fd_sc_hd__nor2_1 _15769_ (.A(_08529_),
    .B(_08312_),
    .Y(_08864_));
 sky130_fd_sc_hd__or2_1 _15770_ (.A(_08476_),
    .B(_08830_),
    .X(_08865_));
 sky130_fd_sc_hd__nand2_1 _15771_ (.A(_08832_),
    .B(_08865_),
    .Y(_08866_));
 sky130_fd_sc_hd__nor3_1 _15772_ (.A(_08341_),
    .B(_08831_),
    .C(_08865_),
    .Y(_08867_));
 sky130_fd_sc_hd__a21oi_1 _15773_ (.A1(_08864_),
    .A2(_08866_),
    .B1(_08867_),
    .Y(_08868_));
 sky130_fd_sc_hd__nor2_1 _15774_ (.A(_08863_),
    .B(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__and2_1 _15775_ (.A(_08863_),
    .B(_08868_),
    .X(_08870_));
 sky130_fd_sc_hd__nor2_1 _15776_ (.A(_08869_),
    .B(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__or2_1 _15777_ (.A(_08288_),
    .B(_08555_),
    .X(_08872_));
 sky130_fd_sc_hd__nand2_1 _15778_ (.A(_08260_),
    .B(_08679_),
    .Y(_08873_));
 sky130_fd_sc_hd__or2_2 _15779_ (.A(_08271_),
    .B(_08522_),
    .X(_08874_));
 sky130_fd_sc_hd__or2_1 _15780_ (.A(_08259_),
    .B(_08521_),
    .X(_08875_));
 sky130_fd_sc_hd__o21a_1 _15781_ (.A1(_08271_),
    .A2(_08529_),
    .B1(_08875_),
    .X(_08876_));
 sky130_fd_sc_hd__o21ba_1 _15782_ (.A1(_08873_),
    .A2(_08874_),
    .B1_N(_08876_),
    .X(_08877_));
 sky130_fd_sc_hd__xnor2_1 _15783_ (.A(_08872_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__a21o_1 _15784_ (.A1(_08871_),
    .A2(_08878_),
    .B1(_08869_),
    .X(_08879_));
 sky130_fd_sc_hd__nand2_1 _15785_ (.A(_08860_),
    .B(_08861_),
    .Y(_08880_));
 sky130_fd_sc_hd__xnor2_1 _15786_ (.A(_08880_),
    .B(_08879_),
    .Y(_08881_));
 sky130_fd_sc_hd__o22ai_4 _15787_ (.A1(_08872_),
    .A2(_08876_),
    .B1(_08874_),
    .B2(_08873_),
    .Y(_08882_));
 sky130_fd_sc_hd__o22a_1 _15788_ (.A1(_08438_),
    .A2(_08555_),
    .B1(_08694_),
    .B2(_08409_),
    .X(_08883_));
 sky130_fd_sc_hd__or2_1 _15789_ (.A(_08826_),
    .B(_08883_),
    .X(_08884_));
 sky130_fd_sc_hd__xnor2_1 _15790_ (.A(_08882_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__a32oi_2 _15791_ (.A1(_08860_),
    .A2(_08861_),
    .A3(_08879_),
    .B1(_08881_),
    .B2(_08885_),
    .Y(_08886_));
 sky130_fd_sc_hd__or2_1 _15792_ (.A(_08859_),
    .B(_08886_),
    .X(_08887_));
 sky130_fd_sc_hd__xnor2_1 _15793_ (.A(_08859_),
    .B(_08886_),
    .Y(_08888_));
 sky130_fd_sc_hd__or3b_1 _15794_ (.A(_08884_),
    .B(_08888_),
    .C_N(_08882_),
    .X(_08889_));
 sky130_fd_sc_hd__or2_1 _15795_ (.A(_08847_),
    .B(_08848_),
    .X(_08890_));
 sky130_fd_sc_hd__nand2_1 _15796_ (.A(_08849_),
    .B(_08890_),
    .Y(_08891_));
 sky130_fd_sc_hd__a21o_1 _15797_ (.A1(_08887_),
    .A2(_08889_),
    .B1(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__inv_2 _15798_ (.A(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__and3_1 _15799_ (.A(_08857_),
    .B(_08858_),
    .C(_08893_),
    .X(_08894_));
 sky130_fd_sc_hd__nor2_1 _15800_ (.A(_08854_),
    .B(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__xnor2_1 _15801_ (.A(_08855_),
    .B(_08895_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand2_1 _15802_ (.A(_08858_),
    .B(_08893_),
    .Y(_08897_));
 sky130_fd_sc_hd__xor2_1 _15803_ (.A(_08857_),
    .B(_08897_),
    .X(_08898_));
 sky130_fd_sc_hd__nand2_1 _15804_ (.A(_08891_),
    .B(_08887_),
    .Y(_08899_));
 sky130_fd_sc_hd__xnor2_1 _15805_ (.A(_08881_),
    .B(_08885_),
    .Y(_08900_));
 sky130_fd_sc_hd__xnor2_1 _15806_ (.A(_08871_),
    .B(_08878_),
    .Y(_08901_));
 sky130_fd_sc_hd__or2_1 _15807_ (.A(_08288_),
    .B(_08694_),
    .X(_08902_));
 sky130_fd_sc_hd__nor2_1 _15808_ (.A(_08272_),
    .B(_08555_),
    .Y(_08903_));
 sky130_fd_sc_hd__xnor2_1 _15809_ (.A(_08874_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__xnor2_1 _15810_ (.A(_08902_),
    .B(_08904_),
    .Y(_08905_));
 sky130_fd_sc_hd__and2b_1 _15811_ (.A_N(_08867_),
    .B(_08866_),
    .X(_08906_));
 sky130_fd_sc_hd__xnor2_1 _15812_ (.A(_08864_),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__or2_1 _15813_ (.A(_08522_),
    .B(_08312_),
    .X(_08908_));
 sky130_fd_sc_hd__or3_1 _15814_ (.A(_08341_),
    .B(_08678_),
    .C(_08865_),
    .X(_08909_));
 sky130_fd_sc_hd__o22ai_1 _15815_ (.A1(_08476_),
    .A2(_08354_),
    .B1(_08830_),
    .B2(_08678_),
    .Y(_08910_));
 sky130_fd_sc_hd__nand2_1 _15816_ (.A(_08909_),
    .B(_08910_),
    .Y(_08911_));
 sky130_fd_sc_hd__o21a_1 _15817_ (.A1(_08908_),
    .A2(_08911_),
    .B1(_08909_),
    .X(_08912_));
 sky130_fd_sc_hd__nor2_1 _15818_ (.A(_08907_),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__and2_1 _15819_ (.A(_08907_),
    .B(_08912_),
    .X(_08914_));
 sky130_fd_sc_hd__nor2_1 _15820_ (.A(_08913_),
    .B(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__a21oi_1 _15821_ (.A1(_08905_),
    .A2(_08915_),
    .B1(_08913_),
    .Y(_08916_));
 sky130_fd_sc_hd__xor2_1 _15822_ (.A(_08901_),
    .B(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__clkbuf_4 _15823_ (.A(_08271_),
    .X(_08918_));
 sky130_fd_sc_hd__or2_1 _15824_ (.A(_08918_),
    .B(_08555_),
    .X(_08919_));
 sky130_fd_sc_hd__or2b_1 _15825_ (.A(_08902_),
    .B_N(_08904_),
    .X(_08920_));
 sky130_fd_sc_hd__o21a_1 _15826_ (.A1(_08875_),
    .A2(_08919_),
    .B1(_08920_),
    .X(_08921_));
 sky130_fd_sc_hd__or2_1 _15827_ (.A(_08818_),
    .B(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__nand2_1 _15828_ (.A(_08818_),
    .B(_08921_),
    .Y(_08923_));
 sky130_fd_sc_hd__and2_1 _15829_ (.A(_08922_),
    .B(_08923_),
    .X(_08924_));
 sky130_fd_sc_hd__nand2_1 _15830_ (.A(_08917_),
    .B(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__o21a_1 _15831_ (.A1(_08901_),
    .A2(_08916_),
    .B1(_08925_),
    .X(_08926_));
 sky130_fd_sc_hd__or2_1 _15832_ (.A(_08900_),
    .B(_08926_),
    .X(_08927_));
 sky130_fd_sc_hd__xnor2_1 _15833_ (.A(_08900_),
    .B(_08926_),
    .Y(_08928_));
 sky130_fd_sc_hd__or2_1 _15834_ (.A(_08922_),
    .B(_08928_),
    .X(_08929_));
 sky130_fd_sc_hd__and2b_1 _15835_ (.A_N(_08884_),
    .B(_08882_),
    .X(_08930_));
 sky130_fd_sc_hd__xor2_1 _15836_ (.A(_08930_),
    .B(_08888_),
    .X(_08931_));
 sky130_fd_sc_hd__a21oi_1 _15837_ (.A1(_08927_),
    .A2(_08929_),
    .B1(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__and4_1 _15838_ (.A(_08858_),
    .B(_08892_),
    .C(_08899_),
    .D(_08932_),
    .X(_08933_));
 sky130_fd_sc_hd__xnor2_1 _15839_ (.A(_08898_),
    .B(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__inv_2 _15840_ (.A(_08889_),
    .Y(_08935_));
 sky130_fd_sc_hd__o22a_1 _15841_ (.A1(_08935_),
    .A2(_08899_),
    .B1(_08927_),
    .B2(_08931_),
    .X(_08936_));
 sky130_fd_sc_hd__or2_1 _15842_ (.A(_08917_),
    .B(_08924_),
    .X(_08937_));
 sky130_fd_sc_hd__nand2_1 _15843_ (.A(_08925_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__xnor2_1 _15844_ (.A(_08905_),
    .B(_08915_),
    .Y(_08939_));
 sky130_fd_sc_hd__xnor2_1 _15845_ (.A(_08908_),
    .B(_08911_),
    .Y(_08940_));
 sky130_fd_sc_hd__clkbuf_4 _15846_ (.A(_08312_),
    .X(_08941_));
 sky130_fd_sc_hd__o22a_1 _15847_ (.A1(_08678_),
    .A2(_08354_),
    .B1(_08830_),
    .B2(_08567_),
    .X(_08942_));
 sky130_fd_sc_hd__nor2_1 _15848_ (.A(_08520_),
    .B(_08354_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand2_1 _15849_ (.A(_08355_),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__or2_1 _15850_ (.A(_08678_),
    .B(_08944_),
    .X(_08945_));
 sky130_fd_sc_hd__o31a_1 _15851_ (.A1(_08555_),
    .A2(_08941_),
    .A3(_08942_),
    .B1(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__xor2_1 _15852_ (.A(_08940_),
    .B(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__nor2_1 _15853_ (.A(_08362_),
    .B(_08694_),
    .Y(_08948_));
 sky130_fd_sc_hd__xnor2_1 _15854_ (.A(_08919_),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__nand2_1 _15855_ (.A(_08947_),
    .B(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__o21a_1 _15856_ (.A1(_08940_),
    .A2(_08946_),
    .B1(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__nor2_1 _15857_ (.A(_08918_),
    .B(_08694_),
    .Y(_08952_));
 sky130_fd_sc_hd__xor2_1 _15858_ (.A(_08939_),
    .B(_08951_),
    .X(_08953_));
 sky130_fd_sc_hd__and3_1 _15859_ (.A(_08903_),
    .B(_08952_),
    .C(_08953_),
    .X(_08954_));
 sky130_fd_sc_hd__o21ba_1 _15860_ (.A1(_08939_),
    .A2(_08951_),
    .B1_N(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__or2_1 _15861_ (.A(_08947_),
    .B(_08949_),
    .X(_08956_));
 sky130_fd_sc_hd__nand2_1 _15862_ (.A(_08950_),
    .B(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__nor2_1 _15863_ (.A(_08555_),
    .B(_08941_),
    .Y(_08958_));
 sky130_fd_sc_hd__clkbuf_4 _15864_ (.A(_08678_),
    .X(_08959_));
 sky130_fd_sc_hd__o21ba_1 _15865_ (.A1(_08959_),
    .A2(_08944_),
    .B1_N(_08942_),
    .X(_08960_));
 sky130_fd_sc_hd__xnor2_1 _15866_ (.A(_08958_),
    .B(_08960_),
    .Y(_08961_));
 sky130_fd_sc_hd__nor2_1 _15867_ (.A(_08505_),
    .B(_08830_),
    .Y(_08962_));
 sky130_fd_sc_hd__xnor2_1 _15868_ (.A(_08943_),
    .B(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__or3_1 _15869_ (.A(_08694_),
    .B(_08941_),
    .C(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__a21boi_1 _15870_ (.A1(_08943_),
    .A2(_08962_),
    .B1_N(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__nor2_1 _15871_ (.A(_08961_),
    .B(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__and2_1 _15872_ (.A(_08961_),
    .B(_08965_),
    .X(_08967_));
 sky130_fd_sc_hd__nor2_1 _15873_ (.A(_08966_),
    .B(_08967_),
    .Y(_08968_));
 sky130_fd_sc_hd__and2_1 _15874_ (.A(_08952_),
    .B(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__nor2_1 _15875_ (.A(_08966_),
    .B(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__and3_1 _15876_ (.A(_08630_),
    .B(_08342_),
    .C(_08962_),
    .X(_08971_));
 sky130_fd_sc_hd__o21ai_1 _15877_ (.A1(_08694_),
    .A2(_08941_),
    .B1(_08963_),
    .Y(_08972_));
 sky130_fd_sc_hd__o2111a_1 _15878_ (.A1(_08952_),
    .A2(_08968_),
    .B1(_08971_),
    .C1(_08972_),
    .D1(_08964_),
    .X(_08973_));
 sky130_fd_sc_hd__a21bo_1 _15879_ (.A1(_08957_),
    .A2(_08970_),
    .B1_N(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__o22a_1 _15880_ (.A1(_08957_),
    .A2(_08970_),
    .B1(_08974_),
    .B2(_08969_),
    .X(_08975_));
 sky130_fd_sc_hd__a21oi_1 _15881_ (.A1(_08903_),
    .A2(_08952_),
    .B1(_08953_),
    .Y(_08976_));
 sky130_fd_sc_hd__a211o_1 _15882_ (.A1(_08938_),
    .A2(_08955_),
    .B1(_08976_),
    .C1(_08954_),
    .X(_08977_));
 sky130_fd_sc_hd__o22a_1 _15883_ (.A1(_08938_),
    .A2(_08955_),
    .B1(_08975_),
    .B2(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__a21oi_1 _15884_ (.A1(_08931_),
    .A2(_08927_),
    .B1(_08893_),
    .Y(_08979_));
 sky130_fd_sc_hd__nand2_1 _15885_ (.A(_08922_),
    .B(_08928_),
    .Y(_08980_));
 sky130_fd_sc_hd__and4b_1 _15886_ (.A_N(_08978_),
    .B(_08979_),
    .C(_08980_),
    .D(_08929_),
    .X(_08981_));
 sky130_fd_sc_hd__and3_1 _15887_ (.A(_08858_),
    .B(_08936_),
    .C(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__and2b_1 _15888_ (.A_N(_08898_),
    .B(_08933_),
    .X(_08983_));
 sky130_fd_sc_hd__a21o_1 _15889_ (.A1(_08934_),
    .A2(_08982_),
    .B1(_08983_),
    .X(_08984_));
 sky130_fd_sc_hd__a22o_2 _15890_ (.A1(_08855_),
    .A2(_08894_),
    .B1(_08896_),
    .B2(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__nor2_1 _15891_ (.A(_08801_),
    .B(_08856_),
    .Y(_08986_));
 sky130_fd_sc_hd__xnor2_2 _15892_ (.A(_08805_),
    .B(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__a22o_2 _15893_ (.A1(_08805_),
    .A2(_08856_),
    .B1(_08985_),
    .B2(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__nor2_1 _15894_ (.A(_08802_),
    .B(_08804_),
    .Y(_08989_));
 sky130_fd_sc_hd__inv_2 _15895_ (.A(_08989_),
    .Y(_08990_));
 sky130_fd_sc_hd__nand2_1 _15896_ (.A(_08990_),
    .B(_08806_),
    .Y(_08991_));
 sky130_fd_sc_hd__xnor2_2 _15897_ (.A(_08713_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__a2bb2o_2 _15898_ (.A1_N(_08713_),
    .A2_N(_08806_),
    .B1(_08988_),
    .B2(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__nand2_1 _15899_ (.A(_08437_),
    .B(_08441_),
    .Y(_08994_));
 sky130_fd_sc_hd__or2_1 _15900_ (.A(_08288_),
    .B(_08295_),
    .X(_08995_));
 sky130_fd_sc_hd__o21ba_1 _15901_ (.A1(_08273_),
    .A2(_08995_),
    .B1_N(_08270_),
    .X(_08996_));
 sky130_fd_sc_hd__or2_1 _15902_ (.A(_08396_),
    .B(_08294_),
    .X(_08997_));
 sky130_fd_sc_hd__xnor2_1 _15903_ (.A(_08436_),
    .B(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__or3_1 _15904_ (.A(_08430_),
    .B(_08429_),
    .C(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__o21ai_1 _15905_ (.A1(_08430_),
    .A2(_08429_),
    .B1(_08998_),
    .Y(_09000_));
 sky130_fd_sc_hd__nand2_1 _15906_ (.A(_08999_),
    .B(_09000_),
    .Y(_09001_));
 sky130_fd_sc_hd__or2_1 _15907_ (.A(_08996_),
    .B(_09001_),
    .X(_09002_));
 sky130_fd_sc_hd__nand2_1 _15908_ (.A(_08996_),
    .B(_09001_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand2_1 _15909_ (.A(_09002_),
    .B(_09003_),
    .Y(_09004_));
 sky130_fd_sc_hd__xnor2_1 _15910_ (.A(_08994_),
    .B(_09004_),
    .Y(_09005_));
 sky130_fd_sc_hd__or4_1 _15911_ (.A(_08272_),
    .B(_08271_),
    .C(_08233_),
    .D(_08306_),
    .X(_09006_));
 sky130_fd_sc_hd__clkbuf_4 _15912_ (.A(_08233_),
    .X(_09007_));
 sky130_fd_sc_hd__o22ai_1 _15913_ (.A1(_08362_),
    .A2(_09007_),
    .B1(_08307_),
    .B2(_08918_),
    .Y(_09008_));
 sky130_fd_sc_hd__nand2_1 _15914_ (.A(_09006_),
    .B(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__nor2_1 _15915_ (.A(_08288_),
    .B(_08244_),
    .Y(_09010_));
 sky130_fd_sc_hd__xnor2_1 _15916_ (.A(_09009_),
    .B(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__a22oi_2 _15917_ (.A1(\rbzero.wall_tracer.stepDistX[2] ),
    .A2(_08231_),
    .B1(_08304_),
    .B2(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_09012_));
 sky130_fd_sc_hd__and2_2 _15918_ (.A(_08320_),
    .B(_09012_),
    .X(_09013_));
 sky130_fd_sc_hd__a21oi_4 _15919_ (.A1(_08210_),
    .A2(_08326_),
    .B1(_08216_),
    .Y(_09014_));
 sky130_fd_sc_hd__inv_2 _15920_ (.A(_08102_),
    .Y(_09015_));
 sky130_fd_sc_hd__nor4_1 _15921_ (.A(_08084_),
    .B(_08090_),
    .C(_08097_),
    .D(_08217_),
    .Y(_09016_));
 sky130_fd_sc_hd__o41a_1 _15922_ (.A1(_08084_),
    .A2(_08090_),
    .A3(_08097_),
    .A4(_08217_),
    .B1(_08103_),
    .X(_09017_));
 sky130_fd_sc_hd__a211o_1 _15923_ (.A1(_09015_),
    .A2(_09016_),
    .B1(_09017_),
    .C1(_08210_),
    .X(_09018_));
 sky130_fd_sc_hd__a22o_2 _15924_ (.A1(\rbzero.wall_tracer.stepDistY[4] ),
    .A2(_08304_),
    .B1(_09014_),
    .B2(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__or4b_1 _15925_ (.A(_08322_),
    .B(_08330_),
    .C(_08830_),
    .D_N(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__nand2_1 _15926_ (.A(_08131_),
    .B(_08321_),
    .Y(_09021_));
 sky130_fd_sc_hd__a2bb2o_1 _15927_ (.A1_N(_08330_),
    .A2_N(_09021_),
    .B1(_09019_),
    .B2(_08349_),
    .X(_09022_));
 sky130_fd_sc_hd__or4bb_1 _15928_ (.A(_08312_),
    .B(_09013_),
    .C_N(_09020_),
    .D_N(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__a2bb2o_1 _15929_ (.A1_N(_08941_),
    .A2_N(_09013_),
    .B1(_09020_),
    .B2(_09022_),
    .X(_09024_));
 sky130_fd_sc_hd__a21o_1 _15930_ (.A1(_08313_),
    .A2(_08332_),
    .B1(_08331_),
    .X(_09025_));
 sky130_fd_sc_hd__nand3_1 _15931_ (.A(_09023_),
    .B(_09024_),
    .C(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__a21o_1 _15932_ (.A1(_09023_),
    .A2(_09024_),
    .B1(_09025_),
    .X(_09027_));
 sky130_fd_sc_hd__nand3_1 _15933_ (.A(_09011_),
    .B(_09026_),
    .C(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__a21o_1 _15934_ (.A1(_09026_),
    .A2(_09027_),
    .B1(_09011_),
    .X(_09029_));
 sky130_fd_sc_hd__and2_1 _15935_ (.A(_08334_),
    .B(_08345_),
    .X(_09030_));
 sky130_fd_sc_hd__a21o_1 _15936_ (.A1(_08297_),
    .A2(_08346_),
    .B1(_09030_),
    .X(_09031_));
 sky130_fd_sc_hd__nand3_1 _15937_ (.A(_09028_),
    .B(_09029_),
    .C(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__a21o_1 _15938_ (.A1(_09028_),
    .A2(_09029_),
    .B1(_09031_),
    .X(_09033_));
 sky130_fd_sc_hd__and3_1 _15939_ (.A(_09005_),
    .B(_09032_),
    .C(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__a21oi_1 _15940_ (.A1(_09032_),
    .A2(_09033_),
    .B1(_09005_),
    .Y(_09035_));
 sky130_fd_sc_hd__or2_1 _15941_ (.A(_09034_),
    .B(_09035_),
    .X(_09036_));
 sky130_fd_sc_hd__nor2_1 _15942_ (.A(_08347_),
    .B(_08375_),
    .Y(_09037_));
 sky130_fd_sc_hd__a21oi_1 _15943_ (.A1(_08376_),
    .A2(_08446_),
    .B1(_09037_),
    .Y(_09038_));
 sky130_fd_sc_hd__xor2_1 _15944_ (.A(_09036_),
    .B(_09038_),
    .X(_09039_));
 sky130_fd_sc_hd__or2b_1 _15945_ (.A(_08584_),
    .B_N(_08582_),
    .X(_09040_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(_09040_),
    .B(_08586_),
    .Y(_09041_));
 sky130_fd_sc_hd__or2_1 _15947_ (.A(_08435_),
    .B(_08444_),
    .X(_09042_));
 sky130_fd_sc_hd__or2b_1 _15948_ (.A(_08445_),
    .B_N(_08434_),
    .X(_09043_));
 sky130_fd_sc_hd__o22ai_1 _15949_ (.A1(_08494_),
    .A2(_08959_),
    .B1(_08567_),
    .B2(_08510_),
    .Y(_09044_));
 sky130_fd_sc_hd__or4_1 _15950_ (.A(_08494_),
    .B(_08506_),
    .C(_08678_),
    .D(_08520_),
    .X(_09045_));
 sky130_fd_sc_hd__nand2_1 _15951_ (.A(_09044_),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__or3_1 _15952_ (.A(_08509_),
    .B(_08573_),
    .C(_09046_),
    .X(_09047_));
 sky130_fd_sc_hd__o21ai_1 _15953_ (.A1(_08509_),
    .A2(_08573_),
    .B1(_09046_),
    .Y(_09048_));
 sky130_fd_sc_hd__and2_1 _15954_ (.A(_09047_),
    .B(_09048_),
    .X(_09049_));
 sky130_fd_sc_hd__or3_1 _15955_ (.A(_08529_),
    .B(_08551_),
    .C(_08580_),
    .X(_09050_));
 sky130_fd_sc_hd__nor2_1 _15956_ (.A(_08387_),
    .B(_08547_),
    .Y(_09051_));
 sky130_fd_sc_hd__xnor2_1 _15957_ (.A(_08577_),
    .B(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__nor2_1 _15958_ (.A(_08478_),
    .B(_08517_),
    .Y(_09053_));
 sky130_fd_sc_hd__xnor2_1 _15959_ (.A(_09052_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__a21oi_1 _15960_ (.A1(_08578_),
    .A2(_09050_),
    .B1(_09054_),
    .Y(_09055_));
 sky130_fd_sc_hd__and3_1 _15961_ (.A(_08578_),
    .B(_09050_),
    .C(_09054_),
    .X(_09056_));
 sky130_fd_sc_hd__nor2_1 _15962_ (.A(_09055_),
    .B(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__xnor2_1 _15963_ (.A(_09049_),
    .B(_09057_),
    .Y(_09058_));
 sky130_fd_sc_hd__a21o_1 _15964_ (.A1(_09042_),
    .A2(_09043_),
    .B1(_09058_),
    .X(_09059_));
 sky130_fd_sc_hd__nand3_1 _15965_ (.A(_09042_),
    .B(_09043_),
    .C(_09058_),
    .Y(_09060_));
 sky130_fd_sc_hd__nand2_1 _15966_ (.A(_09059_),
    .B(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__xnor2_1 _15967_ (.A(_09041_),
    .B(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__xnor2_1 _15968_ (.A(_09039_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__a21oi_1 _15969_ (.A1(_08492_),
    .A2(_08592_),
    .B1(_08490_),
    .Y(_09064_));
 sky130_fd_sc_hd__nor2_1 _15970_ (.A(_09063_),
    .B(_09064_),
    .Y(_09065_));
 sky130_fd_sc_hd__and2_1 _15971_ (.A(_09063_),
    .B(_09064_),
    .X(_09066_));
 sky130_fd_sc_hd__nor2_1 _15972_ (.A(_09065_),
    .B(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__or2b_1 _15973_ (.A(_08591_),
    .B_N(_08565_),
    .X(_09068_));
 sky130_fd_sc_hd__nand2_2 _15974_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08493_),
    .Y(_09069_));
 sky130_fd_sc_hd__clkbuf_4 _15975_ (.A(_09069_),
    .X(_09070_));
 sky130_fd_sc_hd__or2_1 _15976_ (.A(_08511_),
    .B(_09070_),
    .X(_09071_));
 sky130_fd_sc_hd__clkbuf_4 _15977_ (.A(_08573_),
    .X(_09072_));
 sky130_fd_sc_hd__o31a_1 _15978_ (.A1(_08511_),
    .A2(_08571_),
    .A3(_09072_),
    .B1(_08570_),
    .X(_09073_));
 sky130_fd_sc_hd__nor2_1 _15979_ (.A(_09071_),
    .B(_09073_),
    .Y(_09074_));
 sky130_fd_sc_hd__and2_1 _15980_ (.A(_09071_),
    .B(_09073_),
    .X(_09075_));
 sky130_fd_sc_hd__or2_1 _15981_ (.A(_09074_),
    .B(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__a21oi_2 _15982_ (.A1(_08589_),
    .A2(_09068_),
    .B1(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__and3_1 _15983_ (.A(_08589_),
    .B(_09068_),
    .C(_09076_),
    .X(_09078_));
 sky130_fd_sc_hd__nor2_1 _15984_ (.A(_09077_),
    .B(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__xnor2_2 _15985_ (.A(_09067_),
    .B(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__a2bb2o_1 _15986_ (.A1_N(_08593_),
    .A2_N(_08646_),
    .B1(_08647_),
    .B2(_08651_),
    .X(_09081_));
 sky130_fd_sc_hd__xnor2_2 _15987_ (.A(_09080_),
    .B(_09081_),
    .Y(_09082_));
 sky130_fd_sc_hd__xnor2_4 _15988_ (.A(_08649_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__nor2_1 _15989_ (.A(_08990_),
    .B(_08713_),
    .Y(_09084_));
 sky130_fd_sc_hd__or2_2 _15990_ (.A(_08711_),
    .B(_09084_),
    .X(_09085_));
 sky130_fd_sc_hd__xnor2_4 _15991_ (.A(_09083_),
    .B(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__and2b_1 _15992_ (.A_N(_09083_),
    .B(_09084_),
    .X(_09087_));
 sky130_fd_sc_hd__a21o_2 _15993_ (.A1(_08993_),
    .A2(_09086_),
    .B1(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__a21o_1 _15994_ (.A1(_09049_),
    .A2(_09057_),
    .B1(_09055_),
    .X(_09089_));
 sky130_fd_sc_hd__or2b_1 _15995_ (.A(_09004_),
    .B_N(_08994_),
    .X(_09090_));
 sky130_fd_sc_hd__or2_1 _15996_ (.A(_08506_),
    .B(_08476_),
    .X(_09091_));
 sky130_fd_sc_hd__or2_1 _15997_ (.A(_06420_),
    .B(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__or2_1 _15998_ (.A(_08678_),
    .B(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__clkbuf_4 _15999_ (.A(_08476_),
    .X(_09094_));
 sky130_fd_sc_hd__o22ai_1 _16000_ (.A1(_08494_),
    .A2(_09094_),
    .B1(_08959_),
    .B2(_08510_),
    .Y(_09095_));
 sky130_fd_sc_hd__nand2_1 _16001_ (.A(_09093_),
    .B(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__nor2_1 _16002_ (.A(_08567_),
    .B(_09072_),
    .Y(_09097_));
 sky130_fd_sc_hd__xnor2_1 _16003_ (.A(_09096_),
    .B(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__nor2_2 _16004_ (.A(_08430_),
    .B(_08546_),
    .Y(_09099_));
 sky130_fd_sc_hd__o22a_1 _16005_ (.A1(_08430_),
    .A2(_08547_),
    .B1(_08546_),
    .B2(_08387_),
    .X(_09100_));
 sky130_fd_sc_hd__a21oi_1 _16006_ (.A1(_09051_),
    .A2(_09099_),
    .B1(_09100_),
    .Y(_09101_));
 sky130_fd_sc_hd__nor2_1 _16007_ (.A(_08417_),
    .B(_08551_),
    .Y(_09102_));
 sky130_fd_sc_hd__xnor2_1 _16008_ (.A(_09101_),
    .B(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__or3_1 _16009_ (.A(_08387_),
    .B(_08808_),
    .C(_08577_),
    .X(_09104_));
 sky130_fd_sc_hd__a21boi_1 _16010_ (.A1(_09052_),
    .A2(_09053_),
    .B1_N(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__nor2_1 _16011_ (.A(_09103_),
    .B(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__and2_1 _16012_ (.A(_09103_),
    .B(_09105_),
    .X(_09107_));
 sky130_fd_sc_hd__nor2_1 _16013_ (.A(_09106_),
    .B(_09107_),
    .Y(_09108_));
 sky130_fd_sc_hd__xnor2_1 _16014_ (.A(_09098_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__a21o_1 _16015_ (.A1(_09002_),
    .A2(_09090_),
    .B1(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__nand3_1 _16016_ (.A(_09002_),
    .B(_09090_),
    .C(_09109_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand2_1 _16017_ (.A(_09110_),
    .B(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__xnor2_1 _16018_ (.A(_09089_),
    .B(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__o21ai_1 _16019_ (.A1(_08436_),
    .A2(_08997_),
    .B1(_08999_),
    .Y(_09114_));
 sky130_fd_sc_hd__a21bo_1 _16020_ (.A1(_09008_),
    .A2(_09010_),
    .B1_N(_09006_),
    .X(_09115_));
 sky130_fd_sc_hd__or2_1 _16021_ (.A(_08409_),
    .B(_08243_),
    .X(_09116_));
 sky130_fd_sc_hd__or2_1 _16022_ (.A(_08997_),
    .B(_09116_),
    .X(_09117_));
 sky130_fd_sc_hd__o22ai_1 _16023_ (.A1(_08438_),
    .A2(_08244_),
    .B1(_08295_),
    .B2(_08409_),
    .Y(_09118_));
 sky130_fd_sc_hd__nand2_1 _16024_ (.A(_09117_),
    .B(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__nor2_1 _16025_ (.A(_08370_),
    .B(_08442_),
    .Y(_09120_));
 sky130_fd_sc_hd__xor2_1 _16026_ (.A(_09119_),
    .B(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__xnor2_1 _16027_ (.A(_09115_),
    .B(_09121_),
    .Y(_09122_));
 sky130_fd_sc_hd__xor2_1 _16028_ (.A(_09114_),
    .B(_09122_),
    .X(_09123_));
 sky130_fd_sc_hd__or2_1 _16029_ (.A(_08272_),
    .B(_08306_),
    .X(_09124_));
 sky130_fd_sc_hd__or3_1 _16030_ (.A(_08271_),
    .B(_09124_),
    .C(_09013_),
    .X(_09125_));
 sky130_fd_sc_hd__clkbuf_4 _16031_ (.A(_09013_),
    .X(_09126_));
 sky130_fd_sc_hd__o21ai_1 _16032_ (.A1(_08918_),
    .A2(_09126_),
    .B1(_09124_),
    .Y(_09127_));
 sky130_fd_sc_hd__nand2_1 _16033_ (.A(_09125_),
    .B(_09127_),
    .Y(_09128_));
 sky130_fd_sc_hd__nor2_1 _16034_ (.A(_08371_),
    .B(_09007_),
    .Y(_09129_));
 sky130_fd_sc_hd__xnor2_1 _16035_ (.A(_09128_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__a21boi_4 _16036_ (.A1(\rbzero.wall_tracer.stepDistX[3] ),
    .A2(_08629_),
    .B1_N(_08330_),
    .Y(_09131_));
 sky130_fd_sc_hd__nor2_1 _16037_ (.A(_08312_),
    .B(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__nand2_1 _16038_ (.A(_08355_),
    .B(_09019_),
    .Y(_09133_));
 sky130_fd_sc_hd__o21ai_1 _16039_ (.A1(_08103_),
    .A2(_08324_),
    .B1(_08106_),
    .Y(_09134_));
 sky130_fd_sc_hd__o31a_1 _16040_ (.A1(_08103_),
    .A2(_08106_),
    .A3(_08324_),
    .B1(_08214_),
    .X(_09135_));
 sky130_fd_sc_hd__a21oi_4 _16041_ (.A1(_09134_),
    .A2(_09135_),
    .B1(_08327_),
    .Y(_09136_));
 sky130_fd_sc_hd__and3_2 _16042_ (.A(_04494_),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .C(_08239_),
    .X(_09137_));
 sky130_fd_sc_hd__o211a_1 _16043_ (.A1(_09136_),
    .A2(_09137_),
    .B1(\rbzero.wall_tracer.visualWallDist[-11] ),
    .C1(_08493_),
    .X(_09138_));
 sky130_fd_sc_hd__xnor2_1 _16044_ (.A(_09133_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__xor2_1 _16045_ (.A(_09132_),
    .B(_09139_),
    .X(_09140_));
 sky130_fd_sc_hd__and2_1 _16046_ (.A(_09020_),
    .B(_09023_),
    .X(_09141_));
 sky130_fd_sc_hd__xnor2_1 _16047_ (.A(_09140_),
    .B(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__xnor2_1 _16048_ (.A(_09130_),
    .B(_09142_),
    .Y(_09143_));
 sky130_fd_sc_hd__and2_1 _16049_ (.A(_09026_),
    .B(_09028_),
    .X(_09144_));
 sky130_fd_sc_hd__xor2_1 _16050_ (.A(_09143_),
    .B(_09144_),
    .X(_09145_));
 sky130_fd_sc_hd__xnor2_1 _16051_ (.A(_09123_),
    .B(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__a21boi_1 _16052_ (.A1(_09005_),
    .A2(_09033_),
    .B1_N(_09032_),
    .Y(_09147_));
 sky130_fd_sc_hd__nor2_1 _16053_ (.A(_09146_),
    .B(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__and2_1 _16054_ (.A(_09146_),
    .B(_09147_),
    .X(_09149_));
 sky130_fd_sc_hd__nor2_1 _16055_ (.A(_09148_),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__xnor2_1 _16056_ (.A(_09113_),
    .B(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__nor2_1 _16057_ (.A(_09036_),
    .B(_09038_),
    .Y(_09152_));
 sky130_fd_sc_hd__a21oi_1 _16058_ (.A1(_09039_),
    .A2(_09062_),
    .B1(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__xor2_1 _16059_ (.A(_09151_),
    .B(_09153_),
    .X(_09154_));
 sky130_fd_sc_hd__or2b_1 _16060_ (.A(_09061_),
    .B_N(_09041_),
    .X(_09155_));
 sky130_fd_sc_hd__nand2_4 _16061_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08493_),
    .Y(_09156_));
 sky130_fd_sc_hd__or2_1 _16062_ (.A(_08505_),
    .B(_09156_),
    .X(_09157_));
 sky130_fd_sc_hd__nor2_1 _16063_ (.A(_09071_),
    .B(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__clkbuf_4 _16064_ (.A(_09156_),
    .X(_09159_));
 sky130_fd_sc_hd__nor2_1 _16065_ (.A(_08509_),
    .B(_09070_),
    .Y(_09160_));
 sky130_fd_sc_hd__o21ba_1 _16066_ (.A1(_08511_),
    .A2(_09159_),
    .B1_N(_09160_),
    .X(_09161_));
 sky130_fd_sc_hd__or2_1 _16067_ (.A(_09158_),
    .B(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__a21oi_1 _16068_ (.A1(_09045_),
    .A2(_09047_),
    .B1(_09162_),
    .Y(_09163_));
 sky130_fd_sc_hd__and3_1 _16069_ (.A(_09045_),
    .B(_09047_),
    .C(_09162_),
    .X(_09164_));
 sky130_fd_sc_hd__nor2_1 _16070_ (.A(_09163_),
    .B(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(_09074_),
    .B(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__or2_1 _16072_ (.A(_09074_),
    .B(_09165_),
    .X(_09167_));
 sky130_fd_sc_hd__nand2_1 _16073_ (.A(_09166_),
    .B(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__a21oi_2 _16074_ (.A1(_09059_),
    .A2(_09155_),
    .B1(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__and3_1 _16075_ (.A(_09059_),
    .B(_09155_),
    .C(_09168_),
    .X(_09170_));
 sky130_fd_sc_hd__nor2_1 _16076_ (.A(_09169_),
    .B(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__xnor2_1 _16077_ (.A(_09154_),
    .B(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__a21oi_1 _16078_ (.A1(_09067_),
    .A2(_09079_),
    .B1(_09065_),
    .Y(_09173_));
 sky130_fd_sc_hd__xor2_1 _16079_ (.A(_09172_),
    .B(_09173_),
    .X(_09174_));
 sky130_fd_sc_hd__xnor2_1 _16080_ (.A(_09077_),
    .B(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__or2b_1 _16081_ (.A(_09080_),
    .B_N(_09081_),
    .X(_09176_));
 sky130_fd_sc_hd__a21boi_1 _16082_ (.A1(_08649_),
    .A2(_09082_),
    .B1_N(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__xor2_1 _16083_ (.A(_09175_),
    .B(_09177_),
    .X(_09178_));
 sky130_fd_sc_hd__and2b_1 _16084_ (.A_N(_09083_),
    .B(_08711_),
    .X(_09179_));
 sky130_fd_sc_hd__nand2_1 _16085_ (.A(_09178_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__or2_1 _16086_ (.A(_09178_),
    .B(_09179_),
    .X(_09181_));
 sky130_fd_sc_hd__and2_2 _16087_ (.A(_09180_),
    .B(_09181_),
    .X(_09182_));
 sky130_fd_sc_hd__xnor2_4 _16088_ (.A(_09088_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__mux2_1 _16089_ (.A0(_08275_),
    .A1(_08284_),
    .S(_08206_),
    .X(_09184_));
 sky130_fd_sc_hd__xor2_1 _16090_ (.A(_09183_),
    .B(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__xnor2_4 _16091_ (.A(_08993_),
    .B(_09086_),
    .Y(_09186_));
 sky130_fd_sc_hd__and2b_1 _16092_ (.A_N(_04536_),
    .B(\rbzero.debug_overlay.playerY[-7] ),
    .X(_09187_));
 sky130_fd_sc_hd__a21oi_1 _16093_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_08206_),
    .B1(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__xor2_4 _16094_ (.A(_08985_),
    .B(_08987_),
    .X(_09189_));
 sky130_fd_sc_hd__mux2_1 _16095_ (.A0(\rbzero.debug_overlay.playerY[-9] ),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_04536_),
    .X(_09190_));
 sky130_fd_sc_hd__nand2_1 _16096_ (.A(_09189_),
    .B(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__mux2_1 _16097_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_04536_),
    .X(_09192_));
 sky130_fd_sc_hd__xor2_4 _16098_ (.A(_08988_),
    .B(_08992_),
    .X(_09193_));
 sky130_fd_sc_hd__nor2_1 _16099_ (.A(_09192_),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__nand2_1 _16100_ (.A(_09192_),
    .B(_09193_),
    .Y(_09195_));
 sky130_fd_sc_hd__o221a_1 _16101_ (.A1(_09186_),
    .A2(_09188_),
    .B1(_09191_),
    .B2(_09194_),
    .C1(_09195_),
    .X(_09196_));
 sky130_fd_sc_hd__a21oi_1 _16102_ (.A1(_09186_),
    .A2(_09188_),
    .B1(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__xnor2_1 _16103_ (.A(_09185_),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__buf_4 _16104_ (.A(_08285_),
    .X(_09199_));
 sky130_fd_sc_hd__clkbuf_4 _16105_ (.A(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__mux2_1 _16106_ (.A0(_09200_),
    .A1(_06137_),
    .S(_08206_),
    .X(_09201_));
 sky130_fd_sc_hd__buf_2 _16107_ (.A(_09201_),
    .X(_09202_));
 sky130_fd_sc_hd__and2_1 _16108_ (.A(_09198_),
    .B(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__nor2_1 _16109_ (.A(_09198_),
    .B(_09202_),
    .Y(_09204_));
 sky130_fd_sc_hd__or3_1 _16110_ (.A(_08214_),
    .B(_09203_),
    .C(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__o211a_1 _16111_ (.A1(\rbzero.texu_hot[0] ),
    .A2(_08211_),
    .B1(_09205_),
    .C1(_04500_),
    .X(_00466_));
 sky130_fd_sc_hd__a21bo_2 _16112_ (.A1(_09088_),
    .A2(_09182_),
    .B1_N(_09180_),
    .X(_09206_));
 sky130_fd_sc_hd__or2_2 _16113_ (.A(_09175_),
    .B(_09177_),
    .X(_09207_));
 sky130_fd_sc_hd__or2b_1 _16114_ (.A(_09112_),
    .B_N(_09089_),
    .X(_09208_));
 sky130_fd_sc_hd__or3_1 _16115_ (.A(_08567_),
    .B(_08573_),
    .C(_09096_),
    .X(_09209_));
 sky130_fd_sc_hd__nor2_1 _16116_ (.A(_08520_),
    .B(_09069_),
    .Y(_09210_));
 sky130_fd_sc_hd__xnor2_1 _16117_ (.A(_09157_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand2_4 _16118_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08496_),
    .Y(_09212_));
 sky130_fd_sc_hd__buf_4 _16119_ (.A(_09212_),
    .X(_09213_));
 sky130_fd_sc_hd__nor2_1 _16120_ (.A(_08500_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__xnor2_1 _16121_ (.A(_09211_),
    .B(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__and3_1 _16122_ (.A(_09093_),
    .B(_09209_),
    .C(_09215_),
    .X(_09216_));
 sky130_fd_sc_hd__a21oi_2 _16123_ (.A1(_09093_),
    .A2(_09209_),
    .B1(_09215_),
    .Y(_09217_));
 sky130_fd_sc_hd__nor4_1 _16124_ (.A(_09158_),
    .B(_09163_),
    .C(_09216_),
    .D(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__o22a_1 _16125_ (.A1(_09158_),
    .A2(_09163_),
    .B1(_09216_),
    .B2(_09217_),
    .X(_09219_));
 sky130_fd_sc_hd__nor2_1 _16126_ (.A(_09218_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__a21oi_1 _16127_ (.A1(_09110_),
    .A2(_09208_),
    .B1(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__and3_1 _16128_ (.A(_09110_),
    .B(_09208_),
    .C(_09220_),
    .X(_09222_));
 sky130_fd_sc_hd__nor2_1 _16129_ (.A(_09221_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__xnor2_1 _16130_ (.A(_09166_),
    .B(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__a21o_1 _16131_ (.A1(_09098_),
    .A2(_09108_),
    .B1(_09106_),
    .X(_09225_));
 sky130_fd_sc_hd__or2b_1 _16132_ (.A(_09121_),
    .B_N(_09115_),
    .X(_09226_));
 sky130_fd_sc_hd__nand2_1 _16133_ (.A(_09114_),
    .B(_09122_),
    .Y(_09227_));
 sky130_fd_sc_hd__clkbuf_4 _16134_ (.A(_08831_),
    .X(_09228_));
 sky130_fd_sc_hd__o21ai_1 _16135_ (.A1(_08495_),
    .A2(_08831_),
    .B1(_09091_),
    .Y(_09229_));
 sky130_fd_sc_hd__o21ai_1 _16136_ (.A1(_09228_),
    .A2(_09092_),
    .B1(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__nor2_1 _16137_ (.A(_08959_),
    .B(_08573_),
    .Y(_09231_));
 sky130_fd_sc_hd__xnor2_1 _16138_ (.A(_09230_),
    .B(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__nor2_1 _16139_ (.A(_08370_),
    .B(_08547_),
    .Y(_09233_));
 sky130_fd_sc_hd__xnor2_1 _16140_ (.A(_09099_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__nor2_1 _16141_ (.A(_08387_),
    .B(_08551_),
    .Y(_09235_));
 sky130_fd_sc_hd__xnor2_1 _16142_ (.A(_09234_),
    .B(_09235_),
    .Y(_09236_));
 sky130_fd_sc_hd__a22oi_2 _16143_ (.A1(_09051_),
    .A2(_09099_),
    .B1(_09101_),
    .B2(_09102_),
    .Y(_09237_));
 sky130_fd_sc_hd__xnor2_1 _16144_ (.A(_09236_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__xnor2_1 _16145_ (.A(_09232_),
    .B(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__a21o_1 _16146_ (.A1(_09226_),
    .A2(_09227_),
    .B1(_09239_),
    .X(_09240_));
 sky130_fd_sc_hd__nand3_1 _16147_ (.A(_09226_),
    .B(_09227_),
    .C(_09239_),
    .Y(_09241_));
 sky130_fd_sc_hd__nand2_1 _16148_ (.A(_09240_),
    .B(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__xnor2_1 _16149_ (.A(_09225_),
    .B(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__a21bo_1 _16150_ (.A1(_09118_),
    .A2(_09120_),
    .B1_N(_09117_),
    .X(_09244_));
 sky130_fd_sc_hd__o31ai_2 _16151_ (.A1(_08371_),
    .A2(_09007_),
    .A3(_09128_),
    .B1(_09125_),
    .Y(_09245_));
 sky130_fd_sc_hd__or3_1 _16152_ (.A(_08396_),
    .B(_08233_),
    .C(_09116_),
    .X(_09246_));
 sky130_fd_sc_hd__o21ai_1 _16153_ (.A1(_08438_),
    .A2(_09007_),
    .B1(_09116_),
    .Y(_09247_));
 sky130_fd_sc_hd__and2_1 _16154_ (.A(_09246_),
    .B(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__nor2_1 _16155_ (.A(_08442_),
    .B(_08295_),
    .Y(_09249_));
 sky130_fd_sc_hd__xor2_1 _16156_ (.A(_09248_),
    .B(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__xnor2_1 _16157_ (.A(_09245_),
    .B(_09250_),
    .Y(_09251_));
 sky130_fd_sc_hd__xnor2_1 _16158_ (.A(_09244_),
    .B(_09251_),
    .Y(_09252_));
 sky130_fd_sc_hd__nor2_1 _16159_ (.A(_08371_),
    .B(_08307_),
    .Y(_09253_));
 sky130_fd_sc_hd__nor2_1 _16160_ (.A(_08918_),
    .B(_09126_),
    .Y(_09254_));
 sky130_fd_sc_hd__nor2_2 _16161_ (.A(_08272_),
    .B(_09131_),
    .Y(_09255_));
 sky130_fd_sc_hd__o22a_1 _16162_ (.A1(_08362_),
    .A2(_09013_),
    .B1(_09131_),
    .B2(_08918_),
    .X(_09256_));
 sky130_fd_sc_hd__a21oi_2 _16163_ (.A1(_09254_),
    .A2(_09255_),
    .B1(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__xor2_2 _16164_ (.A(_09253_),
    .B(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__and2_1 _16165_ (.A(\rbzero.wall_tracer.stepDistX[4] ),
    .B(_08231_),
    .X(_09259_));
 sky130_fd_sc_hd__a21oi_2 _16166_ (.A1(_06340_),
    .A2(_09019_),
    .B1(_09259_),
    .Y(_09260_));
 sky130_fd_sc_hd__nor2_1 _16167_ (.A(_08312_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__nand2_1 _16168_ (.A(\rbzero.wall_tracer.stepDistY[6] ),
    .B(_08304_),
    .Y(_09262_));
 sky130_fd_sc_hd__o31a_1 _16169_ (.A1(_08103_),
    .A2(_08106_),
    .A3(_08324_),
    .B1(_08110_),
    .X(_09263_));
 sky130_fd_sc_hd__or2_1 _16170_ (.A(_08106_),
    .B(_08110_),
    .X(_09264_));
 sky130_fd_sc_hd__nor3_1 _16171_ (.A(_08103_),
    .B(_08324_),
    .C(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__o31ai_4 _16172_ (.A1(_08210_),
    .A2(_09263_),
    .A3(_09265_),
    .B1(_09014_),
    .Y(_09266_));
 sky130_fd_sc_hd__nand2_1 _16173_ (.A(_09262_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__or3_1 _16174_ (.A(_08341_),
    .B(_08298_),
    .C(_09266_),
    .X(_09268_));
 sky130_fd_sc_hd__o211ai_2 _16175_ (.A1(_09136_),
    .A2(_09137_),
    .B1(_08131_),
    .C1(_08493_),
    .Y(_09269_));
 sky130_fd_sc_hd__a32oi_4 _16176_ (.A1(_08355_),
    .A2(_09138_),
    .A3(_09267_),
    .B1(_09268_),
    .B2(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__xnor2_2 _16177_ (.A(_09261_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__and3_1 _16178_ (.A(_08355_),
    .B(_09019_),
    .C(_09138_),
    .X(_09272_));
 sky130_fd_sc_hd__a21oi_2 _16179_ (.A1(_09132_),
    .A2(_09139_),
    .B1(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__xor2_2 _16180_ (.A(_09271_),
    .B(_09273_),
    .X(_09274_));
 sky130_fd_sc_hd__xnor2_2 _16181_ (.A(_09258_),
    .B(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__and2b_1 _16182_ (.A_N(_09141_),
    .B(_09140_),
    .X(_09276_));
 sky130_fd_sc_hd__a21o_1 _16183_ (.A1(_09130_),
    .A2(_09142_),
    .B1(_09276_),
    .X(_09277_));
 sky130_fd_sc_hd__xnor2_1 _16184_ (.A(_09275_),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__xnor2_1 _16185_ (.A(_09252_),
    .B(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__nor2_1 _16186_ (.A(_09143_),
    .B(_09144_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21oi_1 _16187_ (.A1(_09123_),
    .A2(_09145_),
    .B1(_09280_),
    .Y(_09281_));
 sky130_fd_sc_hd__nor2_1 _16188_ (.A(_09279_),
    .B(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__and2_1 _16189_ (.A(_09279_),
    .B(_09281_),
    .X(_09283_));
 sky130_fd_sc_hd__nor2_1 _16190_ (.A(_09282_),
    .B(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__xnor2_1 _16191_ (.A(_09243_),
    .B(_09284_),
    .Y(_09285_));
 sky130_fd_sc_hd__a21oi_1 _16192_ (.A1(_09113_),
    .A2(_09150_),
    .B1(_09148_),
    .Y(_09286_));
 sky130_fd_sc_hd__nor2_1 _16193_ (.A(_09285_),
    .B(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__and2_1 _16194_ (.A(_09285_),
    .B(_09286_),
    .X(_09288_));
 sky130_fd_sc_hd__nor2_1 _16195_ (.A(_09287_),
    .B(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__xnor2_1 _16196_ (.A(_09224_),
    .B(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__nor2_1 _16197_ (.A(_09151_),
    .B(_09153_),
    .Y(_09291_));
 sky130_fd_sc_hd__a21oi_1 _16198_ (.A1(_09154_),
    .A2(_09171_),
    .B1(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__nor2_1 _16199_ (.A(_09290_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__and2_1 _16200_ (.A(_09290_),
    .B(_09292_),
    .X(_09294_));
 sky130_fd_sc_hd__nor2_1 _16201_ (.A(_09293_),
    .B(_09294_),
    .Y(_09295_));
 sky130_fd_sc_hd__xnor2_2 _16202_ (.A(_09169_),
    .B(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__nor2_1 _16203_ (.A(_09172_),
    .B(_09173_),
    .Y(_09297_));
 sky130_fd_sc_hd__a21oi_2 _16204_ (.A1(_09077_),
    .A2(_09174_),
    .B1(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__xnor2_4 _16205_ (.A(_09296_),
    .B(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__xor2_4 _16206_ (.A(_09207_),
    .B(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__xnor2_4 _16207_ (.A(_09206_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__inv_2 _16208_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .Y(_09302_));
 sky130_fd_sc_hd__mux2_1 _16209_ (.A0(_09302_),
    .A1(_08388_),
    .S(_08206_),
    .X(_09303_));
 sky130_fd_sc_hd__xnor2_1 _16210_ (.A(_09301_),
    .B(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__nor2_1 _16211_ (.A(_09183_),
    .B(_09184_),
    .Y(_09305_));
 sky130_fd_sc_hd__a21oi_1 _16212_ (.A1(_09185_),
    .A2(_09197_),
    .B1(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__xnor2_1 _16213_ (.A(_09304_),
    .B(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__o21ai_1 _16214_ (.A1(_09202_),
    .A2(_09307_),
    .B1(_08211_),
    .Y(_09308_));
 sky130_fd_sc_hd__a21o_1 _16215_ (.A1(_09202_),
    .A2(_09307_),
    .B1(_09308_),
    .X(_09309_));
 sky130_fd_sc_hd__o211a_1 _16216_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_08211_),
    .B1(_09309_),
    .C1(_04500_),
    .X(_00467_));
 sky130_fd_sc_hd__or2_2 _16217_ (.A(_09296_),
    .B(_09298_),
    .X(_09310_));
 sky130_fd_sc_hd__a31o_1 _16218_ (.A1(_09074_),
    .A2(_09165_),
    .A3(_09223_),
    .B1(_09221_),
    .X(_09311_));
 sky130_fd_sc_hd__or2b_1 _16219_ (.A(_09242_),
    .B_N(_09225_),
    .X(_09312_));
 sky130_fd_sc_hd__nand2_4 _16220_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08493_),
    .Y(_09313_));
 sky130_fd_sc_hd__buf_4 _16221_ (.A(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__nor2_2 _16222_ (.A(_08511_),
    .B(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__nor2_1 _16223_ (.A(_08520_),
    .B(_09156_),
    .Y(_09316_));
 sky130_fd_sc_hd__nand2_1 _16224_ (.A(_09160_),
    .B(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__a21bo_1 _16225_ (.A1(_09211_),
    .A2(_09214_),
    .B1_N(_09317_),
    .X(_09318_));
 sky130_fd_sc_hd__nor2_1 _16226_ (.A(_08678_),
    .B(_09156_),
    .Y(_09319_));
 sky130_fd_sc_hd__nor2_1 _16227_ (.A(_08678_),
    .B(_09069_),
    .Y(_09320_));
 sky130_fd_sc_hd__nor2_1 _16228_ (.A(_09316_),
    .B(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__a21o_1 _16229_ (.A1(_09210_),
    .A2(_09319_),
    .B1(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__or3_1 _16230_ (.A(_08509_),
    .B(_09212_),
    .C(_09322_),
    .X(_09323_));
 sky130_fd_sc_hd__o21ai_1 _16231_ (.A1(_08509_),
    .A2(_09212_),
    .B1(_09322_),
    .Y(_09324_));
 sky130_fd_sc_hd__nand2_1 _16232_ (.A(_09323_),
    .B(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__a2bb2o_1 _16233_ (.A1_N(_08831_),
    .A2_N(_09092_),
    .B1(_09229_),
    .B2(_09231_),
    .X(_09326_));
 sky130_fd_sc_hd__and2b_1 _16234_ (.A_N(_09325_),
    .B(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__and2b_1 _16235_ (.A_N(_09326_),
    .B(_09325_),
    .X(_09328_));
 sky130_fd_sc_hd__nor2_1 _16236_ (.A(_09327_),
    .B(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__xnor2_1 _16237_ (.A(_09318_),
    .B(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__o21bai_1 _16238_ (.A1(_09158_),
    .A2(_09217_),
    .B1_N(_09216_),
    .Y(_09331_));
 sky130_fd_sc_hd__xor2_1 _16239_ (.A(_09330_),
    .B(_09331_),
    .X(_09332_));
 sky130_fd_sc_hd__nand2_1 _16240_ (.A(_09315_),
    .B(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__or2_1 _16241_ (.A(_09315_),
    .B(_09332_),
    .X(_09334_));
 sky130_fd_sc_hd__nand2_1 _16242_ (.A(_09333_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__a21oi_1 _16243_ (.A1(_09240_),
    .A2(_09312_),
    .B1(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand3_1 _16244_ (.A(_09240_),
    .B(_09312_),
    .C(_09335_),
    .Y(_09337_));
 sky130_fd_sc_hd__or2b_1 _16245_ (.A(_09336_),
    .B_N(_09337_),
    .X(_09338_));
 sky130_fd_sc_hd__nor3b_1 _16246_ (.A(_09216_),
    .B(_09217_),
    .C_N(_09163_),
    .Y(_09339_));
 sky130_fd_sc_hd__xnor2_1 _16247_ (.A(_09338_),
    .B(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__or2b_1 _16248_ (.A(_09237_),
    .B_N(_09236_),
    .X(_09341_));
 sky130_fd_sc_hd__a21bo_1 _16249_ (.A1(_09232_),
    .A2(_09238_),
    .B1_N(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__or2b_1 _16250_ (.A(_09251_),
    .B_N(_09244_),
    .X(_09343_));
 sky130_fd_sc_hd__a21bo_1 _16251_ (.A1(_09245_),
    .A2(_09250_),
    .B1_N(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__or4_1 _16252_ (.A(_06420_),
    .B(_08506_),
    .C(_08783_),
    .D(_08831_),
    .X(_09345_));
 sky130_fd_sc_hd__inv_2 _16253_ (.A(_09345_),
    .Y(_09346_));
 sky130_fd_sc_hd__buf_2 _16254_ (.A(_08783_),
    .X(_09347_));
 sky130_fd_sc_hd__o22a_1 _16255_ (.A1(_08495_),
    .A2(_09347_),
    .B1(_09228_),
    .B2(_08510_),
    .X(_09348_));
 sky130_fd_sc_hd__nor2_1 _16256_ (.A(_09346_),
    .B(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__nor2_1 _16257_ (.A(_09094_),
    .B(_09072_),
    .Y(_09350_));
 sky130_fd_sc_hd__xor2_2 _16258_ (.A(_09349_),
    .B(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__nor2_1 _16259_ (.A(_08546_),
    .B(_08295_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_1 _16260_ (.A(_09233_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__o22ai_1 _16261_ (.A1(_08370_),
    .A2(_08559_),
    .B1(_08295_),
    .B2(_08808_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_1 _16262_ (.A(_09353_),
    .B(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__or2_1 _16263_ (.A(_08430_),
    .B(_08551_),
    .X(_09356_));
 sky130_fd_sc_hd__xnor2_1 _16264_ (.A(_09355_),
    .B(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__clkbuf_4 _16265_ (.A(_08551_),
    .X(_09358_));
 sky130_fd_sc_hd__nand2_1 _16266_ (.A(_09099_),
    .B(_09233_),
    .Y(_09359_));
 sky130_fd_sc_hd__o31a_1 _16267_ (.A1(_08387_),
    .A2(_09358_),
    .A3(_09234_),
    .B1(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__nor2_1 _16268_ (.A(_09357_),
    .B(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__nand2_1 _16269_ (.A(_09357_),
    .B(_09360_),
    .Y(_09362_));
 sky130_fd_sc_hd__and2b_1 _16270_ (.A_N(_09361_),
    .B(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__xor2_1 _16271_ (.A(_09351_),
    .B(_09363_),
    .X(_09364_));
 sky130_fd_sc_hd__xnor2_1 _16272_ (.A(_09344_),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__xnor2_1 _16273_ (.A(_09342_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__a21bo_1 _16274_ (.A1(_09247_),
    .A2(_09249_),
    .B1_N(_09246_),
    .X(_09367_));
 sky130_fd_sc_hd__a22o_1 _16275_ (.A1(_09254_),
    .A2(_09255_),
    .B1(_09257_),
    .B2(_09253_),
    .X(_09368_));
 sky130_fd_sc_hd__or2_1 _16276_ (.A(_08409_),
    .B(_08306_),
    .X(_09369_));
 sky130_fd_sc_hd__or3_1 _16277_ (.A(_08438_),
    .B(_09007_),
    .C(_09369_),
    .X(_09370_));
 sky130_fd_sc_hd__clkbuf_4 _16278_ (.A(_08409_),
    .X(_09371_));
 sky130_fd_sc_hd__clkbuf_4 _16279_ (.A(_08438_),
    .X(_09372_));
 sky130_fd_sc_hd__o22ai_2 _16280_ (.A1(_09371_),
    .A2(_09007_),
    .B1(_08307_),
    .B2(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand2_1 _16281_ (.A(_09370_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__nor2_1 _16282_ (.A(_08442_),
    .B(_08244_),
    .Y(_09375_));
 sky130_fd_sc_hd__xnor2_2 _16283_ (.A(_09374_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__xor2_2 _16284_ (.A(_09368_),
    .B(_09376_),
    .X(_09377_));
 sky130_fd_sc_hd__xor2_2 _16285_ (.A(_09367_),
    .B(_09377_),
    .X(_09378_));
 sky130_fd_sc_hd__nor2_1 _16286_ (.A(_08371_),
    .B(_09126_),
    .Y(_09379_));
 sky130_fd_sc_hd__nor2_1 _16287_ (.A(_08271_),
    .B(_09260_),
    .Y(_09380_));
 sky130_fd_sc_hd__xnor2_1 _16288_ (.A(_09255_),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__xnor2_2 _16289_ (.A(_09379_),
    .B(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__o21ai_4 _16290_ (.A1(_09136_),
    .A2(_09137_),
    .B1(_06340_),
    .Y(_09383_));
 sky130_fd_sc_hd__nand2_4 _16291_ (.A(\rbzero.wall_tracer.stepDistX[5] ),
    .B(_08629_),
    .Y(_09384_));
 sky130_fd_sc_hd__a21oi_2 _16292_ (.A1(_09383_),
    .A2(_09384_),
    .B1(_08312_),
    .Y(_09385_));
 sky130_fd_sc_hd__or3_1 _16293_ (.A(_08314_),
    .B(_08298_),
    .C(_09266_),
    .X(_09386_));
 sky130_fd_sc_hd__nor4_1 _16294_ (.A(_08103_),
    .B(_08114_),
    .C(_08324_),
    .D(_09264_),
    .Y(_09387_));
 sky130_fd_sc_hd__o31a_1 _16295_ (.A1(_08103_),
    .A2(_08324_),
    .A3(_09264_),
    .B1(_08114_),
    .X(_09388_));
 sky130_fd_sc_hd__o31a_2 _16296_ (.A1(_08210_),
    .A2(_09387_),
    .A3(_09388_),
    .B1(_09014_),
    .X(_09389_));
 sky130_fd_sc_hd__and3_1 _16297_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08493_),
    .C(_09389_),
    .X(_09390_));
 sky130_fd_sc_hd__xnor2_2 _16298_ (.A(_09386_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__xor2_2 _16299_ (.A(_09385_),
    .B(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__and3_1 _16300_ (.A(_08355_),
    .B(_09138_),
    .C(_09267_),
    .X(_09393_));
 sky130_fd_sc_hd__a21o_1 _16301_ (.A1(_09261_),
    .A2(_09270_),
    .B1(_09393_),
    .X(_09394_));
 sky130_fd_sc_hd__xor2_2 _16302_ (.A(_09392_),
    .B(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__xnor2_2 _16303_ (.A(_09382_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__nor2_1 _16304_ (.A(_09271_),
    .B(_09273_),
    .Y(_09397_));
 sky130_fd_sc_hd__a21oi_2 _16305_ (.A1(_09258_),
    .A2(_09274_),
    .B1(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__xor2_2 _16306_ (.A(_09396_),
    .B(_09398_),
    .X(_09399_));
 sky130_fd_sc_hd__xnor2_2 _16307_ (.A(_09378_),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__and2b_1 _16308_ (.A_N(_09275_),
    .B(_09277_),
    .X(_09401_));
 sky130_fd_sc_hd__a21oi_1 _16309_ (.A1(_09252_),
    .A2(_09278_),
    .B1(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__nor2_1 _16310_ (.A(_09400_),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__and2_1 _16311_ (.A(_09400_),
    .B(_09402_),
    .X(_09404_));
 sky130_fd_sc_hd__nor2_1 _16312_ (.A(_09403_),
    .B(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__xnor2_1 _16313_ (.A(_09366_),
    .B(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__a21oi_1 _16314_ (.A1(_09243_),
    .A2(_09284_),
    .B1(_09282_),
    .Y(_09407_));
 sky130_fd_sc_hd__nor2_1 _16315_ (.A(_09406_),
    .B(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__and2_1 _16316_ (.A(_09406_),
    .B(_09407_),
    .X(_09409_));
 sky130_fd_sc_hd__nor2_1 _16317_ (.A(_09408_),
    .B(_09409_),
    .Y(_09410_));
 sky130_fd_sc_hd__xnor2_1 _16318_ (.A(_09340_),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__a21oi_1 _16319_ (.A1(_09224_),
    .A2(_09289_),
    .B1(_09287_),
    .Y(_09412_));
 sky130_fd_sc_hd__nor2_1 _16320_ (.A(_09411_),
    .B(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__and2_1 _16321_ (.A(_09411_),
    .B(_09412_),
    .X(_09414_));
 sky130_fd_sc_hd__nor2_1 _16322_ (.A(_09413_),
    .B(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__xnor2_2 _16323_ (.A(_09311_),
    .B(_09415_),
    .Y(_09416_));
 sky130_fd_sc_hd__a21oi_1 _16324_ (.A1(_09169_),
    .A2(_09295_),
    .B1(_09293_),
    .Y(_09417_));
 sky130_fd_sc_hd__xor2_2 _16325_ (.A(_09416_),
    .B(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__xor2_4 _16326_ (.A(_09310_),
    .B(_09418_),
    .X(_09419_));
 sky130_fd_sc_hd__a21oi_1 _16327_ (.A1(_09207_),
    .A2(_09180_),
    .B1(_09299_),
    .Y(_09420_));
 sky130_fd_sc_hd__a31oi_4 _16328_ (.A1(_09088_),
    .A2(_09182_),
    .A3(_09300_),
    .B1(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__xnor2_4 _16329_ (.A(_09419_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__inv_2 _16330_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_09423_));
 sky130_fd_sc_hd__mux2_1 _16331_ (.A0(_09423_),
    .A1(_08406_),
    .S(_08206_),
    .X(_09424_));
 sky130_fd_sc_hd__nor2_1 _16332_ (.A(_09422_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__nand2_1 _16333_ (.A(_09422_),
    .B(_09424_),
    .Y(_09426_));
 sky130_fd_sc_hd__or2b_1 _16334_ (.A(_09425_),
    .B_N(_09426_),
    .X(_09427_));
 sky130_fd_sc_hd__or2_1 _16335_ (.A(_09301_),
    .B(_09303_),
    .X(_09428_));
 sky130_fd_sc_hd__o21ai_1 _16336_ (.A1(_09304_),
    .A2(_09306_),
    .B1(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__xor2_1 _16337_ (.A(_09427_),
    .B(_09429_),
    .X(_09430_));
 sky130_fd_sc_hd__o21ai_1 _16338_ (.A1(_09202_),
    .A2(_09430_),
    .B1(_08211_),
    .Y(_09431_));
 sky130_fd_sc_hd__a21o_1 _16339_ (.A1(_09202_),
    .A2(_09430_),
    .B1(_09431_),
    .X(_09432_));
 sky130_fd_sc_hd__o211a_1 _16340_ (.A1(\rbzero.texu_hot[2] ),
    .A2(_08211_),
    .B1(_09432_),
    .C1(_04500_),
    .X(_00468_));
 sky130_fd_sc_hd__or2b_1 _16341_ (.A(_09310_),
    .B_N(_09418_),
    .X(_09433_));
 sky130_fd_sc_hd__o21ai_4 _16342_ (.A1(_09419_),
    .A2(_09421_),
    .B1(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__or2_2 _16343_ (.A(_09416_),
    .B(_09417_),
    .X(_09435_));
 sky130_fd_sc_hd__a21o_1 _16344_ (.A1(_09337_),
    .A2(_09339_),
    .B1(_09336_),
    .X(_09436_));
 sky130_fd_sc_hd__o21ai_1 _16345_ (.A1(_09330_),
    .A2(_09331_),
    .B1(_09333_),
    .Y(_09437_));
 sky130_fd_sc_hd__or2b_1 _16346_ (.A(_09365_),
    .B_N(_09342_),
    .X(_09438_));
 sky130_fd_sc_hd__a21bo_1 _16347_ (.A1(_09344_),
    .A2(_09364_),
    .B1_N(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__nand2_4 _16348_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08496_),
    .Y(_09440_));
 sky130_fd_sc_hd__clkbuf_4 _16349_ (.A(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__nor2_1 _16350_ (.A(_08509_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__nor2_1 _16351_ (.A(_08509_),
    .B(_09313_),
    .Y(_09443_));
 sky130_fd_sc_hd__o21ba_1 _16352_ (.A1(_08511_),
    .A2(_09441_),
    .B1_N(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__a21oi_1 _16353_ (.A1(_09315_),
    .A2(_09442_),
    .B1(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__a21bo_1 _16354_ (.A1(_09316_),
    .A2(_09320_),
    .B1_N(_09323_),
    .X(_09446_));
 sky130_fd_sc_hd__nor2_1 _16355_ (.A(_09094_),
    .B(_09070_),
    .Y(_09447_));
 sky130_fd_sc_hd__or2_1 _16356_ (.A(_09319_),
    .B(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__nand2_1 _16357_ (.A(_09319_),
    .B(_09447_),
    .Y(_09449_));
 sky130_fd_sc_hd__and2_1 _16358_ (.A(_09448_),
    .B(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__nor2_1 _16359_ (.A(_08567_),
    .B(_09213_),
    .Y(_09451_));
 sky130_fd_sc_hd__xnor2_1 _16360_ (.A(_09450_),
    .B(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__a21o_1 _16361_ (.A1(_09349_),
    .A2(_09350_),
    .B1(_09346_),
    .X(_09453_));
 sky130_fd_sc_hd__and2b_1 _16362_ (.A_N(_09452_),
    .B(_09453_),
    .X(_09454_));
 sky130_fd_sc_hd__and2b_1 _16363_ (.A_N(_09453_),
    .B(_09452_),
    .X(_09455_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__xnor2_1 _16365_ (.A(_09446_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__a21oi_1 _16366_ (.A1(_09318_),
    .A2(_09329_),
    .B1(_09327_),
    .Y(_09458_));
 sky130_fd_sc_hd__xor2_1 _16367_ (.A(_09457_),
    .B(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__xor2_1 _16368_ (.A(_09445_),
    .B(_09459_),
    .X(_09460_));
 sky130_fd_sc_hd__xnor2_1 _16369_ (.A(_09439_),
    .B(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__xnor2_1 _16370_ (.A(_09437_),
    .B(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__a21o_1 _16371_ (.A1(_09351_),
    .A2(_09362_),
    .B1(_09361_),
    .X(_09463_));
 sky130_fd_sc_hd__nand2_1 _16372_ (.A(_09368_),
    .B(_09376_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand2_1 _16373_ (.A(_09367_),
    .B(_09377_),
    .Y(_09465_));
 sky130_fd_sc_hd__clkbuf_4 _16374_ (.A(_08737_),
    .X(_09466_));
 sky130_fd_sc_hd__o22a_1 _16375_ (.A1(_08495_),
    .A2(_09466_),
    .B1(_08783_),
    .B2(_08510_),
    .X(_09467_));
 sky130_fd_sc_hd__or4_1 _16376_ (.A(_06420_),
    .B(_08510_),
    .C(_08737_),
    .D(_08783_),
    .X(_09468_));
 sky130_fd_sc_hd__or2b_1 _16377_ (.A(_09467_),
    .B_N(_09468_),
    .X(_09469_));
 sky130_fd_sc_hd__nor2_1 _16378_ (.A(_09228_),
    .B(_08573_),
    .Y(_09470_));
 sky130_fd_sc_hd__xnor2_1 _16379_ (.A(_09469_),
    .B(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__nor2_2 _16380_ (.A(_08547_),
    .B(_08244_),
    .Y(_09472_));
 sky130_fd_sc_hd__xnor2_1 _16381_ (.A(_09352_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__or2_1 _16382_ (.A(_08370_),
    .B(_08517_),
    .X(_09474_));
 sky130_fd_sc_hd__xnor2_1 _16383_ (.A(_09473_),
    .B(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__o31a_1 _16384_ (.A1(_08430_),
    .A2(_08551_),
    .A3(_09355_),
    .B1(_09353_),
    .X(_09476_));
 sky130_fd_sc_hd__xor2_1 _16385_ (.A(_09475_),
    .B(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__nand2_1 _16386_ (.A(_09471_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__or2_1 _16387_ (.A(_09471_),
    .B(_09477_),
    .X(_09479_));
 sky130_fd_sc_hd__nand2_1 _16388_ (.A(_09478_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__a21oi_2 _16389_ (.A1(_09464_),
    .A2(_09465_),
    .B1(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__and3_1 _16390_ (.A(_09464_),
    .B(_09465_),
    .C(_09480_),
    .X(_09482_));
 sky130_fd_sc_hd__nor2_1 _16391_ (.A(_09481_),
    .B(_09482_),
    .Y(_09483_));
 sky130_fd_sc_hd__xor2_1 _16392_ (.A(_09463_),
    .B(_09483_),
    .X(_09484_));
 sky130_fd_sc_hd__a21bo_1 _16393_ (.A1(_09373_),
    .A2(_09375_),
    .B1_N(_09370_),
    .X(_09485_));
 sky130_fd_sc_hd__nand2_1 _16394_ (.A(_09255_),
    .B(_09380_),
    .Y(_09486_));
 sky130_fd_sc_hd__o31a_1 _16395_ (.A1(_08371_),
    .A2(_09126_),
    .A3(_09381_),
    .B1(_09486_),
    .X(_09487_));
 sky130_fd_sc_hd__or3_1 _16396_ (.A(_08438_),
    .B(_09013_),
    .C(_09369_),
    .X(_09488_));
 sky130_fd_sc_hd__o21ai_1 _16397_ (.A1(_08438_),
    .A2(_09013_),
    .B1(_09369_),
    .Y(_09489_));
 sky130_fd_sc_hd__nand2_1 _16398_ (.A(_09488_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__or2_1 _16399_ (.A(_08429_),
    .B(_09007_),
    .X(_09491_));
 sky130_fd_sc_hd__xnor2_1 _16400_ (.A(_09490_),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__xor2_1 _16401_ (.A(_09487_),
    .B(_09492_),
    .X(_09493_));
 sky130_fd_sc_hd__xor2_1 _16402_ (.A(_09485_),
    .B(_09493_),
    .X(_09494_));
 sky130_fd_sc_hd__buf_2 _16403_ (.A(_09131_),
    .X(_09495_));
 sky130_fd_sc_hd__nor2_1 _16404_ (.A(_08371_),
    .B(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__buf_2 _16405_ (.A(_09260_),
    .X(_09497_));
 sky130_fd_sc_hd__nor2_1 _16406_ (.A(_08362_),
    .B(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__a21oi_1 _16407_ (.A1(_09383_),
    .A2(_09384_),
    .B1(_08918_),
    .Y(_09499_));
 sky130_fd_sc_hd__xor2_1 _16408_ (.A(_09498_),
    .B(_09499_),
    .X(_09500_));
 sky130_fd_sc_hd__xor2_1 _16409_ (.A(_09496_),
    .B(_09500_),
    .X(_09501_));
 sky130_fd_sc_hd__a21o_2 _16410_ (.A1(_09262_),
    .A2(_09266_),
    .B1(_08629_),
    .X(_09502_));
 sky130_fd_sc_hd__nand2_1 _16411_ (.A(\rbzero.wall_tracer.stepDistX[6] ),
    .B(_08629_),
    .Y(_09503_));
 sky130_fd_sc_hd__and2_1 _16412_ (.A(_09502_),
    .B(_09503_),
    .X(_09504_));
 sky130_fd_sc_hd__o41a_1 _16413_ (.A1(_08103_),
    .A2(_08114_),
    .A3(_08324_),
    .A4(_09264_),
    .B1(_08118_),
    .X(_09505_));
 sky130_fd_sc_hd__a211o_1 _16414_ (.A1(_08117_),
    .A2(_09387_),
    .B1(_09505_),
    .C1(_08210_),
    .X(_09506_));
 sky130_fd_sc_hd__a22oi_4 _16415_ (.A1(\rbzero.wall_tracer.stepDistY[8] ),
    .A2(_08304_),
    .B1(_09014_),
    .B2(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__and3_1 _16416_ (.A(_08131_),
    .B(_08234_),
    .C(_09389_),
    .X(_09508_));
 sky130_fd_sc_hd__or4b_1 _16417_ (.A(_08341_),
    .B(_08298_),
    .C(_09507_),
    .D_N(_09508_),
    .X(_09509_));
 sky130_fd_sc_hd__a22o_2 _16418_ (.A1(\rbzero.wall_tracer.stepDistY[8] ),
    .A2(_08304_),
    .B1(_09014_),
    .B2(_09506_),
    .X(_09510_));
 sky130_fd_sc_hd__a31o_1 _16419_ (.A1(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A2(_08496_),
    .A3(_09510_),
    .B1(_09508_),
    .X(_09511_));
 sky130_fd_sc_hd__or4bb_1 _16420_ (.A(_08941_),
    .B(_09504_),
    .C_N(_09509_),
    .D_N(_09511_),
    .X(_09512_));
 sky130_fd_sc_hd__a2bb2o_1 _16421_ (.A1_N(_08941_),
    .A2_N(_09504_),
    .B1(_09509_),
    .B2(_09511_),
    .X(_09513_));
 sky130_fd_sc_hd__and3_1 _16422_ (.A(_04494_),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .C(_08239_),
    .X(_09514_));
 sky130_fd_sc_hd__o21ai_4 _16423_ (.A1(_09514_),
    .A2(_09389_),
    .B1(_06340_),
    .Y(_09515_));
 sky130_fd_sc_hd__or3_1 _16424_ (.A(_08322_),
    .B(_09386_),
    .C(_09515_),
    .X(_09516_));
 sky130_fd_sc_hd__a21bo_1 _16425_ (.A1(_09385_),
    .A2(_09391_),
    .B1_N(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__nand3_1 _16426_ (.A(_09512_),
    .B(_09513_),
    .C(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__a21o_1 _16427_ (.A1(_09512_),
    .A2(_09513_),
    .B1(_09517_),
    .X(_09519_));
 sky130_fd_sc_hd__nand3_1 _16428_ (.A(_09501_),
    .B(_09518_),
    .C(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__a21o_1 _16429_ (.A1(_09518_),
    .A2(_09519_),
    .B1(_09501_),
    .X(_09521_));
 sky130_fd_sc_hd__and2_1 _16430_ (.A(_09392_),
    .B(_09394_),
    .X(_09522_));
 sky130_fd_sc_hd__a21o_1 _16431_ (.A1(_09382_),
    .A2(_09395_),
    .B1(_09522_),
    .X(_09523_));
 sky130_fd_sc_hd__nand3_1 _16432_ (.A(_09520_),
    .B(_09521_),
    .C(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__a21o_1 _16433_ (.A1(_09520_),
    .A2(_09521_),
    .B1(_09523_),
    .X(_09525_));
 sky130_fd_sc_hd__and3_1 _16434_ (.A(_09494_),
    .B(_09524_),
    .C(_09525_),
    .X(_09526_));
 sky130_fd_sc_hd__a21oi_1 _16435_ (.A1(_09524_),
    .A2(_09525_),
    .B1(_09494_),
    .Y(_09527_));
 sky130_fd_sc_hd__or2_1 _16436_ (.A(_09526_),
    .B(_09527_),
    .X(_09528_));
 sky130_fd_sc_hd__nor2_1 _16437_ (.A(_09396_),
    .B(_09398_),
    .Y(_09529_));
 sky130_fd_sc_hd__a21oi_1 _16438_ (.A1(_09378_),
    .A2(_09399_),
    .B1(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__xor2_1 _16439_ (.A(_09528_),
    .B(_09530_),
    .X(_09531_));
 sky130_fd_sc_hd__nand2_1 _16440_ (.A(_09484_),
    .B(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__or2_1 _16441_ (.A(_09484_),
    .B(_09531_),
    .X(_09533_));
 sky130_fd_sc_hd__nand2_1 _16442_ (.A(_09532_),
    .B(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__a21oi_1 _16443_ (.A1(_09366_),
    .A2(_09405_),
    .B1(_09403_),
    .Y(_09535_));
 sky130_fd_sc_hd__nor2_1 _16444_ (.A(_09534_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__and2_1 _16445_ (.A(_09534_),
    .B(_09535_),
    .X(_09537_));
 sky130_fd_sc_hd__nor2_1 _16446_ (.A(_09536_),
    .B(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__xnor2_1 _16447_ (.A(_09462_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__a21oi_1 _16448_ (.A1(_09340_),
    .A2(_09410_),
    .B1(_09408_),
    .Y(_09540_));
 sky130_fd_sc_hd__xnor2_1 _16449_ (.A(_09539_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__xor2_2 _16450_ (.A(_09436_),
    .B(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__a21oi_2 _16451_ (.A1(_09311_),
    .A2(_09415_),
    .B1(_09413_),
    .Y(_09543_));
 sky130_fd_sc_hd__xnor2_2 _16452_ (.A(_09542_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__xor2_4 _16453_ (.A(_09435_),
    .B(_09544_),
    .X(_09545_));
 sky130_fd_sc_hd__xnor2_4 _16454_ (.A(_09434_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__mux2_1 _16455_ (.A0(_04752_),
    .A1(_04749_),
    .S(_08206_),
    .X(_09547_));
 sky130_fd_sc_hd__nor2_1 _16456_ (.A(_09546_),
    .B(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__and2_1 _16457_ (.A(_09546_),
    .B(_09547_),
    .X(_09549_));
 sky130_fd_sc_hd__or2_1 _16458_ (.A(_09548_),
    .B(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__a21oi_1 _16459_ (.A1(_09426_),
    .A2(_09429_),
    .B1(_09425_),
    .Y(_09551_));
 sky130_fd_sc_hd__nor2_1 _16460_ (.A(_09550_),
    .B(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__and2_1 _16461_ (.A(_09550_),
    .B(_09551_),
    .X(_09553_));
 sky130_fd_sc_hd__or2_1 _16462_ (.A(_09552_),
    .B(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__o21ai_1 _16463_ (.A1(_09202_),
    .A2(_09554_),
    .B1(_08211_),
    .Y(_09555_));
 sky130_fd_sc_hd__a21o_1 _16464_ (.A1(_09202_),
    .A2(_09554_),
    .B1(_09555_),
    .X(_09556_));
 sky130_fd_sc_hd__o211a_1 _16465_ (.A1(\rbzero.texu_hot[3] ),
    .A2(_08211_),
    .B1(_09556_),
    .C1(_04500_),
    .X(_00469_));
 sky130_fd_sc_hd__nor2_1 _16466_ (.A(_09548_),
    .B(_09552_),
    .Y(_09557_));
 sky130_fd_sc_hd__inv_2 _16467_ (.A(_09545_),
    .Y(_09558_));
 sky130_fd_sc_hd__a21o_1 _16468_ (.A1(_09435_),
    .A2(_09433_),
    .B1(_09544_),
    .X(_09559_));
 sky130_fd_sc_hd__o31a_2 _16469_ (.A1(_09419_),
    .A2(_09421_),
    .A3(_09558_),
    .B1(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__nor2_1 _16470_ (.A(_09542_),
    .B(_09543_),
    .Y(_09561_));
 sky130_fd_sc_hd__or2b_1 _16471_ (.A(_09541_),
    .B_N(_09436_),
    .X(_09562_));
 sky130_fd_sc_hd__o21ai_1 _16472_ (.A1(_09539_),
    .A2(_09540_),
    .B1(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__or2b_1 _16473_ (.A(_09461_),
    .B_N(_09437_),
    .X(_09564_));
 sky130_fd_sc_hd__a21bo_1 _16474_ (.A1(_09439_),
    .A2(_09460_),
    .B1_N(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__a2bb2o_1 _16475_ (.A1_N(_09457_),
    .A2_N(_09458_),
    .B1(_09459_),
    .B2(_09445_),
    .X(_09566_));
 sky130_fd_sc_hd__and2_1 _16476_ (.A(_09463_),
    .B(_09483_),
    .X(_09567_));
 sky130_fd_sc_hd__nor2_1 _16477_ (.A(_08567_),
    .B(_09440_),
    .Y(_09568_));
 sky130_fd_sc_hd__o22a_1 _16478_ (.A1(_08567_),
    .A2(_09313_),
    .B1(_09441_),
    .B2(_08509_),
    .X(_09569_));
 sky130_fd_sc_hd__a21o_1 _16479_ (.A1(_09443_),
    .A2(_09568_),
    .B1(_09569_),
    .X(_09570_));
 sky130_fd_sc_hd__nand2_8 _16480_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_08496_),
    .Y(_09571_));
 sky130_fd_sc_hd__nor2_1 _16481_ (.A(_08511_),
    .B(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__xnor2_1 _16482_ (.A(_09570_),
    .B(_09572_),
    .Y(_09573_));
 sky130_fd_sc_hd__nand3_1 _16483_ (.A(_09315_),
    .B(_09442_),
    .C(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__a21o_1 _16484_ (.A1(_09315_),
    .A2(_09442_),
    .B1(_09573_),
    .X(_09575_));
 sky130_fd_sc_hd__nand2_1 _16485_ (.A(_09574_),
    .B(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__a21bo_1 _16486_ (.A1(_09450_),
    .A2(_09451_),
    .B1_N(_09449_),
    .X(_09577_));
 sky130_fd_sc_hd__nor2_1 _16487_ (.A(_08959_),
    .B(_09212_),
    .Y(_09578_));
 sky130_fd_sc_hd__nor2_1 _16488_ (.A(_08831_),
    .B(_09159_),
    .Y(_09579_));
 sky130_fd_sc_hd__o22a_1 _16489_ (.A1(_08831_),
    .A2(_09070_),
    .B1(_09159_),
    .B2(_09094_),
    .X(_09580_));
 sky130_fd_sc_hd__a21oi_1 _16490_ (.A1(_09447_),
    .A2(_09579_),
    .B1(_09580_),
    .Y(_09581_));
 sky130_fd_sc_hd__xnor2_1 _16491_ (.A(_09578_),
    .B(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__o31ai_1 _16492_ (.A1(_09228_),
    .A2(_09072_),
    .A3(_09467_),
    .B1(_09468_),
    .Y(_09583_));
 sky130_fd_sc_hd__and2b_1 _16493_ (.A_N(_09582_),
    .B(_09583_),
    .X(_09584_));
 sky130_fd_sc_hd__and2b_1 _16494_ (.A_N(_09583_),
    .B(_09582_),
    .X(_09585_));
 sky130_fd_sc_hd__nor2_1 _16495_ (.A(_09584_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__xnor2_2 _16496_ (.A(_09577_),
    .B(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__a21oi_2 _16497_ (.A1(_09446_),
    .A2(_09456_),
    .B1(_09454_),
    .Y(_09588_));
 sky130_fd_sc_hd__xor2_1 _16498_ (.A(_09587_),
    .B(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__xnor2_1 _16499_ (.A(_09576_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__o21a_1 _16500_ (.A1(_09481_),
    .A2(_09567_),
    .B1(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__nor3_1 _16501_ (.A(_09481_),
    .B(_09567_),
    .C(_09590_),
    .Y(_09592_));
 sky130_fd_sc_hd__nor2_1 _16502_ (.A(_09591_),
    .B(_09592_),
    .Y(_09593_));
 sky130_fd_sc_hd__xor2_1 _16503_ (.A(_09566_),
    .B(_09593_),
    .X(_09594_));
 sky130_fd_sc_hd__or2_1 _16504_ (.A(_09528_),
    .B(_09530_),
    .X(_09595_));
 sky130_fd_sc_hd__o21ai_1 _16505_ (.A1(_09475_),
    .A2(_09476_),
    .B1(_09478_),
    .Y(_09596_));
 sky130_fd_sc_hd__or2_1 _16506_ (.A(_09487_),
    .B(_09492_),
    .X(_09597_));
 sky130_fd_sc_hd__a21bo_1 _16507_ (.A1(_09485_),
    .A2(_09493_),
    .B1_N(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__o22ai_1 _16508_ (.A1(_08495_),
    .A2(_08661_),
    .B1(_09466_),
    .B2(_08510_),
    .Y(_09599_));
 sky130_fd_sc_hd__or4_1 _16509_ (.A(_08494_),
    .B(_08506_),
    .C(_08661_),
    .D(_08737_),
    .X(_09600_));
 sky130_fd_sc_hd__nand2_1 _16510_ (.A(_09599_),
    .B(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__or3_1 _16511_ (.A(_09347_),
    .B(_08573_),
    .C(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__o21ai_1 _16512_ (.A1(_09347_),
    .A2(_09072_),
    .B1(_09601_),
    .Y(_09603_));
 sky130_fd_sc_hd__and2_1 _16513_ (.A(_09602_),
    .B(_09603_),
    .X(_09604_));
 sky130_fd_sc_hd__nor2_2 _16514_ (.A(_08559_),
    .B(_09007_),
    .Y(_09605_));
 sky130_fd_sc_hd__o22a_1 _16515_ (.A1(_08808_),
    .A2(_09007_),
    .B1(_08244_),
    .B2(_08559_),
    .X(_09606_));
 sky130_fd_sc_hd__a21oi_1 _16516_ (.A1(_09472_),
    .A2(_09605_),
    .B1(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__nor2_1 _16517_ (.A(_08551_),
    .B(_08295_),
    .Y(_09608_));
 sky130_fd_sc_hd__xnor2_1 _16518_ (.A(_09607_),
    .B(_09608_),
    .Y(_09609_));
 sky130_fd_sc_hd__nand2_1 _16519_ (.A(_09352_),
    .B(_09472_),
    .Y(_09610_));
 sky130_fd_sc_hd__o31a_1 _16520_ (.A1(_08370_),
    .A2(_09358_),
    .A3(_09473_),
    .B1(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__nor2_1 _16521_ (.A(_09609_),
    .B(_09611_),
    .Y(_09612_));
 sky130_fd_sc_hd__and2_1 _16522_ (.A(_09609_),
    .B(_09611_),
    .X(_09613_));
 sky130_fd_sc_hd__nor2_1 _16523_ (.A(_09612_),
    .B(_09613_),
    .Y(_09614_));
 sky130_fd_sc_hd__xor2_1 _16524_ (.A(_09604_),
    .B(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__nand2_1 _16525_ (.A(_09598_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__or2_1 _16526_ (.A(_09598_),
    .B(_09615_),
    .X(_09617_));
 sky130_fd_sc_hd__nand2_1 _16527_ (.A(_09616_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__xnor2_1 _16528_ (.A(_09596_),
    .B(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__o21ai_1 _16529_ (.A1(_09490_),
    .A2(_09491_),
    .B1(_09488_),
    .Y(_09620_));
 sky130_fd_sc_hd__a22o_1 _16530_ (.A1(_09498_),
    .A2(_09499_),
    .B1(_09500_),
    .B2(_09496_),
    .X(_09621_));
 sky130_fd_sc_hd__nor2_1 _16531_ (.A(_09372_),
    .B(_09126_),
    .Y(_09622_));
 sky130_fd_sc_hd__nor2_1 _16532_ (.A(_09371_),
    .B(_09495_),
    .Y(_09623_));
 sky130_fd_sc_hd__o22a_1 _16533_ (.A1(_09371_),
    .A2(_09126_),
    .B1(_09495_),
    .B2(_09372_),
    .X(_09624_));
 sky130_fd_sc_hd__a21o_1 _16534_ (.A1(_09622_),
    .A2(_09623_),
    .B1(_09624_),
    .X(_09625_));
 sky130_fd_sc_hd__or2_1 _16535_ (.A(_08429_),
    .B(_08307_),
    .X(_09626_));
 sky130_fd_sc_hd__xor2_1 _16536_ (.A(_09625_),
    .B(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__xor2_1 _16537_ (.A(_09621_),
    .B(_09627_),
    .X(_09628_));
 sky130_fd_sc_hd__xor2_1 _16538_ (.A(_09620_),
    .B(_09628_),
    .X(_09629_));
 sky130_fd_sc_hd__clkbuf_4 _16539_ (.A(_09504_),
    .X(_09630_));
 sky130_fd_sc_hd__or3b_1 _16540_ (.A(_08362_),
    .B(_09630_),
    .C_N(_09499_),
    .X(_09631_));
 sky130_fd_sc_hd__and2_1 _16541_ (.A(_09383_),
    .B(_09384_),
    .X(_09632_));
 sky130_fd_sc_hd__buf_2 _16542_ (.A(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__o22ai_1 _16543_ (.A1(_08362_),
    .A2(_09633_),
    .B1(_09630_),
    .B2(_08918_),
    .Y(_09634_));
 sky130_fd_sc_hd__nand2_1 _16544_ (.A(_09631_),
    .B(_09634_),
    .Y(_09635_));
 sky130_fd_sc_hd__nor2_1 _16545_ (.A(_08371_),
    .B(_09497_),
    .Y(_09636_));
 sky130_fd_sc_hd__xnor2_1 _16546_ (.A(_09635_),
    .B(_09636_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand2_1 _16547_ (.A(\rbzero.wall_tracer.stepDistX[7] ),
    .B(_08629_),
    .Y(_09638_));
 sky130_fd_sc_hd__and2_1 _16548_ (.A(_09515_),
    .B(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__nor2_1 _16549_ (.A(_08941_),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__or4_1 _16550_ (.A(_08102_),
    .B(_08114_),
    .C(_08324_),
    .D(_09264_),
    .X(_09641_));
 sky130_fd_sc_hd__or3_1 _16551_ (.A(_08118_),
    .B(_08120_),
    .C(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__o21ai_1 _16552_ (.A1(_08118_),
    .A2(_09641_),
    .B1(_08120_),
    .Y(_09643_));
 sky130_fd_sc_hd__a31o_1 _16553_ (.A1(_08214_),
    .A2(_09642_),
    .A3(_09643_),
    .B1(_08327_),
    .X(_09644_));
 sky130_fd_sc_hd__or3_1 _16554_ (.A(_08341_),
    .B(_08298_),
    .C(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__nor2_1 _16555_ (.A(_08830_),
    .B(_09507_),
    .Y(_09646_));
 sky130_fd_sc_hd__xnor2_1 _16556_ (.A(_09645_),
    .B(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__xnor2_1 _16557_ (.A(_09640_),
    .B(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__and2_1 _16558_ (.A(_09509_),
    .B(_09512_),
    .X(_09649_));
 sky130_fd_sc_hd__xor2_1 _16559_ (.A(_09648_),
    .B(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__xnor2_1 _16560_ (.A(_09637_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__and2_1 _16561_ (.A(_09518_),
    .B(_09520_),
    .X(_09652_));
 sky130_fd_sc_hd__xor2_1 _16562_ (.A(_09651_),
    .B(_09652_),
    .X(_09653_));
 sky130_fd_sc_hd__xnor2_1 _16563_ (.A(_09629_),
    .B(_09653_),
    .Y(_09654_));
 sky130_fd_sc_hd__a21boi_1 _16564_ (.A1(_09494_),
    .A2(_09525_),
    .B1_N(_09524_),
    .Y(_09655_));
 sky130_fd_sc_hd__nor2_1 _16565_ (.A(_09654_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_1 _16566_ (.A(_09654_),
    .B(_09655_),
    .Y(_09657_));
 sky130_fd_sc_hd__and2b_1 _16567_ (.A_N(_09656_),
    .B(_09657_),
    .X(_09658_));
 sky130_fd_sc_hd__xnor2_1 _16568_ (.A(_09619_),
    .B(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__a21oi_1 _16569_ (.A1(_09595_),
    .A2(_09532_),
    .B1(_09659_),
    .Y(_09660_));
 sky130_fd_sc_hd__and3_1 _16570_ (.A(_09595_),
    .B(_09532_),
    .C(_09659_),
    .X(_09661_));
 sky130_fd_sc_hd__nor2_1 _16571_ (.A(_09660_),
    .B(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__xnor2_1 _16572_ (.A(_09594_),
    .B(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__a21oi_1 _16573_ (.A1(_09462_),
    .A2(_09538_),
    .B1(_09536_),
    .Y(_09664_));
 sky130_fd_sc_hd__nor2_1 _16574_ (.A(_09663_),
    .B(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__nand2_1 _16575_ (.A(_09663_),
    .B(_09664_),
    .Y(_09666_));
 sky130_fd_sc_hd__and2b_1 _16576_ (.A_N(_09665_),
    .B(_09666_),
    .X(_09667_));
 sky130_fd_sc_hd__xnor2_1 _16577_ (.A(_09565_),
    .B(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__xnor2_1 _16578_ (.A(_09563_),
    .B(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__nand2_1 _16579_ (.A(_09561_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__or2_1 _16580_ (.A(_09561_),
    .B(_09669_),
    .X(_09671_));
 sky130_fd_sc_hd__nand2_2 _16581_ (.A(_09670_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__xor2_4 _16582_ (.A(_09560_),
    .B(_09672_),
    .X(_09673_));
 sky130_fd_sc_hd__mux2_1 _16583_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_08206_),
    .X(_09674_));
 sky130_fd_sc_hd__nor2_1 _16584_ (.A(_09673_),
    .B(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__and2_1 _16585_ (.A(_09673_),
    .B(_09674_),
    .X(_09676_));
 sky130_fd_sc_hd__nor2_1 _16586_ (.A(_09675_),
    .B(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__xor2_1 _16587_ (.A(_09202_),
    .B(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__nor2_1 _16588_ (.A(_09557_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__a21o_1 _16589_ (.A1(_09557_),
    .A2(_09678_),
    .B1(_08214_),
    .X(_09680_));
 sky130_fd_sc_hd__or2_1 _16590_ (.A(\rbzero.texu_hot[4] ),
    .B(_08211_),
    .X(_09681_));
 sky130_fd_sc_hd__o211a_1 _16591_ (.A1(_09679_),
    .A2(_09680_),
    .B1(_09681_),
    .C1(_04500_),
    .X(_00470_));
 sky130_fd_sc_hd__inv_2 _16592_ (.A(_09675_),
    .Y(_09682_));
 sky130_fd_sc_hd__o31a_1 _16593_ (.A1(_09548_),
    .A2(_09552_),
    .A3(_09676_),
    .B1(_09682_),
    .X(_09683_));
 sky130_fd_sc_hd__o21a_1 _16594_ (.A1(_09560_),
    .A2(_09672_),
    .B1(_09670_),
    .X(_09684_));
 sky130_fd_sc_hd__or2b_2 _16595_ (.A(_09668_),
    .B_N(_09563_),
    .X(_09685_));
 sky130_fd_sc_hd__a21oi_1 _16596_ (.A1(_09566_),
    .A2(_09593_),
    .B1(_09591_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand2_4 _16597_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_08496_),
    .Y(_09687_));
 sky130_fd_sc_hd__or3_1 _16598_ (.A(_08630_),
    .B(_09686_),
    .C(_09687_),
    .X(_09688_));
 sky130_fd_sc_hd__or2_1 _16599_ (.A(_09574_),
    .B(_09686_),
    .X(_09689_));
 sky130_fd_sc_hd__nand2_1 _16600_ (.A(_09574_),
    .B(_09686_),
    .Y(_09690_));
 sky130_fd_sc_hd__nor2_4 _16601_ (.A(_06270_),
    .B(_08298_),
    .Y(_09691_));
 sky130_fd_sc_hd__a22o_1 _16602_ (.A1(_09689_),
    .A2(_09690_),
    .B1(_09691_),
    .B2(_08511_),
    .X(_09692_));
 sky130_fd_sc_hd__and2_2 _16603_ (.A(_09688_),
    .B(_09692_),
    .X(_09693_));
 sky130_fd_sc_hd__or2b_1 _16604_ (.A(_09576_),
    .B_N(_09589_),
    .X(_09694_));
 sky130_fd_sc_hd__o21ai_2 _16605_ (.A1(_09587_),
    .A2(_09588_),
    .B1(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__or2b_1 _16606_ (.A(_09618_),
    .B_N(_09596_),
    .X(_09696_));
 sky130_fd_sc_hd__nor2_1 _16607_ (.A(_09094_),
    .B(_09313_),
    .Y(_09697_));
 sky130_fd_sc_hd__o22a_1 _16608_ (.A1(_09094_),
    .A2(_09212_),
    .B1(_09313_),
    .B2(_08959_),
    .X(_09698_));
 sky130_fd_sc_hd__a21oi_1 _16609_ (.A1(_09578_),
    .A2(_09697_),
    .B1(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__and2_1 _16610_ (.A(_09568_),
    .B(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__nor2_1 _16611_ (.A(_09568_),
    .B(_09699_),
    .Y(_09701_));
 sky130_fd_sc_hd__or2_1 _16612_ (.A(_09700_),
    .B(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__nand2_1 _16613_ (.A(_09443_),
    .B(_09568_),
    .Y(_09703_));
 sky130_fd_sc_hd__o31a_1 _16614_ (.A1(_08511_),
    .A2(_09570_),
    .A3(_09571_),
    .B1(_09703_),
    .X(_09704_));
 sky130_fd_sc_hd__xor2_1 _16615_ (.A(_09702_),
    .B(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__buf_4 _16616_ (.A(_09571_),
    .X(_09706_));
 sky130_fd_sc_hd__nor2_1 _16617_ (.A(_08509_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__xor2_1 _16618_ (.A(_09705_),
    .B(_09707_),
    .X(_09708_));
 sky130_fd_sc_hd__nand2_1 _16619_ (.A(_09447_),
    .B(_09579_),
    .Y(_09709_));
 sky130_fd_sc_hd__a21bo_1 _16620_ (.A1(_09578_),
    .A2(_09581_),
    .B1_N(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__o22a_1 _16621_ (.A1(_08737_),
    .A2(_08573_),
    .B1(_09070_),
    .B2(_09347_),
    .X(_09711_));
 sky130_fd_sc_hd__or2_1 _16622_ (.A(_08737_),
    .B(_09069_),
    .X(_09712_));
 sky130_fd_sc_hd__or3_1 _16623_ (.A(_08783_),
    .B(_08572_),
    .C(_09712_),
    .X(_09713_));
 sky130_fd_sc_hd__and2b_1 _16624_ (.A_N(_09711_),
    .B(_09713_),
    .X(_09714_));
 sky130_fd_sc_hd__xnor2_1 _16625_ (.A(_09579_),
    .B(_09714_),
    .Y(_09715_));
 sky130_fd_sc_hd__a21oi_1 _16626_ (.A1(_09600_),
    .A2(_09602_),
    .B1(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__and3_1 _16627_ (.A(_09600_),
    .B(_09602_),
    .C(_09715_),
    .X(_09717_));
 sky130_fd_sc_hd__nor2_1 _16628_ (.A(_09716_),
    .B(_09717_),
    .Y(_09718_));
 sky130_fd_sc_hd__xnor2_1 _16629_ (.A(_09710_),
    .B(_09718_),
    .Y(_09719_));
 sky130_fd_sc_hd__a21oi_1 _16630_ (.A1(_09577_),
    .A2(_09586_),
    .B1(_09584_),
    .Y(_09720_));
 sky130_fd_sc_hd__nor2_1 _16631_ (.A(_09719_),
    .B(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__and2_1 _16632_ (.A(_09719_),
    .B(_09720_),
    .X(_09722_));
 sky130_fd_sc_hd__nor2_1 _16633_ (.A(_09721_),
    .B(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__xnor2_1 _16634_ (.A(_09708_),
    .B(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__a21o_1 _16635_ (.A1(_09616_),
    .A2(_09696_),
    .B1(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__nand3_1 _16636_ (.A(_09616_),
    .B(_09696_),
    .C(_09724_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand2_1 _16637_ (.A(_09725_),
    .B(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__xnor2_2 _16638_ (.A(_09695_),
    .B(_09727_),
    .Y(_09728_));
 sky130_fd_sc_hd__a21o_1 _16639_ (.A1(_09604_),
    .A2(_09614_),
    .B1(_09612_),
    .X(_09729_));
 sky130_fd_sc_hd__nand2_1 _16640_ (.A(_09621_),
    .B(_09627_),
    .Y(_09730_));
 sky130_fd_sc_hd__a21bo_1 _16641_ (.A1(_09620_),
    .A2(_09628_),
    .B1_N(_09730_),
    .X(_09731_));
 sky130_fd_sc_hd__nor2_1 _16642_ (.A(_08510_),
    .B(_08661_),
    .Y(_09732_));
 sky130_fd_sc_hd__nor2_1 _16643_ (.A(_08517_),
    .B(_08244_),
    .Y(_09733_));
 sky130_fd_sc_hd__nor2_1 _16644_ (.A(_08494_),
    .B(_08293_),
    .Y(_09734_));
 sky130_fd_sc_hd__xor2_1 _16645_ (.A(_09733_),
    .B(_09734_),
    .X(_09735_));
 sky130_fd_sc_hd__xor2_1 _16646_ (.A(_09732_),
    .B(_09735_),
    .X(_09736_));
 sky130_fd_sc_hd__a21o_1 _16647_ (.A1(_08336_),
    .A2(_09012_),
    .B1(_08547_),
    .X(_09737_));
 sky130_fd_sc_hd__nor2_1 _16648_ (.A(_09626_),
    .B(_09737_),
    .Y(_09738_));
 sky130_fd_sc_hd__or2_1 _16649_ (.A(_08808_),
    .B(_08307_),
    .X(_09739_));
 sky130_fd_sc_hd__o21ai_1 _16650_ (.A1(_08442_),
    .A2(_09126_),
    .B1(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__and2b_1 _16651_ (.A_N(_09738_),
    .B(_09740_),
    .X(_09741_));
 sky130_fd_sc_hd__xnor2_1 _16652_ (.A(_09605_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__a22oi_2 _16653_ (.A1(_09472_),
    .A2(_09605_),
    .B1(_09607_),
    .B2(_09608_),
    .Y(_09743_));
 sky130_fd_sc_hd__nor2_1 _16654_ (.A(_09742_),
    .B(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__nand2_1 _16655_ (.A(_09742_),
    .B(_09743_),
    .Y(_09745_));
 sky130_fd_sc_hd__and2b_1 _16656_ (.A_N(_09744_),
    .B(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__xnor2_1 _16657_ (.A(_09736_),
    .B(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__xor2_1 _16658_ (.A(_09731_),
    .B(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__xnor2_2 _16659_ (.A(_09729_),
    .B(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__a2bb2o_1 _16660_ (.A1_N(_09624_),
    .A2_N(_09626_),
    .B1(_09622_),
    .B2(_09623_),
    .X(_09750_));
 sky130_fd_sc_hd__clkbuf_4 _16661_ (.A(_08371_),
    .X(_09751_));
 sky130_fd_sc_hd__o31a_1 _16662_ (.A1(_09751_),
    .A2(_09497_),
    .A3(_09635_),
    .B1(_09631_),
    .X(_09752_));
 sky130_fd_sc_hd__a21oi_2 _16663_ (.A1(_09383_),
    .A2(_09384_),
    .B1(_08438_),
    .Y(_09753_));
 sky130_fd_sc_hd__o22a_1 _16664_ (.A1(_09372_),
    .A2(_09497_),
    .B1(_09633_),
    .B2(_08371_),
    .X(_09754_));
 sky130_fd_sc_hd__a21oi_1 _16665_ (.A1(_09636_),
    .A2(_09753_),
    .B1(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__xor2_1 _16666_ (.A(_09623_),
    .B(_09755_),
    .X(_09756_));
 sky130_fd_sc_hd__xnor2_1 _16667_ (.A(_09752_),
    .B(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__xor2_2 _16668_ (.A(_09750_),
    .B(_09757_),
    .X(_09758_));
 sky130_fd_sc_hd__or2_1 _16669_ (.A(_08362_),
    .B(_09504_),
    .X(_09759_));
 sky130_fd_sc_hd__mux2_2 _16670_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_09510_),
    .S(_06340_),
    .X(_09760_));
 sky130_fd_sc_hd__a21oi_1 _16671_ (.A1(_09515_),
    .A2(_09638_),
    .B1(_08271_),
    .Y(_09761_));
 sky130_fd_sc_hd__and3_1 _16672_ (.A(_08350_),
    .B(_09760_),
    .C(_09761_),
    .X(_09762_));
 sky130_fd_sc_hd__buf_2 _16673_ (.A(_09760_),
    .X(_09763_));
 sky130_fd_sc_hd__a21oi_1 _16674_ (.A1(_08350_),
    .A2(_09763_),
    .B1(_09761_),
    .Y(_09764_));
 sky130_fd_sc_hd__or3_1 _16675_ (.A(_09759_),
    .B(_09762_),
    .C(_09764_),
    .X(_09765_));
 sky130_fd_sc_hd__o21ai_1 _16676_ (.A1(_09762_),
    .A2(_09764_),
    .B1(_09759_),
    .Y(_09766_));
 sky130_fd_sc_hd__and2_1 _16677_ (.A(_09765_),
    .B(_09766_),
    .X(_09767_));
 sky130_fd_sc_hd__or4_1 _16678_ (.A(_08118_),
    .B(_08120_),
    .C(_08122_),
    .D(_09641_),
    .X(_09768_));
 sky130_fd_sc_hd__a21o_1 _16679_ (.A1(_08214_),
    .A2(_09768_),
    .B1(_08327_),
    .X(_09769_));
 sky130_fd_sc_hd__or3_2 _16680_ (.A(_08341_),
    .B(_08298_),
    .C(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__mux2_1 _16681_ (.A0(\rbzero.wall_tracer.visualWallDist[10] ),
    .A1(_09687_),
    .S(_09770_),
    .X(_09771_));
 sky130_fd_sc_hd__nand2_1 _16682_ (.A(\rbzero.wall_tracer.stepDistY[9] ),
    .B(_08304_),
    .Y(_09772_));
 sky130_fd_sc_hd__and2_1 _16683_ (.A(_09772_),
    .B(_09644_),
    .X(_09773_));
 sky130_fd_sc_hd__nor2_1 _16684_ (.A(_08830_),
    .B(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__xor2_1 _16685_ (.A(_09771_),
    .B(_09774_),
    .X(_09775_));
 sky130_fd_sc_hd__or3_1 _16686_ (.A(_08830_),
    .B(_09507_),
    .C(_09645_),
    .X(_09776_));
 sky130_fd_sc_hd__a21bo_1 _16687_ (.A1(_09640_),
    .A2(_09647_),
    .B1_N(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__xnor2_1 _16688_ (.A(_09775_),
    .B(_09777_),
    .Y(_09778_));
 sky130_fd_sc_hd__xnor2_2 _16689_ (.A(_09767_),
    .B(_09778_),
    .Y(_09779_));
 sky130_fd_sc_hd__nor2_1 _16690_ (.A(_09648_),
    .B(_09649_),
    .Y(_09780_));
 sky130_fd_sc_hd__a21o_1 _16691_ (.A1(_09637_),
    .A2(_09650_),
    .B1(_09780_),
    .X(_09781_));
 sky130_fd_sc_hd__xnor2_2 _16692_ (.A(_09779_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__xnor2_2 _16693_ (.A(_09758_),
    .B(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__nor2_1 _16694_ (.A(_09651_),
    .B(_09652_),
    .Y(_09784_));
 sky130_fd_sc_hd__a21o_1 _16695_ (.A1(_09629_),
    .A2(_09653_),
    .B1(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__xnor2_2 _16696_ (.A(_09783_),
    .B(_09785_),
    .Y(_09786_));
 sky130_fd_sc_hd__xnor2_2 _16697_ (.A(_09749_),
    .B(_09786_),
    .Y(_09787_));
 sky130_fd_sc_hd__a21o_1 _16698_ (.A1(_09619_),
    .A2(_09657_),
    .B1(_09656_),
    .X(_09788_));
 sky130_fd_sc_hd__xnor2_2 _16699_ (.A(_09787_),
    .B(_09788_),
    .Y(_09789_));
 sky130_fd_sc_hd__xnor2_2 _16700_ (.A(_09728_),
    .B(_09789_),
    .Y(_09790_));
 sky130_fd_sc_hd__a21oi_1 _16701_ (.A1(_09594_),
    .A2(_09662_),
    .B1(_09660_),
    .Y(_09791_));
 sky130_fd_sc_hd__xor2_2 _16702_ (.A(_09790_),
    .B(_09791_),
    .X(_09792_));
 sky130_fd_sc_hd__xnor2_4 _16703_ (.A(_09693_),
    .B(_09792_),
    .Y(_09793_));
 sky130_fd_sc_hd__a21oi_2 _16704_ (.A1(_09565_),
    .A2(_09666_),
    .B1(_09665_),
    .Y(_09794_));
 sky130_fd_sc_hd__xnor2_4 _16705_ (.A(_09793_),
    .B(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__xor2_4 _16706_ (.A(_09685_),
    .B(_09795_),
    .X(_09796_));
 sky130_fd_sc_hd__xnor2_4 _16707_ (.A(_09684_),
    .B(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__mux2_1 _16708_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_08206_),
    .X(_09798_));
 sky130_fd_sc_hd__xnor2_1 _16709_ (.A(_09202_),
    .B(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__xnor2_1 _16710_ (.A(_09797_),
    .B(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__xnor2_1 _16711_ (.A(_09683_),
    .B(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__nand2_1 _16712_ (.A(_08211_),
    .B(_09801_),
    .Y(_09802_));
 sky130_fd_sc_hd__o211a_1 _16713_ (.A1(\rbzero.texu_hot[5] ),
    .A2(_08211_),
    .B1(_09802_),
    .C1(_04500_),
    .X(_00471_));
 sky130_fd_sc_hd__nor2_1 _16714_ (.A(_05105_),
    .B(_04761_),
    .Y(_09803_));
 sky130_fd_sc_hd__and4_1 _16715_ (.A(_04643_),
    .B(_04709_),
    .C(_09803_),
    .D(_05098_),
    .X(_09804_));
 sky130_fd_sc_hd__buf_4 _16716_ (.A(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__or2_1 _16717_ (.A(_04469_),
    .B(_09805_),
    .X(_09806_));
 sky130_fd_sc_hd__buf_2 _16718_ (.A(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__nor2_1 _16719_ (.A(_04030_),
    .B(_09807_),
    .Y(_00472_));
 sky130_fd_sc_hd__clkbuf_8 _16720_ (.A(_04112_),
    .X(_09808_));
 sky130_fd_sc_hd__and3b_1 _16721_ (.A_N(_04707_),
    .B(_09808_),
    .C(_04509_),
    .X(_09809_));
 sky130_fd_sc_hd__clkbuf_1 _16722_ (.A(_09809_),
    .X(_00473_));
 sky130_fd_sc_hd__buf_4 _16723_ (.A(_04112_),
    .X(_09810_));
 sky130_fd_sc_hd__or2_1 _16724_ (.A(_04506_),
    .B(_04707_),
    .X(_09811_));
 sky130_fd_sc_hd__and3_1 _16725_ (.A(_09810_),
    .B(_04708_),
    .C(_09811_),
    .X(_09812_));
 sky130_fd_sc_hd__clkbuf_1 _16726_ (.A(_09812_),
    .X(_00474_));
 sky130_fd_sc_hd__buf_4 _16727_ (.A(_04470_),
    .X(_09813_));
 sky130_fd_sc_hd__nor2_1 _16728_ (.A(_09813_),
    .B(_05110_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _16729_ (.A(_05125_),
    .B(_09807_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _16730_ (.A(_05130_),
    .B(_09807_),
    .Y(_00477_));
 sky130_fd_sc_hd__nor2_1 _16731_ (.A(_05108_),
    .B(_09807_),
    .Y(_00478_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_05148_),
    .B(_09807_),
    .Y(_00479_));
 sky130_fd_sc_hd__and3_1 _16733_ (.A(_04033_),
    .B(_04696_),
    .C(_05337_),
    .X(_09814_));
 sky130_fd_sc_hd__a21o_1 _16734_ (.A1(_04696_),
    .A2(_05337_),
    .B1(_04033_),
    .X(_09815_));
 sky130_fd_sc_hd__nor2_4 _16735_ (.A(_04469_),
    .B(_09805_),
    .Y(_09816_));
 sky130_fd_sc_hd__and3b_1 _16736_ (.A_N(_09814_),
    .B(_09815_),
    .C(_09816_),
    .X(_09817_));
 sky130_fd_sc_hd__clkbuf_1 _16737_ (.A(_09817_),
    .X(_00480_));
 sky130_fd_sc_hd__a21oi_1 _16738_ (.A1(_04034_),
    .A2(_09814_),
    .B1(_09807_),
    .Y(_09818_));
 sky130_fd_sc_hd__o21a_1 _16739_ (.A1(_04034_),
    .A2(_09814_),
    .B1(_09818_),
    .X(_00481_));
 sky130_fd_sc_hd__and3_1 _16740_ (.A(_04494_),
    .B(_05095_),
    .C(_09805_),
    .X(_09819_));
 sky130_fd_sc_hd__nor2_1 _16741_ (.A(_04489_),
    .B(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__clkbuf_4 _16742_ (.A(_09820_),
    .X(_09821_));
 sky130_fd_sc_hd__buf_4 _16743_ (.A(_09821_),
    .X(_09822_));
 sky130_fd_sc_hd__buf_4 _16744_ (.A(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__and4_1 _16745_ (.A(_04495_),
    .B(_04490_),
    .C(_05095_),
    .D(_09805_),
    .X(_09824_));
 sky130_fd_sc_hd__clkbuf_4 _16746_ (.A(_09824_),
    .X(_09825_));
 sky130_fd_sc_hd__buf_6 _16747_ (.A(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__clkbuf_4 _16748_ (.A(_09826_),
    .X(_09827_));
 sky130_fd_sc_hd__a22o_1 _16749_ (.A1(\rbzero.row_render.side ),
    .A2(_09823_),
    .B1(_09827_),
    .B2(_08206_),
    .X(_00482_));
 sky130_fd_sc_hd__a22o_1 _16750_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_09823_),
    .B1(_09827_),
    .B2(_08005_),
    .X(_00483_));
 sky130_fd_sc_hd__a22o_1 _16751_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_09823_),
    .B1(_09827_),
    .B2(_08017_),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _16752_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_09823_),
    .B1(_09827_),
    .B2(_08030_),
    .X(_00485_));
 sky130_fd_sc_hd__nand4_4 _16753_ (.A(_04495_),
    .B(_04491_),
    .C(_05095_),
    .D(_09805_),
    .Y(_09828_));
 sky130_fd_sc_hd__a2bb2o_1 _16754_ (.A1_N(_08040_),
    .A2_N(_09828_),
    .B1(_09823_),
    .B2(\rbzero.row_render.size[3] ),
    .X(_00486_));
 sky130_fd_sc_hd__a22o_1 _16755_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_09823_),
    .B1(_09827_),
    .B2(_08049_),
    .X(_00487_));
 sky130_fd_sc_hd__a2bb2o_1 _16756_ (.A1_N(_08057_),
    .A2_N(_09828_),
    .B1(_09823_),
    .B2(\rbzero.row_render.size[5] ),
    .X(_00488_));
 sky130_fd_sc_hd__buf_4 _16757_ (.A(_09820_),
    .X(_09829_));
 sky130_fd_sc_hd__clkbuf_4 _16758_ (.A(_09829_),
    .X(_09830_));
 sky130_fd_sc_hd__a22o_1 _16759_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_09830_),
    .B1(_09827_),
    .B2(_08061_),
    .X(_00489_));
 sky130_fd_sc_hd__a22o_1 _16760_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_09830_),
    .B1(_09827_),
    .B2(_08069_),
    .X(_00490_));
 sky130_fd_sc_hd__a22o_1 _16761_ (.A1(\rbzero.row_render.size[8] ),
    .A2(_09830_),
    .B1(_09827_),
    .B2(_08078_),
    .X(_00491_));
 sky130_fd_sc_hd__a22o_1 _16762_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_09830_),
    .B1(_09827_),
    .B2(_08084_),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _16763_ (.A1(\rbzero.row_render.size[10] ),
    .A2(_09830_),
    .B1(_09827_),
    .B2(_08090_),
    .X(_00493_));
 sky130_fd_sc_hd__clkbuf_4 _16764_ (.A(_09826_),
    .X(_09831_));
 sky130_fd_sc_hd__a22o_1 _16765_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_09830_),
    .B1(_09831_),
    .B2(\rbzero.texu_hot[0] ),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _16766_ (.A1(\rbzero.row_render.texu[1] ),
    .A2(_09830_),
    .B1(_09831_),
    .B2(\rbzero.texu_hot[1] ),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _16767_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_09830_),
    .B1(_09831_),
    .B2(net514),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_1 _16768_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(_09830_),
    .B1(_09831_),
    .B2(net515),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _16769_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_09830_),
    .B1(_09831_),
    .B2(net516),
    .X(_00498_));
 sky130_fd_sc_hd__buf_2 _16770_ (.A(_09829_),
    .X(_09832_));
 sky130_fd_sc_hd__a22o_1 _16771_ (.A1(\rbzero.traced_texa[-11] ),
    .A2(_09832_),
    .B1(_09831_),
    .B2(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _16772_ (.A1(\rbzero.traced_texa[-10] ),
    .A2(_09832_),
    .B1(_09831_),
    .B2(_08131_),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _16773_ (.A1(\rbzero.traced_texa[-9] ),
    .A2(_09832_),
    .B1(_09831_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_1 _16774_ (.A1(\rbzero.traced_texa[-8] ),
    .A2(_09832_),
    .B1(_09831_),
    .B2(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _16775_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(_09832_),
    .B1(_09831_),
    .B2(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(_00503_));
 sky130_fd_sc_hd__buf_2 _16776_ (.A(_09825_),
    .X(_09833_));
 sky130_fd_sc_hd__a22o_1 _16777_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(_09832_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _16778_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(_09832_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _16779_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(_09832_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(_00506_));
 sky130_fd_sc_hd__a22o_1 _16780_ (.A1(\rbzero.traced_texa[-3] ),
    .A2(_09832_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _16781_ (.A1(\rbzero.traced_texa[-2] ),
    .A2(_09832_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_00508_));
 sky130_fd_sc_hd__buf_2 _16782_ (.A(_09829_),
    .X(_09834_));
 sky130_fd_sc_hd__a22o_1 _16783_ (.A1(\rbzero.traced_texa[-1] ),
    .A2(_09834_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_00509_));
 sky130_fd_sc_hd__a22o_1 _16784_ (.A1(\rbzero.traced_texa[0] ),
    .A2(_09834_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_00510_));
 sky130_fd_sc_hd__a22o_1 _16785_ (.A1(\rbzero.traced_texa[1] ),
    .A2(_09834_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_00511_));
 sky130_fd_sc_hd__a22o_1 _16786_ (.A1(\rbzero.traced_texa[2] ),
    .A2(_09834_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _16787_ (.A1(\rbzero.traced_texa[3] ),
    .A2(_09834_),
    .B1(_09833_),
    .B2(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(_00513_));
 sky130_fd_sc_hd__clkbuf_4 _16788_ (.A(_09825_),
    .X(_09835_));
 sky130_fd_sc_hd__a22o_1 _16789_ (.A1(\rbzero.traced_texa[4] ),
    .A2(_09834_),
    .B1(_09835_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_1 _16790_ (.A1(\rbzero.traced_texa[5] ),
    .A2(_09834_),
    .B1(_09835_),
    .B2(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _16791_ (.A1(\rbzero.traced_texa[6] ),
    .A2(_09834_),
    .B1(_09835_),
    .B2(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_00516_));
 sky130_fd_sc_hd__a22o_1 _16792_ (.A1(\rbzero.traced_texa[7] ),
    .A2(_09834_),
    .B1(_09835_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _16793_ (.A1(\rbzero.traced_texa[8] ),
    .A2(_09834_),
    .B1(_09835_),
    .B2(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_00518_));
 sky130_fd_sc_hd__buf_2 _16794_ (.A(_09829_),
    .X(_09836_));
 sky130_fd_sc_hd__a22o_1 _16795_ (.A1(\rbzero.traced_texa[9] ),
    .A2(_09836_),
    .B1(_09835_),
    .B2(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_00519_));
 sky130_fd_sc_hd__a22o_1 _16796_ (.A1(\rbzero.traced_texa[10] ),
    .A2(_09836_),
    .B1(_09835_),
    .B2(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _16797_ (.A0(_04603_),
    .A1(\rbzero.row_render.wall[0] ),
    .S(_09828_),
    .X(_09837_));
 sky130_fd_sc_hd__clkbuf_1 _16798_ (.A(_09837_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _16799_ (.A0(\rbzero.wall_hot[1] ),
    .A1(\rbzero.row_render.wall[1] ),
    .S(_09828_),
    .X(_09838_));
 sky130_fd_sc_hd__clkbuf_1 _16800_ (.A(_09838_),
    .X(_00522_));
 sky130_fd_sc_hd__o21a_1 _16801_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(\rbzero.wall_tracer.mapX[5] ),
    .B1(_09199_),
    .X(_09839_));
 sky130_fd_sc_hd__xor2_1 _16802_ (.A(\rbzero.wall_tracer.mapX[5] ),
    .B(_09199_),
    .X(_09840_));
 sky130_fd_sc_hd__xnor2_1 _16803_ (.A(_06241_),
    .B(_09199_),
    .Y(_09841_));
 sky130_fd_sc_hd__or2_1 _16804_ (.A(_06259_),
    .B(_09199_),
    .X(_09842_));
 sky130_fd_sc_hd__xnor2_1 _16805_ (.A(_06286_),
    .B(_08285_),
    .Y(_09843_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(\rbzero.map_rom.f4 ),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__a21bo_1 _16807_ (.A1(\rbzero.map_rom.f3 ),
    .A2(_09199_),
    .B1_N(_09844_),
    .X(_09845_));
 sky130_fd_sc_hd__and2_1 _16808_ (.A(\rbzero.map_rom.f2 ),
    .B(_08285_),
    .X(_09846_));
 sky130_fd_sc_hd__nor2_1 _16809_ (.A(\rbzero.map_rom.f2 ),
    .B(_08285_),
    .Y(_09847_));
 sky130_fd_sc_hd__nor2_1 _16810_ (.A(_09846_),
    .B(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__a21o_1 _16811_ (.A1(_09845_),
    .A2(_09848_),
    .B1(_09846_),
    .X(_09849_));
 sky130_fd_sc_hd__nand2_1 _16812_ (.A(_06259_),
    .B(_09199_),
    .Y(_09850_));
 sky130_fd_sc_hd__or2b_1 _16813_ (.A(_09849_),
    .B_N(_09850_),
    .X(_09851_));
 sky130_fd_sc_hd__and3_2 _16814_ (.A(_09841_),
    .B(_09842_),
    .C(_09851_),
    .X(_09852_));
 sky130_fd_sc_hd__and2_1 _16815_ (.A(_09840_),
    .B(_09852_),
    .X(_09853_));
 sky130_fd_sc_hd__xor2_1 _16816_ (.A(\rbzero.wall_tracer.mapX[6] ),
    .B(_09199_),
    .X(_09854_));
 sky130_fd_sc_hd__o21ai_1 _16817_ (.A1(_09839_),
    .A2(_09853_),
    .B1(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__or3_1 _16818_ (.A(_09854_),
    .B(_09839_),
    .C(_09853_),
    .X(_09856_));
 sky130_fd_sc_hd__nand2_2 _16819_ (.A(_06342_),
    .B(_08125_),
    .Y(_09857_));
 sky130_fd_sc_hd__nor2_2 _16820_ (.A(_06164_),
    .B(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__buf_8 _16821_ (.A(_09857_),
    .X(_09859_));
 sky130_fd_sc_hd__buf_4 _16822_ (.A(_09859_),
    .X(_09860_));
 sky130_fd_sc_hd__a32o_1 _16823_ (.A1(_09855_),
    .A2(_09856_),
    .A3(_09858_),
    .B1(_09860_),
    .B2(\rbzero.wall_tracer.mapX[6] ),
    .X(_00523_));
 sky130_fd_sc_hd__xor2_1 _16824_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(_09199_),
    .X(_09861_));
 sky130_fd_sc_hd__a21boi_1 _16825_ (.A1(\rbzero.wall_tracer.mapX[6] ),
    .A2(_09200_),
    .B1_N(_09855_),
    .Y(_09862_));
 sky130_fd_sc_hd__xnor2_1 _16826_ (.A(_09861_),
    .B(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__a22o_1 _16827_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(_09860_),
    .B1(_09858_),
    .B2(_09863_),
    .X(_00524_));
 sky130_fd_sc_hd__xor2_1 _16828_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(_09200_),
    .X(_09864_));
 sky130_fd_sc_hd__and3_1 _16829_ (.A(_09854_),
    .B(_09853_),
    .C(_09861_),
    .X(_09865_));
 sky130_fd_sc_hd__o21a_1 _16830_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(\rbzero.wall_tracer.mapX[6] ),
    .B1(_09199_),
    .X(_09866_));
 sky130_fd_sc_hd__or3_1 _16831_ (.A(_09839_),
    .B(_09865_),
    .C(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__xor2_1 _16832_ (.A(_09864_),
    .B(_09867_),
    .X(_09868_));
 sky130_fd_sc_hd__a22o_1 _16833_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09860_),
    .B1(_09858_),
    .B2(_09868_),
    .X(_00525_));
 sky130_fd_sc_hd__a22o_1 _16834_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09200_),
    .B1(_09864_),
    .B2(_09867_),
    .X(_09869_));
 sky130_fd_sc_hd__xnor2_1 _16835_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(_09200_),
    .Y(_09870_));
 sky130_fd_sc_hd__xnor2_1 _16836_ (.A(_09869_),
    .B(_09870_),
    .Y(_09871_));
 sky130_fd_sc_hd__a22o_1 _16837_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09860_),
    .B1(_09858_),
    .B2(_09871_),
    .X(_00526_));
 sky130_fd_sc_hd__o21a_1 _16838_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09200_),
    .B1(_09869_),
    .X(_09872_));
 sky130_fd_sc_hd__a21oi_1 _16839_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09200_),
    .B1(_09872_),
    .Y(_09873_));
 sky130_fd_sc_hd__xnor2_1 _16840_ (.A(\rbzero.wall_tracer.mapX[10] ),
    .B(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__nand2_1 _16841_ (.A(_09200_),
    .B(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__or2_1 _16842_ (.A(_09200_),
    .B(_09874_),
    .X(_09876_));
 sky130_fd_sc_hd__a32o_1 _16843_ (.A1(_09858_),
    .A2(_09875_),
    .A3(_09876_),
    .B1(_09860_),
    .B2(\rbzero.wall_tracer.mapX[10] ),
    .X(_00527_));
 sky130_fd_sc_hd__nor2_1 _16844_ (.A(_08934_),
    .B(_08982_),
    .Y(_09877_));
 sky130_fd_sc_hd__a211o_2 _16845_ (.A1(_08934_),
    .A2(_08982_),
    .B1(_09877_),
    .C1(_08195_),
    .X(_09878_));
 sky130_fd_sc_hd__o21ai_1 _16846_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_08194_),
    .Y(_09879_));
 sky130_fd_sc_hd__a21oi_1 _16847_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__nor2_1 _16848_ (.A(_09859_),
    .B(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__inv_2 _16849_ (.A(_09857_),
    .Y(_09882_));
 sky130_fd_sc_hd__clkbuf_8 _16850_ (.A(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__buf_4 _16851_ (.A(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__o2bb2a_1 _16852_ (.A1_N(_09878_),
    .A2_N(_09881_),
    .B1(\rbzero.wall_tracer.trackDistX[-11] ),
    .B2(_09884_),
    .X(_00528_));
 sky130_fd_sc_hd__and2_1 _16853_ (.A(_08896_),
    .B(_08984_),
    .X(_09885_));
 sky130_fd_sc_hd__nor2_1 _16854_ (.A(_08896_),
    .B(_08984_),
    .Y(_09886_));
 sky130_fd_sc_hd__or3_2 _16855_ (.A(_08194_),
    .B(_09885_),
    .C(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__or2_1 _16856_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_09888_));
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_09889_));
 sky130_fd_sc_hd__and4_1 _16858_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .C(_09888_),
    .D(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__a22oi_1 _16859_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09888_),
    .B2(_09889_),
    .Y(_09891_));
 sky130_fd_sc_hd__o31a_1 _16860_ (.A1(_08156_),
    .A2(_09890_),
    .A3(_09891_),
    .B1(_09883_),
    .X(_09892_));
 sky130_fd_sc_hd__o2bb2a_1 _16861_ (.A1_N(_09887_),
    .A2_N(_09892_),
    .B1(\rbzero.wall_tracer.trackDistX[-10] ),
    .B2(_09884_),
    .X(_00529_));
 sky130_fd_sc_hd__a21oi_2 _16862_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(\rbzero.wall_tracer.stepDistX[-10] ),
    .B1(_09890_),
    .Y(_09893_));
 sky130_fd_sc_hd__nor2_1 _16863_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .Y(_09894_));
 sky130_fd_sc_hd__and2_1 _16864_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_09895_));
 sky130_fd_sc_hd__nor3_1 _16865_ (.A(_09893_),
    .B(_09894_),
    .C(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__o21a_1 _16866_ (.A1(_09894_),
    .A2(_09895_),
    .B1(_09893_),
    .X(_09897_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(_06164_),
    .B(_09189_),
    .Y(_09898_));
 sky130_fd_sc_hd__o311a_1 _16868_ (.A1(_06164_),
    .A2(_09896_),
    .A3(_09897_),
    .B1(_09883_),
    .C1(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__a21oi_1 _16869_ (.A1(_06188_),
    .A2(_09860_),
    .B1(_09899_),
    .Y(_00530_));
 sky130_fd_sc_hd__or2_1 _16870_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_09900_));
 sky130_fd_sc_hd__nand2_1 _16871_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_09901_));
 sky130_fd_sc_hd__o21bai_2 _16872_ (.A1(_09893_),
    .A2(_09894_),
    .B1_N(_09895_),
    .Y(_09902_));
 sky130_fd_sc_hd__and3_1 _16873_ (.A(_09900_),
    .B(_09901_),
    .C(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__a21oi_1 _16874_ (.A1(_09900_),
    .A2(_09901_),
    .B1(_09902_),
    .Y(_09904_));
 sky130_fd_sc_hd__buf_6 _16875_ (.A(_06163_),
    .X(_09905_));
 sky130_fd_sc_hd__nand2_1 _16876_ (.A(_09905_),
    .B(_09193_),
    .Y(_09906_));
 sky130_fd_sc_hd__o311a_1 _16877_ (.A1(_06164_),
    .A2(_09903_),
    .A3(_09904_),
    .B1(_09883_),
    .C1(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__a21oi_1 _16878_ (.A1(_06215_),
    .A2(_09860_),
    .B1(_09907_),
    .Y(_00531_));
 sky130_fd_sc_hd__nor2_1 _16879_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09908_));
 sky130_fd_sc_hd__nand2_1 _16880_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09909_));
 sky130_fd_sc_hd__or2b_1 _16881_ (.A(_09908_),
    .B_N(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__a21boi_1 _16882_ (.A1(_09900_),
    .A2(_09902_),
    .B1_N(_09901_),
    .Y(_09911_));
 sky130_fd_sc_hd__nor2_1 _16883_ (.A(_09910_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__a21o_1 _16884_ (.A1(_09910_),
    .A2(_09911_),
    .B1(_08155_),
    .X(_09913_));
 sky130_fd_sc_hd__xor2_2 _16885_ (.A(_08993_),
    .B(_09086_),
    .X(_09914_));
 sky130_fd_sc_hd__nand2_1 _16886_ (.A(_09905_),
    .B(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__o21ai_1 _16887_ (.A1(_09912_),
    .A2(_09913_),
    .B1(_09915_),
    .Y(_09916_));
 sky130_fd_sc_hd__buf_4 _16888_ (.A(_09882_),
    .X(_09917_));
 sky130_fd_sc_hd__mux2_1 _16889_ (.A0(\rbzero.wall_tracer.trackDistX[-7] ),
    .A1(_09916_),
    .S(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__clkbuf_1 _16890_ (.A(_09918_),
    .X(_00532_));
 sky130_fd_sc_hd__or2_1 _16891_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_09919_));
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_09920_));
 sky130_fd_sc_hd__o21ai_1 _16893_ (.A1(_09908_),
    .A2(_09911_),
    .B1(_09909_),
    .Y(_09921_));
 sky130_fd_sc_hd__and3_1 _16894_ (.A(_09919_),
    .B(_09920_),
    .C(_09921_),
    .X(_09922_));
 sky130_fd_sc_hd__a21oi_1 _16895_ (.A1(_09919_),
    .A2(_09920_),
    .B1(_09921_),
    .Y(_09923_));
 sky130_fd_sc_hd__or2_1 _16896_ (.A(_08194_),
    .B(_09183_),
    .X(_09924_));
 sky130_fd_sc_hd__o311a_1 _16897_ (.A1(_06164_),
    .A2(_09922_),
    .A3(_09923_),
    .B1(_09917_),
    .C1(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__a21oi_1 _16898_ (.A1(_06200_),
    .A2(_09860_),
    .B1(_09925_),
    .Y(_00533_));
 sky130_fd_sc_hd__xor2_2 _16899_ (.A(_09206_),
    .B(_09300_),
    .X(_09926_));
 sky130_fd_sc_hd__nand2_1 _16900_ (.A(_08155_),
    .B(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__nor2_1 _16901_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09928_));
 sky130_fd_sc_hd__nand2_1 _16902_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09929_));
 sky130_fd_sc_hd__or2b_1 _16903_ (.A(_09928_),
    .B_N(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__a21boi_1 _16904_ (.A1(_09919_),
    .A2(_09921_),
    .B1_N(_09920_),
    .Y(_09931_));
 sky130_fd_sc_hd__xor2_1 _16905_ (.A(_09930_),
    .B(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__a21oi_1 _16906_ (.A1(_08195_),
    .A2(_09932_),
    .B1(_09859_),
    .Y(_09933_));
 sky130_fd_sc_hd__o2bb2a_1 _16907_ (.A1_N(_09927_),
    .A2_N(_09933_),
    .B1(\rbzero.wall_tracer.trackDistX[-5] ),
    .B2(_09884_),
    .X(_00534_));
 sky130_fd_sc_hd__or2_1 _16908_ (.A(_08195_),
    .B(_09422_),
    .X(_09934_));
 sky130_fd_sc_hd__or2_1 _16909_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(_09935_));
 sky130_fd_sc_hd__nand2_1 _16910_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09936_));
 sky130_fd_sc_hd__o21ai_1 _16911_ (.A1(_09928_),
    .A2(_09931_),
    .B1(_09929_),
    .Y(_09937_));
 sky130_fd_sc_hd__and3_1 _16912_ (.A(_09935_),
    .B(_09936_),
    .C(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__a21oi_1 _16913_ (.A1(_09935_),
    .A2(_09936_),
    .B1(_09937_),
    .Y(_09939_));
 sky130_fd_sc_hd__o31a_1 _16914_ (.A1(_08156_),
    .A2(_09938_),
    .A3(_09939_),
    .B1(_09883_),
    .X(_09940_));
 sky130_fd_sc_hd__o2bb2a_1 _16915_ (.A1_N(_09934_),
    .A2_N(_09940_),
    .B1(\rbzero.wall_tracer.trackDistX[-4] ),
    .B2(_09884_),
    .X(_00535_));
 sky130_fd_sc_hd__nor2_1 _16916_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09942_));
 sky130_fd_sc_hd__or2b_1 _16918_ (.A(_09941_),
    .B_N(_09942_),
    .X(_09943_));
 sky130_fd_sc_hd__a21boi_1 _16919_ (.A1(_09935_),
    .A2(_09937_),
    .B1_N(_09936_),
    .Y(_09944_));
 sky130_fd_sc_hd__nor2_1 _16920_ (.A(_09943_),
    .B(_09944_),
    .Y(_09945_));
 sky130_fd_sc_hd__a21o_1 _16921_ (.A1(_09943_),
    .A2(_09944_),
    .B1(_08155_),
    .X(_09946_));
 sky130_fd_sc_hd__xnor2_4 _16922_ (.A(_09434_),
    .B(_09558_),
    .Y(_09947_));
 sky130_fd_sc_hd__nand2_1 _16923_ (.A(_09905_),
    .B(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__o21ai_1 _16924_ (.A1(_09945_),
    .A2(_09946_),
    .B1(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__mux2_1 _16925_ (.A0(\rbzero.wall_tracer.trackDistX[-3] ),
    .A1(_09949_),
    .S(_09917_),
    .X(_09950_));
 sky130_fd_sc_hd__clkbuf_1 _16926_ (.A(_09950_),
    .X(_00536_));
 sky130_fd_sc_hd__or2_1 _16927_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_09951_));
 sky130_fd_sc_hd__nand2_1 _16928_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_09952_));
 sky130_fd_sc_hd__o21ai_1 _16929_ (.A1(_09941_),
    .A2(_09944_),
    .B1(_09942_),
    .Y(_09953_));
 sky130_fd_sc_hd__and3_1 _16930_ (.A(_09951_),
    .B(_09952_),
    .C(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__a21oi_1 _16931_ (.A1(_09951_),
    .A2(_09952_),
    .B1(_09953_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand2_1 _16932_ (.A(_09905_),
    .B(_09673_),
    .Y(_09956_));
 sky130_fd_sc_hd__o311a_1 _16933_ (.A1(_06164_),
    .A2(_09954_),
    .A3(_09955_),
    .B1(_09917_),
    .C1(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__a21oi_1 _16934_ (.A1(_06170_),
    .A2(_09860_),
    .B1(_09957_),
    .Y(_00537_));
 sky130_fd_sc_hd__nor2_1 _16935_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_09958_));
 sky130_fd_sc_hd__and2_1 _16936_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(_09959_));
 sky130_fd_sc_hd__or2_1 _16937_ (.A(_09958_),
    .B(_09959_),
    .X(_09960_));
 sky130_fd_sc_hd__a21boi_1 _16938_ (.A1(_09951_),
    .A2(_09953_),
    .B1_N(_09952_),
    .Y(_09961_));
 sky130_fd_sc_hd__nor2_1 _16939_ (.A(_09960_),
    .B(_09961_),
    .Y(_09962_));
 sky130_fd_sc_hd__a21o_1 _16940_ (.A1(_09960_),
    .A2(_09961_),
    .B1(_08155_),
    .X(_09963_));
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(_09905_),
    .B(_09797_),
    .Y(_09964_));
 sky130_fd_sc_hd__o21ai_1 _16942_ (.A1(_09962_),
    .A2(_09963_),
    .B1(_09964_),
    .Y(_09965_));
 sky130_fd_sc_hd__mux2_1 _16943_ (.A0(\rbzero.wall_tracer.trackDistX[-1] ),
    .A1(_09965_),
    .S(_09917_),
    .X(_09966_));
 sky130_fd_sc_hd__clkbuf_1 _16944_ (.A(_09966_),
    .X(_00538_));
 sky130_fd_sc_hd__nor2_1 _16945_ (.A(_09793_),
    .B(_09794_),
    .Y(_09967_));
 sky130_fd_sc_hd__o21ai_1 _16946_ (.A1(_09574_),
    .A2(_09686_),
    .B1(_09688_),
    .Y(_09968_));
 sky130_fd_sc_hd__or2b_1 _16947_ (.A(_09727_),
    .B_N(_09695_),
    .X(_09969_));
 sky130_fd_sc_hd__o2bb2a_1 _16948_ (.A1_N(_09705_),
    .A2_N(_09707_),
    .B1(_09702_),
    .B2(_09704_),
    .X(_09970_));
 sky130_fd_sc_hd__a21oi_2 _16949_ (.A1(_09725_),
    .A2(_09969_),
    .B1(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__and3_1 _16950_ (.A(_09725_),
    .B(_09969_),
    .C(_09970_),
    .X(_09972_));
 sky130_fd_sc_hd__nor2_1 _16951_ (.A(_09971_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__a21o_1 _16952_ (.A1(_09708_),
    .A2(_09723_),
    .B1(_09721_),
    .X(_09974_));
 sky130_fd_sc_hd__or2b_1 _16953_ (.A(_09747_),
    .B_N(_09731_),
    .X(_09975_));
 sky130_fd_sc_hd__or2b_1 _16954_ (.A(_09748_),
    .B_N(_09729_),
    .X(_09976_));
 sky130_fd_sc_hd__nor2_1 _16955_ (.A(_08959_),
    .B(_09440_),
    .Y(_09977_));
 sky130_fd_sc_hd__xor2_1 _16956_ (.A(_09697_),
    .B(_09977_),
    .X(_09978_));
 sky130_fd_sc_hd__nor2_1 _16957_ (.A(_08567_),
    .B(_09571_),
    .Y(_09979_));
 sky130_fd_sc_hd__and2_1 _16958_ (.A(_09978_),
    .B(_09979_),
    .X(_09980_));
 sky130_fd_sc_hd__nor2_1 _16959_ (.A(_09978_),
    .B(_09979_),
    .Y(_09981_));
 sky130_fd_sc_hd__or2_1 _16960_ (.A(_09980_),
    .B(_09981_),
    .X(_09982_));
 sky130_fd_sc_hd__a21oi_1 _16961_ (.A1(_09578_),
    .A2(_09697_),
    .B1(_09700_),
    .Y(_09983_));
 sky130_fd_sc_hd__nor2_1 _16962_ (.A(_09982_),
    .B(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__nand2_1 _16963_ (.A(_09982_),
    .B(_09983_),
    .Y(_09985_));
 sky130_fd_sc_hd__or2b_1 _16964_ (.A(_09984_),
    .B_N(_09985_),
    .X(_09986_));
 sky130_fd_sc_hd__nor2_1 _16965_ (.A(_08504_),
    .B(_09687_),
    .Y(_09987_));
 sky130_fd_sc_hd__xnor2_1 _16966_ (.A(_09986_),
    .B(_09987_),
    .Y(_09988_));
 sky130_fd_sc_hd__a21bo_1 _16967_ (.A1(_09579_),
    .A2(_09714_),
    .B1_N(_09713_),
    .X(_09989_));
 sky130_fd_sc_hd__o21a_1 _16968_ (.A1(_08783_),
    .A2(_09156_),
    .B1(_09712_),
    .X(_09990_));
 sky130_fd_sc_hd__or3_1 _16969_ (.A(_08783_),
    .B(_09156_),
    .C(_09712_),
    .X(_09991_));
 sky130_fd_sc_hd__or2b_1 _16970_ (.A(_09990_),
    .B_N(_09991_),
    .X(_09992_));
 sky130_fd_sc_hd__or2_1 _16971_ (.A(_08831_),
    .B(_09212_),
    .X(_09993_));
 sky130_fd_sc_hd__xnor2_1 _16972_ (.A(_09992_),
    .B(_09993_),
    .Y(_09994_));
 sky130_fd_sc_hd__a22o_1 _16973_ (.A1(_09733_),
    .A2(_09734_),
    .B1(_09735_),
    .B2(_09732_),
    .X(_09995_));
 sky130_fd_sc_hd__and2b_1 _16974_ (.A_N(_09994_),
    .B(_09995_),
    .X(_09996_));
 sky130_fd_sc_hd__and2b_1 _16975_ (.A_N(_09995_),
    .B(_09994_),
    .X(_09997_));
 sky130_fd_sc_hd__nor2_1 _16976_ (.A(_09996_),
    .B(_09997_),
    .Y(_09998_));
 sky130_fd_sc_hd__xnor2_1 _16977_ (.A(_09989_),
    .B(_09998_),
    .Y(_09999_));
 sky130_fd_sc_hd__a21oi_1 _16978_ (.A1(_09710_),
    .A2(_09718_),
    .B1(_09716_),
    .Y(_10000_));
 sky130_fd_sc_hd__xor2_1 _16979_ (.A(_09999_),
    .B(_10000_),
    .X(_10001_));
 sky130_fd_sc_hd__nand2_1 _16980_ (.A(_09988_),
    .B(_10001_),
    .Y(_10002_));
 sky130_fd_sc_hd__or2_1 _16981_ (.A(_09988_),
    .B(_10001_),
    .X(_10003_));
 sky130_fd_sc_hd__nand2_1 _16982_ (.A(_10002_),
    .B(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__a21o_1 _16983_ (.A1(_09975_),
    .A2(_09976_),
    .B1(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__nand3_1 _16984_ (.A(_09975_),
    .B(_09976_),
    .C(_10004_),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_1 _16985_ (.A(_10005_),
    .B(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__xnor2_1 _16986_ (.A(_09974_),
    .B(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__a21o_1 _16987_ (.A1(_09736_),
    .A2(_09745_),
    .B1(_09744_),
    .X(_10009_));
 sky130_fd_sc_hd__and2b_1 _16988_ (.A_N(_09752_),
    .B(_09756_),
    .X(_10010_));
 sky130_fd_sc_hd__a21o_1 _16989_ (.A1(_09750_),
    .A2(_09757_),
    .B1(_10010_),
    .X(_10011_));
 sky130_fd_sc_hd__clkbuf_4 _16990_ (.A(_08661_),
    .X(_10012_));
 sky130_fd_sc_hd__a21oi_2 _16991_ (.A1(_08493_),
    .A2(_08238_),
    .B1(_08240_),
    .Y(_10013_));
 sky130_fd_sc_hd__nor2_1 _16992_ (.A(_08510_),
    .B(_10013_),
    .Y(_10014_));
 sky130_fd_sc_hd__o22a_1 _16993_ (.A1(_08495_),
    .A2(_10013_),
    .B1(_08293_),
    .B2(_08510_),
    .X(_10015_));
 sky130_fd_sc_hd__a21o_1 _16994_ (.A1(_09734_),
    .A2(_10014_),
    .B1(_10015_),
    .X(_10016_));
 sky130_fd_sc_hd__or3_1 _16995_ (.A(_10012_),
    .B(_09072_),
    .C(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__o21ai_1 _16996_ (.A1(_10012_),
    .A2(_09072_),
    .B1(_10016_),
    .Y(_10018_));
 sky130_fd_sc_hd__and2_1 _16997_ (.A(_10017_),
    .B(_10018_),
    .X(_10019_));
 sky130_fd_sc_hd__nor2_1 _16998_ (.A(_08559_),
    .B(_08307_),
    .Y(_10020_));
 sky130_fd_sc_hd__xnor2_1 _16999_ (.A(_09737_),
    .B(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__nor2_1 _17000_ (.A(_08551_),
    .B(_09007_),
    .Y(_10022_));
 sky130_fd_sc_hd__nand2_1 _17001_ (.A(_10021_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__or2_1 _17002_ (.A(_10021_),
    .B(_10022_),
    .X(_10024_));
 sky130_fd_sc_hd__nand2_1 _17003_ (.A(_10023_),
    .B(_10024_),
    .Y(_10025_));
 sky130_fd_sc_hd__a21oi_1 _17004_ (.A1(_09605_),
    .A2(_09741_),
    .B1(_09738_),
    .Y(_10026_));
 sky130_fd_sc_hd__nor2_1 _17005_ (.A(_10025_),
    .B(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__and2_1 _17006_ (.A(_10025_),
    .B(_10026_),
    .X(_10028_));
 sky130_fd_sc_hd__nor2_1 _17007_ (.A(_10027_),
    .B(_10028_),
    .Y(_10029_));
 sky130_fd_sc_hd__xnor2_1 _17008_ (.A(_10019_),
    .B(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__xor2_1 _17009_ (.A(_10011_),
    .B(_10030_),
    .X(_10031_));
 sky130_fd_sc_hd__xnor2_1 _17010_ (.A(_10009_),
    .B(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__a22o_1 _17011_ (.A1(_09636_),
    .A2(_09753_),
    .B1(_09755_),
    .B2(_09623_),
    .X(_10033_));
 sky130_fd_sc_hd__o21bai_1 _17012_ (.A1(_09759_),
    .A2(_09764_),
    .B1_N(_09762_),
    .Y(_10034_));
 sky130_fd_sc_hd__nor2_1 _17013_ (.A(_08409_),
    .B(_09497_),
    .Y(_10035_));
 sky130_fd_sc_hd__xnor2_1 _17014_ (.A(_09753_),
    .B(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__nor2_1 _17015_ (.A(_08442_),
    .B(_09495_),
    .Y(_10037_));
 sky130_fd_sc_hd__xnor2_1 _17016_ (.A(_10036_),
    .B(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__nand2_1 _17017_ (.A(_10034_),
    .B(_10038_),
    .Y(_10039_));
 sky130_fd_sc_hd__or2_1 _17018_ (.A(_10034_),
    .B(_10038_),
    .X(_10040_));
 sky130_fd_sc_hd__nand2_1 _17019_ (.A(_10039_),
    .B(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__xnor2_1 _17020_ (.A(_10033_),
    .B(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__nor2_1 _17021_ (.A(_09751_),
    .B(_09630_),
    .Y(_10043_));
 sky130_fd_sc_hd__and3_1 _17022_ (.A(_08260_),
    .B(_09760_),
    .C(_09761_),
    .X(_10044_));
 sky130_fd_sc_hd__a2bb2o_1 _17023_ (.A1_N(_08362_),
    .A2_N(_09639_),
    .B1(_09760_),
    .B2(_08269_),
    .X(_10045_));
 sky130_fd_sc_hd__and2b_1 _17024_ (.A_N(_10044_),
    .B(_10045_),
    .X(_10046_));
 sky130_fd_sc_hd__xor2_1 _17025_ (.A(_10043_),
    .B(_10046_),
    .X(_10047_));
 sky130_fd_sc_hd__o32a_1 _17026_ (.A1(_08830_),
    .A2(_09773_),
    .A3(_09771_),
    .B1(_09770_),
    .B2(_06270_),
    .X(_10048_));
 sky130_fd_sc_hd__nand2_1 _17027_ (.A(\rbzero.wall_tracer.stepDistX[10] ),
    .B(_08629_),
    .Y(_10049_));
 sky130_fd_sc_hd__nand2_1 _17028_ (.A(\rbzero.wall_tracer.stepDistY[10] ),
    .B(_08304_),
    .Y(_10050_));
 sky130_fd_sc_hd__a21o_1 _17029_ (.A1(_09769_),
    .A2(_10050_),
    .B1(_08629_),
    .X(_10051_));
 sky130_fd_sc_hd__a21o_1 _17030_ (.A1(_10049_),
    .A2(_10051_),
    .B1(_08941_),
    .X(_10052_));
 sky130_fd_sc_hd__a21o_1 _17031_ (.A1(_09772_),
    .A2(_09644_),
    .B1(_08629_),
    .X(_10053_));
 sky130_fd_sc_hd__nand2_1 _17032_ (.A(\rbzero.wall_tracer.stepDistX[9] ),
    .B(_08629_),
    .Y(_10054_));
 sky130_fd_sc_hd__a21oi_1 _17033_ (.A1(_10053_),
    .A2(_10054_),
    .B1(_08941_),
    .Y(_10055_));
 sky130_fd_sc_hd__or3_1 _17034_ (.A(_08314_),
    .B(_08298_),
    .C(_09769_),
    .X(_10056_));
 sky130_fd_sc_hd__mux2_1 _17035_ (.A0(_08599_),
    .A1(_10056_),
    .S(_09770_),
    .X(_10057_));
 sky130_fd_sc_hd__mux2_1 _17036_ (.A0(_10052_),
    .A1(_10055_),
    .S(_10057_),
    .X(_10058_));
 sky130_fd_sc_hd__xnor2_1 _17037_ (.A(_10048_),
    .B(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__xnor2_1 _17038_ (.A(_10047_),
    .B(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__or2b_1 _17039_ (.A(_09775_),
    .B_N(_09777_),
    .X(_10061_));
 sky130_fd_sc_hd__a21bo_1 _17040_ (.A1(_09767_),
    .A2(_09778_),
    .B1_N(_10061_),
    .X(_10062_));
 sky130_fd_sc_hd__xnor2_1 _17041_ (.A(_10060_),
    .B(_10062_),
    .Y(_10063_));
 sky130_fd_sc_hd__xnor2_1 _17042_ (.A(_10042_),
    .B(_10063_),
    .Y(_10064_));
 sky130_fd_sc_hd__or2b_1 _17043_ (.A(_09779_),
    .B_N(_09781_),
    .X(_10065_));
 sky130_fd_sc_hd__a21bo_1 _17044_ (.A1(_09758_),
    .A2(_09782_),
    .B1_N(_10065_),
    .X(_10066_));
 sky130_fd_sc_hd__xnor2_1 _17045_ (.A(_10064_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__xnor2_1 _17046_ (.A(_10032_),
    .B(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__and2b_1 _17047_ (.A_N(_09783_),
    .B(_09785_),
    .X(_10069_));
 sky130_fd_sc_hd__a21oi_1 _17048_ (.A1(_09749_),
    .A2(_09786_),
    .B1(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__or2_1 _17049_ (.A(_10068_),
    .B(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__nand2_1 _17050_ (.A(_10068_),
    .B(_10070_),
    .Y(_10072_));
 sky130_fd_sc_hd__and2_1 _17051_ (.A(_10071_),
    .B(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__xnor2_1 _17052_ (.A(_10008_),
    .B(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__or2b_1 _17053_ (.A(_09787_),
    .B_N(_09788_),
    .X(_10075_));
 sky130_fd_sc_hd__a21boi_1 _17054_ (.A1(_09728_),
    .A2(_09789_),
    .B1_N(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__xor2_1 _17055_ (.A(_10074_),
    .B(_10076_),
    .X(_10077_));
 sky130_fd_sc_hd__nand2_1 _17056_ (.A(_09973_),
    .B(_10077_),
    .Y(_10078_));
 sky130_fd_sc_hd__or2_1 _17057_ (.A(_09973_),
    .B(_10077_),
    .X(_10079_));
 sky130_fd_sc_hd__nand2_1 _17058_ (.A(_10078_),
    .B(_10079_),
    .Y(_10080_));
 sky130_fd_sc_hd__o2bb2a_1 _17059_ (.A1_N(_09693_),
    .A2_N(_09792_),
    .B1(_09791_),
    .B2(_09790_),
    .X(_10081_));
 sky130_fd_sc_hd__xor2_1 _17060_ (.A(_10080_),
    .B(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__nand2_1 _17061_ (.A(_09968_),
    .B(_10082_),
    .Y(_10083_));
 sky130_fd_sc_hd__or2_1 _17062_ (.A(_09968_),
    .B(_10082_),
    .X(_10084_));
 sky130_fd_sc_hd__and2_1 _17063_ (.A(_10083_),
    .B(_10084_),
    .X(_10085_));
 sky130_fd_sc_hd__nand2_1 _17064_ (.A(_09967_),
    .B(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__or2_1 _17065_ (.A(_09967_),
    .B(_10085_),
    .X(_10087_));
 sky130_fd_sc_hd__nand2_2 _17066_ (.A(_10086_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__inv_2 _17067_ (.A(_09796_),
    .Y(_10089_));
 sky130_fd_sc_hd__a21o_1 _17068_ (.A1(_09685_),
    .A2(_09670_),
    .B1(_09795_),
    .X(_10090_));
 sky130_fd_sc_hd__o31a_2 _17069_ (.A1(_09560_),
    .A2(_09672_),
    .A3(_10089_),
    .B1(_10090_),
    .X(_10091_));
 sky130_fd_sc_hd__xor2_4 _17070_ (.A(_10088_),
    .B(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__nand2_1 _17071_ (.A(_08156_),
    .B(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__or2_1 _17072_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .X(_10094_));
 sky130_fd_sc_hd__nand2_1 _17073_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_10095_));
 sky130_fd_sc_hd__a211oi_1 _17074_ (.A1(_10094_),
    .A2(_10095_),
    .B1(_09959_),
    .C1(_09962_),
    .Y(_10096_));
 sky130_fd_sc_hd__o211a_1 _17075_ (.A1(_09959_),
    .A2(_09962_),
    .B1(_10094_),
    .C1(_10095_),
    .X(_10097_));
 sky130_fd_sc_hd__o31a_1 _17076_ (.A1(_08156_),
    .A2(_10096_),
    .A3(_10097_),
    .B1(_09883_),
    .X(_10098_));
 sky130_fd_sc_hd__o2bb2a_1 _17077_ (.A1_N(_10093_),
    .A2_N(_10098_),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_09884_),
    .X(_00539_));
 sky130_fd_sc_hd__or2_1 _17078_ (.A(_10080_),
    .B(_10081_),
    .X(_10099_));
 sky130_fd_sc_hd__or2b_1 _17079_ (.A(_10007_),
    .B_N(_09974_),
    .X(_10100_));
 sky130_fd_sc_hd__a21oi_1 _17080_ (.A1(_09985_),
    .A2(_09987_),
    .B1(_09984_),
    .Y(_10101_));
 sky130_fd_sc_hd__a21oi_1 _17081_ (.A1(_10005_),
    .A2(_10100_),
    .B1(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__and3_1 _17082_ (.A(_10005_),
    .B(_10100_),
    .C(_10101_),
    .X(_10103_));
 sky130_fd_sc_hd__nor2_1 _17083_ (.A(_10102_),
    .B(_10103_),
    .Y(_10104_));
 sky130_fd_sc_hd__nand2_1 _17084_ (.A(_10008_),
    .B(_10073_),
    .Y(_10105_));
 sky130_fd_sc_hd__o21ai_1 _17085_ (.A1(_09999_),
    .A2(_10000_),
    .B1(_10002_),
    .Y(_10106_));
 sky130_fd_sc_hd__or2b_1 _17086_ (.A(_10030_),
    .B_N(_10011_),
    .X(_10107_));
 sky130_fd_sc_hd__or2b_1 _17087_ (.A(_10031_),
    .B_N(_10009_),
    .X(_10108_));
 sky130_fd_sc_hd__nand2_1 _17088_ (.A(_10107_),
    .B(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__o22a_1 _17089_ (.A1(_09228_),
    .A2(_09313_),
    .B1(_09441_),
    .B2(_09094_),
    .X(_10110_));
 sky130_fd_sc_hd__or2_1 _17090_ (.A(_08831_),
    .B(_09440_),
    .X(_10111_));
 sky130_fd_sc_hd__or3_1 _17091_ (.A(_09094_),
    .B(_09313_),
    .C(_10111_),
    .X(_10112_));
 sky130_fd_sc_hd__and2b_1 _17092_ (.A_N(_10110_),
    .B(_10112_),
    .X(_10113_));
 sky130_fd_sc_hd__nor2_1 _17093_ (.A(_08959_),
    .B(_09571_),
    .Y(_10114_));
 sky130_fd_sc_hd__xnor2_1 _17094_ (.A(_10113_),
    .B(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__a21oi_1 _17095_ (.A1(_09697_),
    .A2(_09977_),
    .B1(_09980_),
    .Y(_10116_));
 sky130_fd_sc_hd__xor2_1 _17096_ (.A(_10115_),
    .B(_10116_),
    .X(_10117_));
 sky130_fd_sc_hd__and2_1 _17097_ (.A(_08567_),
    .B(_09691_),
    .X(_10118_));
 sky130_fd_sc_hd__xor2_1 _17098_ (.A(_10117_),
    .B(_10118_),
    .X(_10119_));
 sky130_fd_sc_hd__o31ai_2 _17099_ (.A1(_09228_),
    .A2(_09213_),
    .A3(_09990_),
    .B1(_09991_),
    .Y(_10120_));
 sky130_fd_sc_hd__nand2_1 _17100_ (.A(_09734_),
    .B(_10014_),
    .Y(_10121_));
 sky130_fd_sc_hd__nand2_1 _17101_ (.A(_10121_),
    .B(_10017_),
    .Y(_10122_));
 sky130_fd_sc_hd__o22ai_1 _17102_ (.A1(_08661_),
    .A2(_09070_),
    .B1(_09159_),
    .B2(_09466_),
    .Y(_10123_));
 sky130_fd_sc_hd__or3_1 _17103_ (.A(_08661_),
    .B(_09159_),
    .C(_09712_),
    .X(_10124_));
 sky130_fd_sc_hd__nand2_1 _17104_ (.A(_10123_),
    .B(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__nor2_1 _17105_ (.A(_09347_),
    .B(_09213_),
    .Y(_10126_));
 sky130_fd_sc_hd__xor2_1 _17106_ (.A(_10125_),
    .B(_10126_),
    .X(_10127_));
 sky130_fd_sc_hd__xnor2_1 _17107_ (.A(_10122_),
    .B(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__xnor2_1 _17108_ (.A(_10120_),
    .B(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__a21oi_1 _17109_ (.A1(_09989_),
    .A2(_09998_),
    .B1(_09996_),
    .Y(_10130_));
 sky130_fd_sc_hd__nor2_1 _17110_ (.A(_10129_),
    .B(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__and2_1 _17111_ (.A(_10129_),
    .B(_10130_),
    .X(_10132_));
 sky130_fd_sc_hd__nor2_1 _17112_ (.A(_10131_),
    .B(_10132_),
    .Y(_10133_));
 sky130_fd_sc_hd__xor2_1 _17113_ (.A(_10119_),
    .B(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__xnor2_1 _17114_ (.A(_10109_),
    .B(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__xnor2_1 _17115_ (.A(_10106_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__a21o_1 _17116_ (.A1(_10019_),
    .A2(_10029_),
    .B1(_10027_),
    .X(_10137_));
 sky130_fd_sc_hd__a21bo_1 _17117_ (.A1(_10033_),
    .A2(_10040_),
    .B1_N(_10039_),
    .X(_10138_));
 sky130_fd_sc_hd__nand2_1 _17118_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08321_),
    .Y(_10139_));
 sky130_fd_sc_hd__nand2_2 _17119_ (.A(_06340_),
    .B(_08228_),
    .Y(_10140_));
 sky130_fd_sc_hd__nor2_1 _17120_ (.A(_10139_),
    .B(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__xnor2_1 _17121_ (.A(_10014_),
    .B(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__or3_1 _17122_ (.A(_08293_),
    .B(_08573_),
    .C(_10142_),
    .X(_10143_));
 sky130_fd_sc_hd__clkbuf_4 _17123_ (.A(_08293_),
    .X(_10144_));
 sky130_fd_sc_hd__o21ai_1 _17124_ (.A1(_10144_),
    .A2(_09072_),
    .B1(_10142_),
    .Y(_10145_));
 sky130_fd_sc_hd__and2_1 _17125_ (.A(_10143_),
    .B(_10145_),
    .X(_10146_));
 sky130_fd_sc_hd__nor2_1 _17126_ (.A(_08559_),
    .B(_09126_),
    .Y(_10147_));
 sky130_fd_sc_hd__nor2_1 _17127_ (.A(_08808_),
    .B(_09131_),
    .Y(_10148_));
 sky130_fd_sc_hd__xnor2_1 _17128_ (.A(_10147_),
    .B(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__or2_1 _17129_ (.A(_08551_),
    .B(_08307_),
    .X(_10150_));
 sky130_fd_sc_hd__xnor2_1 _17130_ (.A(_10149_),
    .B(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__o31a_1 _17131_ (.A1(_08583_),
    .A2(_08307_),
    .A3(_09737_),
    .B1(_10023_),
    .X(_10152_));
 sky130_fd_sc_hd__nor2_1 _17132_ (.A(_10151_),
    .B(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__nand2_1 _17133_ (.A(_10151_),
    .B(_10152_),
    .Y(_10154_));
 sky130_fd_sc_hd__and2b_1 _17134_ (.A_N(_10153_),
    .B(_10154_),
    .X(_10155_));
 sky130_fd_sc_hd__xor2_1 _17135_ (.A(_10146_),
    .B(_10155_),
    .X(_10156_));
 sky130_fd_sc_hd__xnor2_1 _17136_ (.A(_10138_),
    .B(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__xnor2_1 _17137_ (.A(_10137_),
    .B(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__buf_2 _17138_ (.A(_08442_),
    .X(_10159_));
 sky130_fd_sc_hd__or3_1 _17139_ (.A(_10159_),
    .B(_09495_),
    .C(_10036_),
    .X(_10160_));
 sky130_fd_sc_hd__a21bo_1 _17140_ (.A1(_09753_),
    .A2(_10035_),
    .B1_N(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__a21o_1 _17141_ (.A1(_10043_),
    .A2(_10045_),
    .B1(_10044_),
    .X(_10162_));
 sky130_fd_sc_hd__clkbuf_4 _17142_ (.A(_09383_),
    .X(_10163_));
 sky130_fd_sc_hd__a21oi_1 _17143_ (.A1(_10163_),
    .A2(_09384_),
    .B1(_09371_),
    .Y(_10164_));
 sky130_fd_sc_hd__a21oi_2 _17144_ (.A1(_09502_),
    .A2(_09503_),
    .B1(_09372_),
    .Y(_10165_));
 sky130_fd_sc_hd__xnor2_1 _17145_ (.A(_10164_),
    .B(_10165_),
    .Y(_10166_));
 sky130_fd_sc_hd__nor2_1 _17146_ (.A(_08442_),
    .B(_09497_),
    .Y(_10167_));
 sky130_fd_sc_hd__xnor2_1 _17147_ (.A(_10166_),
    .B(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__and2_1 _17148_ (.A(_10162_),
    .B(_10168_),
    .X(_10169_));
 sky130_fd_sc_hd__or2_1 _17149_ (.A(_10162_),
    .B(_10168_),
    .X(_10170_));
 sky130_fd_sc_hd__or2b_1 _17150_ (.A(_10169_),
    .B_N(_10170_),
    .X(_10171_));
 sky130_fd_sc_hd__xnor2_1 _17151_ (.A(_10161_),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__buf_2 _17152_ (.A(_09639_),
    .X(_10173_));
 sky130_fd_sc_hd__nor2_1 _17153_ (.A(_09751_),
    .B(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__nand2_1 _17154_ (.A(_08260_),
    .B(_09763_),
    .Y(_10175_));
 sky130_fd_sc_hd__a21o_1 _17155_ (.A1(_10053_),
    .A2(_10054_),
    .B1(_08918_),
    .X(_10176_));
 sky130_fd_sc_hd__xnor2_1 _17156_ (.A(_10175_),
    .B(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__xnor2_1 _17157_ (.A(_10174_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand3_1 _17158_ (.A(_09770_),
    .B(_10056_),
    .C(_10052_),
    .Y(_10179_));
 sky130_fd_sc_hd__or3_2 _17159_ (.A(_09021_),
    .B(_09770_),
    .C(_10052_),
    .X(_10180_));
 sky130_fd_sc_hd__and2_1 _17160_ (.A(_10179_),
    .B(_10180_),
    .X(_10181_));
 sky130_fd_sc_hd__buf_2 _17161_ (.A(_10181_),
    .X(_10182_));
 sky130_fd_sc_hd__xnor2_1 _17162_ (.A(_10178_),
    .B(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__and2b_1 _17163_ (.A_N(_10048_),
    .B(_10058_),
    .X(_10184_));
 sky130_fd_sc_hd__a21oi_2 _17164_ (.A1(_10047_),
    .A2(_10059_),
    .B1(_10184_),
    .Y(_10185_));
 sky130_fd_sc_hd__xor2_1 _17165_ (.A(_10183_),
    .B(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__xnor2_1 _17166_ (.A(_10172_),
    .B(_10186_),
    .Y(_10187_));
 sky130_fd_sc_hd__or2b_1 _17167_ (.A(_10060_),
    .B_N(_10062_),
    .X(_10188_));
 sky130_fd_sc_hd__a21bo_1 _17168_ (.A1(_10042_),
    .A2(_10063_),
    .B1_N(_10188_),
    .X(_10189_));
 sky130_fd_sc_hd__xnor2_1 _17169_ (.A(_10187_),
    .B(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__xnor2_1 _17170_ (.A(_10158_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__and2b_1 _17171_ (.A_N(_10064_),
    .B(_10066_),
    .X(_10192_));
 sky130_fd_sc_hd__a21oi_1 _17172_ (.A1(_10032_),
    .A2(_10067_),
    .B1(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__nor2_1 _17173_ (.A(_10191_),
    .B(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__and2_1 _17174_ (.A(_10191_),
    .B(_10193_),
    .X(_10195_));
 sky130_fd_sc_hd__nor2_1 _17175_ (.A(_10194_),
    .B(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__xnor2_1 _17176_ (.A(_10136_),
    .B(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__a21oi_1 _17177_ (.A1(_10071_),
    .A2(_10105_),
    .B1(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__and3_1 _17178_ (.A(_10071_),
    .B(_10105_),
    .C(_10197_),
    .X(_10199_));
 sky130_fd_sc_hd__nor2_1 _17179_ (.A(_10198_),
    .B(_10199_),
    .Y(_10200_));
 sky130_fd_sc_hd__xnor2_1 _17180_ (.A(_10104_),
    .B(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__o21a_1 _17181_ (.A1(_10074_),
    .A2(_10076_),
    .B1(_10078_),
    .X(_10202_));
 sky130_fd_sc_hd__nor2_1 _17182_ (.A(_10201_),
    .B(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__and2_1 _17183_ (.A(_10201_),
    .B(_10202_),
    .X(_10204_));
 sky130_fd_sc_hd__nor2_1 _17184_ (.A(_10203_),
    .B(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__xnor2_2 _17185_ (.A(_09971_),
    .B(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__a21oi_1 _17186_ (.A1(_10099_),
    .A2(_10083_),
    .B1(_10206_),
    .Y(_10207_));
 sky130_fd_sc_hd__and3_1 _17187_ (.A(_10099_),
    .B(_10083_),
    .C(_10206_),
    .X(_10208_));
 sky130_fd_sc_hd__or2_2 _17188_ (.A(_10207_),
    .B(_10208_),
    .X(_10209_));
 sky130_fd_sc_hd__o21ai_2 _17189_ (.A1(_10088_),
    .A2(_10091_),
    .B1(_10086_),
    .Y(_10210_));
 sky130_fd_sc_hd__xnor2_4 _17190_ (.A(_10209_),
    .B(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__nand2_1 _17191_ (.A(_09905_),
    .B(_10211_),
    .Y(_10212_));
 sky130_fd_sc_hd__nand2_1 _17192_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_10213_));
 sky130_fd_sc_hd__or2_1 _17193_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_10214_));
 sky130_fd_sc_hd__a21o_1 _17194_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(\rbzero.wall_tracer.stepDistX[0] ),
    .B1(_10097_),
    .X(_10215_));
 sky130_fd_sc_hd__and3_1 _17195_ (.A(_10213_),
    .B(_10214_),
    .C(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__a21o_1 _17196_ (.A1(_10213_),
    .A2(_10214_),
    .B1(_10215_),
    .X(_10217_));
 sky130_fd_sc_hd__or3b_1 _17197_ (.A(_06163_),
    .B(_10216_),
    .C_N(_10217_),
    .X(_10218_));
 sky130_fd_sc_hd__nand2_1 _17198_ (.A(_10212_),
    .B(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__mux2_1 _17199_ (.A0(\rbzero.wall_tracer.trackDistX[1] ),
    .A1(_10219_),
    .S(_09917_),
    .X(_10220_));
 sky130_fd_sc_hd__clkbuf_1 _17200_ (.A(_10220_),
    .X(_00540_));
 sky130_fd_sc_hd__nand2_1 _17201_ (.A(_10109_),
    .B(_10134_),
    .Y(_10221_));
 sky130_fd_sc_hd__or2b_1 _17202_ (.A(_10135_),
    .B_N(_10106_),
    .X(_10222_));
 sky130_fd_sc_hd__o2bb2a_1 _17203_ (.A1_N(_10117_),
    .A2_N(_10118_),
    .B1(_10115_),
    .B2(_10116_),
    .X(_10223_));
 sky130_fd_sc_hd__a21oi_1 _17204_ (.A1(_10221_),
    .A2(_10222_),
    .B1(_10223_),
    .Y(_10224_));
 sky130_fd_sc_hd__and3_1 _17205_ (.A(_10221_),
    .B(_10222_),
    .C(_10223_),
    .X(_10225_));
 sky130_fd_sc_hd__nor2_1 _17206_ (.A(_10224_),
    .B(_10225_),
    .Y(_10226_));
 sky130_fd_sc_hd__a21o_1 _17207_ (.A1(_10119_),
    .A2(_10133_),
    .B1(_10131_),
    .X(_10227_));
 sky130_fd_sc_hd__or2b_1 _17208_ (.A(_10157_),
    .B_N(_10137_),
    .X(_10228_));
 sky130_fd_sc_hd__a21bo_1 _17209_ (.A1(_10138_),
    .A2(_10156_),
    .B1_N(_10228_),
    .X(_10229_));
 sky130_fd_sc_hd__or2_1 _17210_ (.A(_09347_),
    .B(_09440_),
    .X(_10230_));
 sky130_fd_sc_hd__o21ai_1 _17211_ (.A1(_09347_),
    .A2(_09314_),
    .B1(_10111_),
    .Y(_10231_));
 sky130_fd_sc_hd__o31a_1 _17212_ (.A1(_09228_),
    .A2(_09314_),
    .A3(_10230_),
    .B1(_10231_),
    .X(_10232_));
 sky130_fd_sc_hd__nor2_1 _17213_ (.A(_09094_),
    .B(_09571_),
    .Y(_10233_));
 sky130_fd_sc_hd__nand2_1 _17214_ (.A(_10232_),
    .B(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__or2_1 _17215_ (.A(_10232_),
    .B(_10233_),
    .X(_10235_));
 sky130_fd_sc_hd__nand2_1 _17216_ (.A(_10234_),
    .B(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__o31a_1 _17217_ (.A1(_08959_),
    .A2(_09706_),
    .A3(_10110_),
    .B1(_10112_),
    .X(_10237_));
 sky130_fd_sc_hd__xor2_1 _17218_ (.A(_10236_),
    .B(_10237_),
    .X(_10238_));
 sky130_fd_sc_hd__and2_1 _17219_ (.A(_08959_),
    .B(_09691_),
    .X(_10239_));
 sky130_fd_sc_hd__xor2_1 _17220_ (.A(_10238_),
    .B(_10239_),
    .X(_10240_));
 sky130_fd_sc_hd__a21bo_1 _17221_ (.A1(_10123_),
    .A2(_10126_),
    .B1_N(_10124_),
    .X(_10241_));
 sky130_fd_sc_hd__o22ai_1 _17222_ (.A1(_08293_),
    .A2(_09070_),
    .B1(_09159_),
    .B2(_10012_),
    .Y(_10242_));
 sky130_fd_sc_hd__or4_1 _17223_ (.A(_08661_),
    .B(_08293_),
    .C(_09070_),
    .D(_09159_),
    .X(_10243_));
 sky130_fd_sc_hd__nand2_1 _17224_ (.A(_10242_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__nor2_1 _17225_ (.A(_09466_),
    .B(_09213_),
    .Y(_10245_));
 sky130_fd_sc_hd__xor2_1 _17226_ (.A(_10244_),
    .B(_10245_),
    .X(_10246_));
 sky130_fd_sc_hd__a21bo_1 _17227_ (.A1(_10014_),
    .A2(_10141_),
    .B1_N(_10143_),
    .X(_10247_));
 sky130_fd_sc_hd__and2b_1 _17228_ (.A_N(_10246_),
    .B(_10247_),
    .X(_10248_));
 sky130_fd_sc_hd__and2b_1 _17229_ (.A_N(_10247_),
    .B(_10246_),
    .X(_10249_));
 sky130_fd_sc_hd__nor2_1 _17230_ (.A(_10248_),
    .B(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__xnor2_1 _17231_ (.A(_10241_),
    .B(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__a21oi_1 _17232_ (.A1(_10121_),
    .A2(_10017_),
    .B1(_10127_),
    .Y(_10252_));
 sky130_fd_sc_hd__a21oi_1 _17233_ (.A1(_10120_),
    .A2(_10128_),
    .B1(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__nor2_1 _17234_ (.A(_10251_),
    .B(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__and2_1 _17235_ (.A(_10251_),
    .B(_10253_),
    .X(_10255_));
 sky130_fd_sc_hd__nor2_1 _17236_ (.A(_10254_),
    .B(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__xor2_1 _17237_ (.A(_10240_),
    .B(_10256_),
    .X(_10257_));
 sky130_fd_sc_hd__xnor2_1 _17238_ (.A(_10229_),
    .B(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__xnor2_1 _17239_ (.A(_10227_),
    .B(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__a21o_1 _17240_ (.A1(_10146_),
    .A2(_10154_),
    .B1(_10153_),
    .X(_10260_));
 sky130_fd_sc_hd__a21o_1 _17241_ (.A1(_10161_),
    .A2(_10170_),
    .B1(_10169_),
    .X(_10261_));
 sky130_fd_sc_hd__buf_2 _17242_ (.A(_10013_),
    .X(_10262_));
 sky130_fd_sc_hd__nor2_1 _17243_ (.A(_08495_),
    .B(_08303_),
    .Y(_10263_));
 sky130_fd_sc_hd__a31o_1 _17244_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_08496_),
    .A3(_08228_),
    .B1(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__buf_2 _17245_ (.A(_10139_),
    .X(_10265_));
 sky130_fd_sc_hd__nor2_1 _17246_ (.A(_08506_),
    .B(_08303_),
    .Y(_10266_));
 sky130_fd_sc_hd__or3b_1 _17247_ (.A(_10265_),
    .B(_10140_),
    .C_N(_10266_),
    .X(_10267_));
 sky130_fd_sc_hd__nand2_1 _17248_ (.A(_10264_),
    .B(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__or3_1 _17249_ (.A(_10262_),
    .B(_09072_),
    .C(_10268_),
    .X(_10269_));
 sky130_fd_sc_hd__o21ai_1 _17250_ (.A1(_10262_),
    .A2(_09072_),
    .B1(_10268_),
    .Y(_10270_));
 sky130_fd_sc_hd__and2_1 _17251_ (.A(_10269_),
    .B(_10270_),
    .X(_10271_));
 sky130_fd_sc_hd__or2_1 _17252_ (.A(_08559_),
    .B(_09497_),
    .X(_10272_));
 sky130_fd_sc_hd__o22ai_1 _17253_ (.A1(_08559_),
    .A2(_09495_),
    .B1(_09497_),
    .B2(_08808_),
    .Y(_10273_));
 sky130_fd_sc_hd__o31ai_1 _17254_ (.A1(_08808_),
    .A2(_09495_),
    .A3(_10272_),
    .B1(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__nor2_1 _17255_ (.A(_09358_),
    .B(_09126_),
    .Y(_10275_));
 sky130_fd_sc_hd__xor2_1 _17256_ (.A(_10274_),
    .B(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__nand2_1 _17257_ (.A(_10147_),
    .B(_10148_),
    .Y(_10277_));
 sky130_fd_sc_hd__o31a_1 _17258_ (.A1(_09358_),
    .A2(_08307_),
    .A3(_10149_),
    .B1(_10277_),
    .X(_10278_));
 sky130_fd_sc_hd__nor2_1 _17259_ (.A(_10276_),
    .B(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__nand2_1 _17260_ (.A(_10276_),
    .B(_10278_),
    .Y(_10280_));
 sky130_fd_sc_hd__and2b_1 _17261_ (.A_N(_10279_),
    .B(_10280_),
    .X(_10281_));
 sky130_fd_sc_hd__xor2_1 _17262_ (.A(_10271_),
    .B(_10281_),
    .X(_10282_));
 sky130_fd_sc_hd__xnor2_1 _17263_ (.A(_10261_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__xnor2_1 _17264_ (.A(_10260_),
    .B(_10283_),
    .Y(_10284_));
 sky130_fd_sc_hd__or3_1 _17265_ (.A(_10159_),
    .B(_09497_),
    .C(_10166_),
    .X(_10285_));
 sky130_fd_sc_hd__a21bo_1 _17266_ (.A1(_10164_),
    .A2(_10165_),
    .B1_N(_10285_),
    .X(_10286_));
 sky130_fd_sc_hd__or2_1 _17267_ (.A(_10175_),
    .B(_10176_),
    .X(_10287_));
 sky130_fd_sc_hd__o31a_1 _17268_ (.A1(_09751_),
    .A2(_10173_),
    .A3(_10177_),
    .B1(_10287_),
    .X(_10288_));
 sky130_fd_sc_hd__or3b_1 _17269_ (.A(_09371_),
    .B(_10173_),
    .C_N(_10165_),
    .X(_10289_));
 sky130_fd_sc_hd__o22ai_1 _17270_ (.A1(_09371_),
    .A2(_09630_),
    .B1(_10173_),
    .B2(_09372_),
    .Y(_10290_));
 sky130_fd_sc_hd__nor2_1 _17271_ (.A(_08442_),
    .B(_09633_),
    .Y(_10291_));
 sky130_fd_sc_hd__and3_1 _17272_ (.A(_10289_),
    .B(_10290_),
    .C(_10291_),
    .X(_10292_));
 sky130_fd_sc_hd__a21oi_1 _17273_ (.A1(_10289_),
    .A2(_10290_),
    .B1(_10291_),
    .Y(_10293_));
 sky130_fd_sc_hd__or2_1 _17274_ (.A(_10292_),
    .B(_10293_),
    .X(_10294_));
 sky130_fd_sc_hd__xor2_1 _17275_ (.A(_10288_),
    .B(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__xor2_1 _17276_ (.A(_10286_),
    .B(_10295_),
    .X(_10296_));
 sky130_fd_sc_hd__and2b_1 _17277_ (.A_N(_09751_),
    .B(_09763_),
    .X(_10297_));
 sky130_fd_sc_hd__a21oi_1 _17278_ (.A1(_10053_),
    .A2(_10054_),
    .B1(_08362_),
    .Y(_10298_));
 sky130_fd_sc_hd__a21o_1 _17279_ (.A1(_10049_),
    .A2(_10051_),
    .B1(_08918_),
    .X(_10299_));
 sky130_fd_sc_hd__xnor2_1 _17280_ (.A(_10298_),
    .B(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__xor2_1 _17281_ (.A(_10297_),
    .B(_10300_),
    .X(_10301_));
 sky130_fd_sc_hd__xnor2_1 _17282_ (.A(_10182_),
    .B(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__a21bo_1 _17283_ (.A1(_10178_),
    .A2(_10182_),
    .B1_N(_10180_),
    .X(_10303_));
 sky130_fd_sc_hd__xnor2_1 _17284_ (.A(_10302_),
    .B(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__xnor2_1 _17285_ (.A(_10296_),
    .B(_10304_),
    .Y(_10305_));
 sky130_fd_sc_hd__nor2_1 _17286_ (.A(_10183_),
    .B(_10185_),
    .Y(_10306_));
 sky130_fd_sc_hd__a21o_1 _17287_ (.A1(_10172_),
    .A2(_10186_),
    .B1(_10306_),
    .X(_10307_));
 sky130_fd_sc_hd__xnor2_1 _17288_ (.A(_10305_),
    .B(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__xnor2_1 _17289_ (.A(_10284_),
    .B(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__and2b_1 _17290_ (.A_N(_10187_),
    .B(_10189_),
    .X(_10310_));
 sky130_fd_sc_hd__a21oi_1 _17291_ (.A1(_10158_),
    .A2(_10190_),
    .B1(_10310_),
    .Y(_10311_));
 sky130_fd_sc_hd__nor2_1 _17292_ (.A(_10309_),
    .B(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__and2_1 _17293_ (.A(_10309_),
    .B(_10311_),
    .X(_10313_));
 sky130_fd_sc_hd__nor2_1 _17294_ (.A(_10312_),
    .B(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__xnor2_1 _17295_ (.A(_10259_),
    .B(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__a21oi_1 _17296_ (.A1(_10136_),
    .A2(_10196_),
    .B1(_10194_),
    .Y(_10316_));
 sky130_fd_sc_hd__nor2_1 _17297_ (.A(_10315_),
    .B(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__and2_1 _17298_ (.A(_10315_),
    .B(_10316_),
    .X(_10318_));
 sky130_fd_sc_hd__nor2_1 _17299_ (.A(_10317_),
    .B(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__xnor2_1 _17300_ (.A(_10226_),
    .B(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__a21oi_1 _17301_ (.A1(_10104_),
    .A2(_10200_),
    .B1(_10198_),
    .Y(_10321_));
 sky130_fd_sc_hd__xor2_1 _17302_ (.A(_10320_),
    .B(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__nand2_1 _17303_ (.A(_10102_),
    .B(_10322_),
    .Y(_10323_));
 sky130_fd_sc_hd__or2_1 _17304_ (.A(_10102_),
    .B(_10322_),
    .X(_10324_));
 sky130_fd_sc_hd__nand2_1 _17305_ (.A(_10323_),
    .B(_10324_),
    .Y(_10325_));
 sky130_fd_sc_hd__a21oi_1 _17306_ (.A1(_09971_),
    .A2(_10205_),
    .B1(_10203_),
    .Y(_10326_));
 sky130_fd_sc_hd__or2_1 _17307_ (.A(_10325_),
    .B(_10326_),
    .X(_10327_));
 sky130_fd_sc_hd__nand2_1 _17308_ (.A(_10325_),
    .B(_10326_),
    .Y(_10328_));
 sky130_fd_sc_hd__and2_2 _17309_ (.A(_10327_),
    .B(_10328_),
    .X(_10329_));
 sky130_fd_sc_hd__a21o_1 _17310_ (.A1(_10099_),
    .A2(_10083_),
    .B1(_10206_),
    .X(_10330_));
 sky130_fd_sc_hd__a21o_1 _17311_ (.A1(_10086_),
    .A2(_10330_),
    .B1(_10208_),
    .X(_10331_));
 sky130_fd_sc_hd__o31a_4 _17312_ (.A1(_10088_),
    .A2(_10091_),
    .A3(_10209_),
    .B1(_10331_),
    .X(_10332_));
 sky130_fd_sc_hd__xnor2_4 _17313_ (.A(_10329_),
    .B(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__nand2_1 _17314_ (.A(_06162_),
    .B(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__inv_2 _17315_ (.A(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__nand2_1 _17316_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .Y(_10336_));
 sky130_fd_sc_hd__or2_1 _17317_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_10337_));
 sky130_fd_sc_hd__inv_2 _17318_ (.A(_10213_),
    .Y(_10338_));
 sky130_fd_sc_hd__a211o_1 _17319_ (.A1(_10336_),
    .A2(_10337_),
    .B1(_10338_),
    .C1(_10216_),
    .X(_10339_));
 sky130_fd_sc_hd__o211ai_2 _17320_ (.A1(_10338_),
    .A2(_10216_),
    .B1(_10336_),
    .C1(_10337_),
    .Y(_10340_));
 sky130_fd_sc_hd__a31o_1 _17321_ (.A1(_08195_),
    .A2(_10339_),
    .A3(_10340_),
    .B1(_09859_),
    .X(_10341_));
 sky130_fd_sc_hd__o22a_1 _17322_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_09883_),
    .B1(_10335_),
    .B2(_10341_),
    .X(_00541_));
 sky130_fd_sc_hd__or2_1 _17323_ (.A(_10320_),
    .B(_10321_),
    .X(_10342_));
 sky130_fd_sc_hd__nand2_1 _17324_ (.A(_10229_),
    .B(_10257_),
    .Y(_10343_));
 sky130_fd_sc_hd__or2b_1 _17325_ (.A(_10258_),
    .B_N(_10227_),
    .X(_10344_));
 sky130_fd_sc_hd__o2bb2a_1 _17326_ (.A1_N(_10238_),
    .A2_N(_10239_),
    .B1(_10236_),
    .B2(_10237_),
    .X(_10345_));
 sky130_fd_sc_hd__a21oi_1 _17327_ (.A1(_10343_),
    .A2(_10344_),
    .B1(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__and3_1 _17328_ (.A(_10343_),
    .B(_10344_),
    .C(_10345_),
    .X(_10347_));
 sky130_fd_sc_hd__nor2_1 _17329_ (.A(_10346_),
    .B(_10347_),
    .Y(_10348_));
 sky130_fd_sc_hd__a21o_1 _17330_ (.A1(_10240_),
    .A2(_10256_),
    .B1(_10254_),
    .X(_10349_));
 sky130_fd_sc_hd__or2b_1 _17331_ (.A(_10283_),
    .B_N(_10260_),
    .X(_10350_));
 sky130_fd_sc_hd__a21bo_1 _17332_ (.A1(_10261_),
    .A2(_10282_),
    .B1_N(_10350_),
    .X(_10351_));
 sky130_fd_sc_hd__nor2_1 _17333_ (.A(_09466_),
    .B(_09313_),
    .Y(_10352_));
 sky130_fd_sc_hd__xnor2_1 _17334_ (.A(_10230_),
    .B(_10352_),
    .Y(_10353_));
 sky130_fd_sc_hd__nor2_1 _17335_ (.A(_09228_),
    .B(_09571_),
    .Y(_10354_));
 sky130_fd_sc_hd__nand2_1 _17336_ (.A(_10353_),
    .B(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__or2_1 _17337_ (.A(_10353_),
    .B(_10354_),
    .X(_10356_));
 sky130_fd_sc_hd__nand2_1 _17338_ (.A(_10355_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__o31a_1 _17339_ (.A1(_09228_),
    .A2(_09314_),
    .A3(_10230_),
    .B1(_10234_),
    .X(_10358_));
 sky130_fd_sc_hd__xor2_1 _17340_ (.A(_10357_),
    .B(_10358_),
    .X(_10359_));
 sky130_fd_sc_hd__and2_1 _17341_ (.A(_09094_),
    .B(_09691_),
    .X(_10360_));
 sky130_fd_sc_hd__xor2_1 _17342_ (.A(_10359_),
    .B(_10360_),
    .X(_10361_));
 sky130_fd_sc_hd__a21bo_1 _17343_ (.A1(_10242_),
    .A2(_10245_),
    .B1_N(_10243_),
    .X(_10362_));
 sky130_fd_sc_hd__o22ai_1 _17344_ (.A1(_10262_),
    .A2(_09070_),
    .B1(_09159_),
    .B2(_08293_),
    .Y(_10363_));
 sky130_fd_sc_hd__or4_1 _17345_ (.A(_10262_),
    .B(_08293_),
    .C(_09070_),
    .D(_09159_),
    .X(_10364_));
 sky130_fd_sc_hd__nand2_1 _17346_ (.A(_10363_),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__nor2_1 _17347_ (.A(_08661_),
    .B(_09213_),
    .Y(_10366_));
 sky130_fd_sc_hd__xor2_1 _17348_ (.A(_10365_),
    .B(_10366_),
    .X(_10367_));
 sky130_fd_sc_hd__a21oi_1 _17349_ (.A1(_10267_),
    .A2(_10269_),
    .B1(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__and3_1 _17350_ (.A(_10267_),
    .B(_10269_),
    .C(_10367_),
    .X(_10369_));
 sky130_fd_sc_hd__nor2_1 _17351_ (.A(_10368_),
    .B(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__xnor2_1 _17352_ (.A(_10362_),
    .B(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__a21oi_1 _17353_ (.A1(_10241_),
    .A2(_10250_),
    .B1(_10248_),
    .Y(_10372_));
 sky130_fd_sc_hd__nor2_1 _17354_ (.A(_10371_),
    .B(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__and2_1 _17355_ (.A(_10371_),
    .B(_10372_),
    .X(_10374_));
 sky130_fd_sc_hd__nor2_1 _17356_ (.A(_10373_),
    .B(_10374_),
    .Y(_10375_));
 sky130_fd_sc_hd__xor2_1 _17357_ (.A(_10361_),
    .B(_10375_),
    .X(_10376_));
 sky130_fd_sc_hd__xnor2_1 _17358_ (.A(_10351_),
    .B(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__xnor2_1 _17359_ (.A(_10349_),
    .B(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__a21o_1 _17360_ (.A1(_10271_),
    .A2(_10280_),
    .B1(_10279_),
    .X(_10379_));
 sky130_fd_sc_hd__nor2_1 _17361_ (.A(_10288_),
    .B(_10294_),
    .Y(_10380_));
 sky130_fd_sc_hd__a21o_1 _17362_ (.A1(_10286_),
    .A2(_10295_),
    .B1(_10380_),
    .X(_10381_));
 sky130_fd_sc_hd__nand2_1 _17363_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08321_),
    .Y(_10382_));
 sky130_fd_sc_hd__nor2_1 _17364_ (.A(_06420_),
    .B(_08336_),
    .Y(_10383_));
 sky130_fd_sc_hd__xnor2_1 _17365_ (.A(_10266_),
    .B(_10383_),
    .Y(_10384_));
 sky130_fd_sc_hd__or3_1 _17366_ (.A(_10140_),
    .B(_10382_),
    .C(_10384_),
    .X(_10385_));
 sky130_fd_sc_hd__buf_2 _17367_ (.A(_10382_),
    .X(_10386_));
 sky130_fd_sc_hd__o21ai_1 _17368_ (.A1(_10140_),
    .A2(_10386_),
    .B1(_10384_),
    .Y(_10387_));
 sky130_fd_sc_hd__and2_1 _17369_ (.A(_10385_),
    .B(_10387_),
    .X(_10388_));
 sky130_fd_sc_hd__or3_1 _17370_ (.A(_08808_),
    .B(_09633_),
    .C(_10272_),
    .X(_10389_));
 sky130_fd_sc_hd__o21ai_1 _17371_ (.A1(_08809_),
    .A2(_09633_),
    .B1(_10272_),
    .Y(_10390_));
 sky130_fd_sc_hd__nand2_1 _17372_ (.A(_10389_),
    .B(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__nor2_1 _17373_ (.A(_09358_),
    .B(_09495_),
    .Y(_10392_));
 sky130_fd_sc_hd__xor2_1 _17374_ (.A(_10391_),
    .B(_10392_),
    .X(_10393_));
 sky130_fd_sc_hd__or3_1 _17375_ (.A(_09358_),
    .B(_09126_),
    .C(_10274_),
    .X(_10394_));
 sky130_fd_sc_hd__o31a_1 _17376_ (.A1(_08809_),
    .A2(_09495_),
    .A3(_10272_),
    .B1(_10394_),
    .X(_10395_));
 sky130_fd_sc_hd__xor2_1 _17377_ (.A(_10393_),
    .B(_10395_),
    .X(_10396_));
 sky130_fd_sc_hd__xnor2_1 _17378_ (.A(_10388_),
    .B(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__xor2_1 _17379_ (.A(_10381_),
    .B(_10397_),
    .X(_10398_));
 sky130_fd_sc_hd__xnor2_1 _17380_ (.A(_10379_),
    .B(_10398_),
    .Y(_10399_));
 sky130_fd_sc_hd__nor2_1 _17381_ (.A(_09371_),
    .B(_09639_),
    .Y(_10400_));
 sky130_fd_sc_hd__a21o_1 _17382_ (.A1(_10165_),
    .A2(_10400_),
    .B1(_10292_),
    .X(_10401_));
 sky130_fd_sc_hd__and2_1 _17383_ (.A(_10053_),
    .B(_10054_),
    .X(_10402_));
 sky130_fd_sc_hd__clkbuf_2 _17384_ (.A(_10402_),
    .X(_10403_));
 sky130_fd_sc_hd__a211o_2 _17385_ (.A1(_10049_),
    .A2(_10051_),
    .B1(_08272_),
    .C1(_08271_),
    .X(_10404_));
 sky130_fd_sc_hd__a2bb2o_1 _17386_ (.A1_N(_10403_),
    .A2_N(_10404_),
    .B1(_10300_),
    .B2(_10297_),
    .X(_10405_));
 sky130_fd_sc_hd__and2_1 _17387_ (.A(_08676_),
    .B(_09763_),
    .X(_10406_));
 sky130_fd_sc_hd__xnor2_1 _17388_ (.A(_10400_),
    .B(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__nor2_1 _17389_ (.A(_10159_),
    .B(_09630_),
    .Y(_10408_));
 sky130_fd_sc_hd__xnor2_1 _17390_ (.A(_10407_),
    .B(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__xnor2_1 _17391_ (.A(_10405_),
    .B(_10409_),
    .Y(_10410_));
 sky130_fd_sc_hd__xnor2_1 _17392_ (.A(_10401_),
    .B(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__nor2_1 _17393_ (.A(_08260_),
    .B(_08269_),
    .Y(_10412_));
 sky130_fd_sc_hd__and2_1 _17394_ (.A(_10049_),
    .B(_10051_),
    .X(_10413_));
 sky130_fd_sc_hd__buf_2 _17395_ (.A(_10413_),
    .X(_10414_));
 sky130_fd_sc_hd__or3b_1 _17396_ (.A(_10412_),
    .B(_10414_),
    .C_N(_10404_),
    .X(_10415_));
 sky130_fd_sc_hd__clkbuf_2 _17397_ (.A(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__nor2_1 _17398_ (.A(_09751_),
    .B(_10403_),
    .Y(_10417_));
 sky130_fd_sc_hd__xnor2_1 _17399_ (.A(_10416_),
    .B(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__xnor2_1 _17400_ (.A(_10182_),
    .B(_10418_),
    .Y(_10419_));
 sky130_fd_sc_hd__a21bo_1 _17401_ (.A1(_10182_),
    .A2(_10301_),
    .B1_N(_10180_),
    .X(_10420_));
 sky130_fd_sc_hd__xnor2_1 _17402_ (.A(_10419_),
    .B(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__xnor2_1 _17403_ (.A(_10411_),
    .B(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__or2b_1 _17404_ (.A(_10302_),
    .B_N(_10303_),
    .X(_10423_));
 sky130_fd_sc_hd__a21bo_1 _17405_ (.A1(_10296_),
    .A2(_10304_),
    .B1_N(_10423_),
    .X(_10424_));
 sky130_fd_sc_hd__xnor2_1 _17406_ (.A(_10422_),
    .B(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__xnor2_1 _17407_ (.A(_10399_),
    .B(_10425_),
    .Y(_10426_));
 sky130_fd_sc_hd__and2b_1 _17408_ (.A_N(_10305_),
    .B(_10307_),
    .X(_10427_));
 sky130_fd_sc_hd__a21oi_1 _17409_ (.A1(_10284_),
    .A2(_10308_),
    .B1(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__nor2_1 _17410_ (.A(_10426_),
    .B(_10428_),
    .Y(_10429_));
 sky130_fd_sc_hd__and2_1 _17411_ (.A(_10426_),
    .B(_10428_),
    .X(_10430_));
 sky130_fd_sc_hd__nor2_1 _17412_ (.A(_10429_),
    .B(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__xnor2_1 _17413_ (.A(_10378_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__a21oi_1 _17414_ (.A1(_10259_),
    .A2(_10314_),
    .B1(_10312_),
    .Y(_10433_));
 sky130_fd_sc_hd__xor2_1 _17415_ (.A(_10432_),
    .B(_10433_),
    .X(_10434_));
 sky130_fd_sc_hd__nand2_1 _17416_ (.A(_10348_),
    .B(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__or2_1 _17417_ (.A(_10348_),
    .B(_10434_),
    .X(_10436_));
 sky130_fd_sc_hd__nand2_1 _17418_ (.A(_10435_),
    .B(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__a21oi_1 _17419_ (.A1(_10226_),
    .A2(_10319_),
    .B1(_10317_),
    .Y(_10438_));
 sky130_fd_sc_hd__xor2_1 _17420_ (.A(_10437_),
    .B(_10438_),
    .X(_10439_));
 sky130_fd_sc_hd__nand2_1 _17421_ (.A(_10224_),
    .B(_10439_),
    .Y(_10440_));
 sky130_fd_sc_hd__or2_1 _17422_ (.A(_10224_),
    .B(_10439_),
    .X(_10441_));
 sky130_fd_sc_hd__nand2_1 _17423_ (.A(_10440_),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__a21o_1 _17424_ (.A1(_10342_),
    .A2(_10323_),
    .B1(_10442_),
    .X(_10443_));
 sky130_fd_sc_hd__and3_1 _17425_ (.A(_10342_),
    .B(_10323_),
    .C(_10442_),
    .X(_10444_));
 sky130_fd_sc_hd__inv_2 _17426_ (.A(_10444_),
    .Y(_10445_));
 sky130_fd_sc_hd__nand2_1 _17427_ (.A(_10443_),
    .B(_10445_),
    .Y(_10446_));
 sky130_fd_sc_hd__inv_2 _17428_ (.A(_10329_),
    .Y(_10447_));
 sky130_fd_sc_hd__o21a_1 _17429_ (.A1(_10447_),
    .A2(_10332_),
    .B1(_10327_),
    .X(_01663_));
 sky130_fd_sc_hd__a21oi_1 _17430_ (.A1(_10446_),
    .A2(_01663_),
    .B1(_08195_),
    .Y(_01664_));
 sky130_fd_sc_hd__o21ai_4 _17431_ (.A1(_10446_),
    .A2(_01663_),
    .B1(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__and2_1 _17432_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_01666_));
 sky130_fd_sc_hd__nor2_1 _17433_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_01667_));
 sky130_fd_sc_hd__o211a_1 _17434_ (.A1(_01666_),
    .A2(_01667_),
    .B1(_10336_),
    .C1(_10340_),
    .X(_01668_));
 sky130_fd_sc_hd__a211oi_2 _17435_ (.A1(_10336_),
    .A2(_10340_),
    .B1(_01666_),
    .C1(_01667_),
    .Y(_01669_));
 sky130_fd_sc_hd__o31a_1 _17436_ (.A1(_08156_),
    .A2(_01668_),
    .A3(_01669_),
    .B1(_09883_),
    .X(_01670_));
 sky130_fd_sc_hd__o2bb2a_1 _17437_ (.A1_N(_01665_),
    .A2_N(_01670_),
    .B1(\rbzero.wall_tracer.trackDistX[3] ),
    .B2(_09884_),
    .X(_00542_));
 sky130_fd_sc_hd__nand2_1 _17438_ (.A(_10351_),
    .B(_10376_),
    .Y(_01671_));
 sky130_fd_sc_hd__or2b_1 _17439_ (.A(_10377_),
    .B_N(_10349_),
    .X(_01672_));
 sky130_fd_sc_hd__o2bb2a_1 _17440_ (.A1_N(_10359_),
    .A2_N(_10360_),
    .B1(_10357_),
    .B2(_10358_),
    .X(_01673_));
 sky130_fd_sc_hd__a21oi_2 _17441_ (.A1(_01671_),
    .A2(_01672_),
    .B1(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__and3_1 _17442_ (.A(_01671_),
    .B(_01672_),
    .C(_01673_),
    .X(_01675_));
 sky130_fd_sc_hd__nor2_1 _17443_ (.A(_01674_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21o_1 _17444_ (.A1(_10361_),
    .A2(_10375_),
    .B1(_10373_),
    .X(_01677_));
 sky130_fd_sc_hd__or2b_1 _17445_ (.A(_10397_),
    .B_N(_10381_),
    .X(_01678_));
 sky130_fd_sc_hd__or2b_1 _17446_ (.A(_10398_),
    .B_N(_10379_),
    .X(_01679_));
 sky130_fd_sc_hd__o22ai_1 _17447_ (.A1(_10012_),
    .A2(_09314_),
    .B1(_09441_),
    .B2(_09466_),
    .Y(_01680_));
 sky130_fd_sc_hd__or4_1 _17448_ (.A(_10012_),
    .B(_09466_),
    .C(_09313_),
    .D(_09440_),
    .X(_01681_));
 sky130_fd_sc_hd__nand2_1 _17449_ (.A(_01680_),
    .B(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__nor2_1 _17450_ (.A(_09347_),
    .B(_09571_),
    .Y(_01683_));
 sky130_fd_sc_hd__xor2_1 _17451_ (.A(_01682_),
    .B(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__o31a_1 _17452_ (.A1(_09466_),
    .A2(_09314_),
    .A3(_10230_),
    .B1(_10355_),
    .X(_01685_));
 sky130_fd_sc_hd__xor2_1 _17453_ (.A(_01684_),
    .B(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__and2_1 _17454_ (.A(_09228_),
    .B(_09691_),
    .X(_01687_));
 sky130_fd_sc_hd__xor2_1 _17455_ (.A(_01686_),
    .B(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__a21bo_1 _17456_ (.A1(_10363_),
    .A2(_10366_),
    .B1_N(_10364_),
    .X(_01689_));
 sky130_fd_sc_hd__nand2_1 _17457_ (.A(_10266_),
    .B(_10383_),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _17458_ (.A(_01690_),
    .B(_10385_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_2 _17459_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08321_),
    .Y(_01692_));
 sky130_fd_sc_hd__or2b_1 _17460_ (.A(_09156_),
    .B_N(_08238_),
    .X(_01693_));
 sky130_fd_sc_hd__or3_1 _17461_ (.A(_10140_),
    .B(_01692_),
    .C(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__o21ai_1 _17462_ (.A1(_10140_),
    .A2(_01692_),
    .B1(_01693_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _17463_ (.A(_01694_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__nor2_1 _17464_ (.A(_10144_),
    .B(_09213_),
    .Y(_01697_));
 sky130_fd_sc_hd__xor2_1 _17465_ (.A(_01696_),
    .B(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__xnor2_1 _17466_ (.A(_01691_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__xnor2_1 _17467_ (.A(_01689_),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__a21oi_1 _17468_ (.A1(_10362_),
    .A2(_10370_),
    .B1(_10368_),
    .Y(_01701_));
 sky130_fd_sc_hd__nor2_1 _17469_ (.A(_01700_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__and2_1 _17470_ (.A(_01700_),
    .B(_01701_),
    .X(_01703_));
 sky130_fd_sc_hd__nor2_1 _17471_ (.A(_01702_),
    .B(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__xnor2_1 _17472_ (.A(_01688_),
    .B(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__a21o_1 _17473_ (.A1(_01678_),
    .A2(_01679_),
    .B1(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__nand3_1 _17474_ (.A(_01678_),
    .B(_01679_),
    .C(_01705_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _17475_ (.A(_01706_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__xnor2_1 _17476_ (.A(_01677_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__nor2_1 _17477_ (.A(_10393_),
    .B(_10395_),
    .Y(_01710_));
 sky130_fd_sc_hd__a21o_1 _17478_ (.A1(_10388_),
    .A2(_10396_),
    .B1(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__or2b_1 _17479_ (.A(_10410_),
    .B_N(_10401_),
    .X(_01712_));
 sky130_fd_sc_hd__a21bo_1 _17480_ (.A1(_10405_),
    .A2(_10409_),
    .B1_N(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__inv_2 _17481_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .Y(_01714_));
 sky130_fd_sc_hd__nand2_1 _17482_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08321_),
    .Y(_01715_));
 sky130_fd_sc_hd__buf_2 _17483_ (.A(_08330_),
    .X(_01716_));
 sky130_fd_sc_hd__or4_1 _17484_ (.A(_10265_),
    .B(_01715_),
    .C(_08336_),
    .D(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__buf_2 _17485_ (.A(_01715_),
    .X(_01718_));
 sky130_fd_sc_hd__o22ai_1 _17486_ (.A1(_01718_),
    .A2(_08336_),
    .B1(_01716_),
    .B2(_10265_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _17487_ (.A(_01717_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__or3_1 _17488_ (.A(_01714_),
    .B(_08335_),
    .C(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__o21ai_1 _17489_ (.A1(_01714_),
    .A2(_08335_),
    .B1(_01720_),
    .Y(_01722_));
 sky130_fd_sc_hd__and2_1 _17490_ (.A(_01721_),
    .B(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__nor2_1 _17491_ (.A(_08583_),
    .B(_09633_),
    .Y(_01724_));
 sky130_fd_sc_hd__nor2_1 _17492_ (.A(_08808_),
    .B(_09630_),
    .Y(_01725_));
 sky130_fd_sc_hd__xnor2_1 _17493_ (.A(_01724_),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__or2_1 _17494_ (.A(_09358_),
    .B(_09497_),
    .X(_01727_));
 sky130_fd_sc_hd__xnor2_1 _17495_ (.A(_01726_),
    .B(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__buf_2 _17496_ (.A(_09358_),
    .X(_01729_));
 sky130_fd_sc_hd__o31a_1 _17497_ (.A1(_01729_),
    .A2(_09495_),
    .A3(_10391_),
    .B1(_10389_),
    .X(_01730_));
 sky130_fd_sc_hd__xor2_1 _17498_ (.A(_01728_),
    .B(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__xnor2_1 _17499_ (.A(_01723_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__xor2_1 _17500_ (.A(_01713_),
    .B(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__xnor2_1 _17501_ (.A(_01711_),
    .B(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__or3_1 _17502_ (.A(_10159_),
    .B(_09630_),
    .C(_10407_),
    .X(_01735_));
 sky130_fd_sc_hd__a21bo_1 _17503_ (.A1(_10400_),
    .A2(_10406_),
    .B1_N(_01735_),
    .X(_01736_));
 sky130_fd_sc_hd__buf_2 _17504_ (.A(_10403_),
    .X(_01737_));
 sky130_fd_sc_hd__o31ai_1 _17505_ (.A1(_09751_),
    .A2(_01737_),
    .A3(_10416_),
    .B1(_10404_),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _17506_ (.A(_08469_),
    .B(_09763_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _17507_ (.A(_09372_),
    .B(_10403_),
    .Y(_01740_));
 sky130_fd_sc_hd__xor2_1 _17508_ (.A(_01739_),
    .B(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__nor2_1 _17509_ (.A(_10159_),
    .B(_10173_),
    .Y(_01742_));
 sky130_fd_sc_hd__xor2_1 _17510_ (.A(_01741_),
    .B(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__xnor2_1 _17511_ (.A(_01738_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__xor2_1 _17512_ (.A(_01736_),
    .B(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__nand2_1 _17513_ (.A(_10182_),
    .B(_10418_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _17514_ (.A(_09751_),
    .B(_10414_),
    .Y(_01747_));
 sky130_fd_sc_hd__mux2_1 _17515_ (.A0(_09751_),
    .A1(_01747_),
    .S(_10416_),
    .X(_01748_));
 sky130_fd_sc_hd__xnor2_1 _17516_ (.A(_10182_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__a21oi_1 _17517_ (.A1(_10180_),
    .A2(_01746_),
    .B1(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__and3_1 _17518_ (.A(_10180_),
    .B(_01746_),
    .C(_01749_),
    .X(_01751_));
 sky130_fd_sc_hd__nor2_1 _17519_ (.A(_01750_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__xnor2_1 _17520_ (.A(_01745_),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__and2b_1 _17521_ (.A_N(_10419_),
    .B(_10420_),
    .X(_01754_));
 sky130_fd_sc_hd__a21oi_1 _17522_ (.A1(_10411_),
    .A2(_10421_),
    .B1(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__xor2_1 _17523_ (.A(_01753_),
    .B(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__xnor2_1 _17524_ (.A(_01734_),
    .B(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__and2b_1 _17525_ (.A_N(_10422_),
    .B(_10424_),
    .X(_01758_));
 sky130_fd_sc_hd__a21oi_1 _17526_ (.A1(_10399_),
    .A2(_10425_),
    .B1(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__xor2_1 _17527_ (.A(_01757_),
    .B(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__xnor2_1 _17528_ (.A(_01709_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__a21oi_1 _17529_ (.A1(_10378_),
    .A2(_10431_),
    .B1(_10429_),
    .Y(_01762_));
 sky130_fd_sc_hd__nor2_1 _17530_ (.A(_01761_),
    .B(_01762_),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _17531_ (.A(_01761_),
    .B(_01762_),
    .Y(_01764_));
 sky130_fd_sc_hd__and2b_1 _17532_ (.A_N(_01763_),
    .B(_01764_),
    .X(_01765_));
 sky130_fd_sc_hd__xnor2_1 _17533_ (.A(_01676_),
    .B(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__o21a_1 _17534_ (.A1(_10432_),
    .A2(_10433_),
    .B1(_10435_),
    .X(_01767_));
 sky130_fd_sc_hd__xor2_1 _17535_ (.A(_01766_),
    .B(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__nand2_1 _17536_ (.A(_10346_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__or2_1 _17537_ (.A(_10346_),
    .B(_01768_),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_1 _17538_ (.A(_01769_),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__o21a_1 _17539_ (.A1(_10437_),
    .A2(_10438_),
    .B1(_10440_),
    .X(_01772_));
 sky130_fd_sc_hd__xor2_2 _17540_ (.A(_01771_),
    .B(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__nand3_1 _17541_ (.A(_10329_),
    .B(_10443_),
    .C(_10445_),
    .Y(_01774_));
 sky130_fd_sc_hd__a21oi_1 _17542_ (.A1(_10327_),
    .A2(_10443_),
    .B1(_10444_),
    .Y(_01775_));
 sky130_fd_sc_hd__o21bai_2 _17543_ (.A1(_10332_),
    .A2(_01774_),
    .B1_N(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__a21oi_1 _17544_ (.A1(_01773_),
    .A2(_01776_),
    .B1(_08195_),
    .Y(_01777_));
 sky130_fd_sc_hd__o21ai_4 _17545_ (.A1(_01773_),
    .A2(_01776_),
    .B1(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__buf_4 _17546_ (.A(_08155_),
    .X(_01779_));
 sky130_fd_sc_hd__nand2_1 _17547_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_01780_));
 sky130_fd_sc_hd__or2_1 _17548_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_01781_));
 sky130_fd_sc_hd__o211a_1 _17549_ (.A1(_01666_),
    .A2(_01669_),
    .B1(_01780_),
    .C1(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__a211oi_1 _17550_ (.A1(_01780_),
    .A2(_01781_),
    .B1(_01666_),
    .C1(_01669_),
    .Y(_01783_));
 sky130_fd_sc_hd__o31a_1 _17551_ (.A1(_01779_),
    .A2(_01782_),
    .A3(_01783_),
    .B1(_09883_),
    .X(_01784_));
 sky130_fd_sc_hd__o2bb2a_1 _17552_ (.A1_N(_01778_),
    .A2_N(_01784_),
    .B1(\rbzero.wall_tracer.trackDistX[4] ),
    .B2(_09884_),
    .X(_00543_));
 sky130_fd_sc_hd__nor2_1 _17553_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_01785_));
 sky130_fd_sc_hd__and2_1 _17554_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_01786_));
 sky130_fd_sc_hd__a21oi_1 _17555_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(\rbzero.wall_tracer.stepDistX[4] ),
    .B1(_01782_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor3_1 _17556_ (.A(_01785_),
    .B(_01786_),
    .C(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__o21a_1 _17557_ (.A1(_01785_),
    .A2(_01786_),
    .B1(_01787_),
    .X(_01789_));
 sky130_fd_sc_hd__or2_1 _17558_ (.A(_01766_),
    .B(_01767_),
    .X(_01790_));
 sky130_fd_sc_hd__or2b_1 _17559_ (.A(_01708_),
    .B_N(_01677_),
    .X(_01791_));
 sky130_fd_sc_hd__o2bb2a_1 _17560_ (.A1_N(_01686_),
    .A2_N(_01687_),
    .B1(_01684_),
    .B2(_01685_),
    .X(_01792_));
 sky130_fd_sc_hd__a21oi_4 _17561_ (.A1(_01706_),
    .A2(_01791_),
    .B1(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__and3_1 _17562_ (.A(_01706_),
    .B(_01791_),
    .C(_01792_),
    .X(_01794_));
 sky130_fd_sc_hd__nor2_1 _17563_ (.A(_01793_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21o_1 _17564_ (.A1(_01688_),
    .A2(_01704_),
    .B1(_01702_),
    .X(_01796_));
 sky130_fd_sc_hd__or2b_1 _17565_ (.A(_01732_),
    .B_N(_01713_),
    .X(_01797_));
 sky130_fd_sc_hd__or2b_1 _17566_ (.A(_01733_),
    .B_N(_01711_),
    .X(_01798_));
 sky130_fd_sc_hd__o22ai_1 _17567_ (.A1(_10144_),
    .A2(_09314_),
    .B1(_09441_),
    .B2(_10012_),
    .Y(_01799_));
 sky130_fd_sc_hd__or4_1 _17568_ (.A(_10012_),
    .B(_10144_),
    .C(_09313_),
    .D(_09441_),
    .X(_01800_));
 sky130_fd_sc_hd__nand2_1 _17569_ (.A(_01799_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__nor2_1 _17570_ (.A(_09466_),
    .B(_09571_),
    .Y(_01802_));
 sky130_fd_sc_hd__xor2_1 _17571_ (.A(_01801_),
    .B(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__o31a_1 _17572_ (.A1(_09347_),
    .A2(_09571_),
    .A3(_01682_),
    .B1(_01681_),
    .X(_01804_));
 sky130_fd_sc_hd__xor2_1 _17573_ (.A(_01803_),
    .B(_01804_),
    .X(_01805_));
 sky130_fd_sc_hd__and2_1 _17574_ (.A(_09347_),
    .B(_09691_),
    .X(_01806_));
 sky130_fd_sc_hd__xor2_1 _17575_ (.A(_01805_),
    .B(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__o31ai_2 _17576_ (.A1(_10144_),
    .A2(_09213_),
    .A3(_01696_),
    .B1(_01694_),
    .Y(_01808_));
 sky130_fd_sc_hd__inv_2 _17577_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_1 _17578_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08321_),
    .Y(_01810_));
 sky130_fd_sc_hd__or4_1 _17579_ (.A(_01809_),
    .B(_10140_),
    .C(_08335_),
    .D(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__a32o_1 _17580_ (.A1(\rbzero.wall_tracer.visualWallDist[5] ),
    .A2(_08496_),
    .A3(_08228_),
    .B1(_08339_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_01812_));
 sky130_fd_sc_hd__nand2_1 _17581_ (.A(_01811_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__nor2_1 _17582_ (.A(_10262_),
    .B(_09213_),
    .Y(_01814_));
 sky130_fd_sc_hd__xor2_1 _17583_ (.A(_01813_),
    .B(_01814_),
    .X(_01815_));
 sky130_fd_sc_hd__a21oi_1 _17584_ (.A1(_01717_),
    .A2(_01721_),
    .B1(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__and3_1 _17585_ (.A(_01717_),
    .B(_01721_),
    .C(_01815_),
    .X(_01817_));
 sky130_fd_sc_hd__nor2_1 _17586_ (.A(_01816_),
    .B(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__xnor2_1 _17587_ (.A(_01808_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__a21oi_1 _17588_ (.A1(_01690_),
    .A2(_10385_),
    .B1(_01698_),
    .Y(_01820_));
 sky130_fd_sc_hd__a21oi_1 _17589_ (.A1(_01689_),
    .A2(_01699_),
    .B1(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__nor2_1 _17590_ (.A(_01819_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__and2_1 _17591_ (.A(_01819_),
    .B(_01821_),
    .X(_01823_));
 sky130_fd_sc_hd__nor2_1 _17592_ (.A(_01822_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__xnor2_1 _17593_ (.A(_01807_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__a21o_1 _17594_ (.A1(_01797_),
    .A2(_01798_),
    .B1(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__nand3_1 _17595_ (.A(_01797_),
    .B(_01798_),
    .C(_01825_),
    .Y(_01827_));
 sky130_fd_sc_hd__nand2_1 _17596_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__xnor2_1 _17597_ (.A(_01796_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__nor2_1 _17598_ (.A(_01728_),
    .B(_01730_),
    .Y(_01830_));
 sky130_fd_sc_hd__a21o_1 _17599_ (.A1(_01723_),
    .A2(_01731_),
    .B1(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__or2b_1 _17600_ (.A(_01743_),
    .B_N(_01738_),
    .X(_01832_));
 sky130_fd_sc_hd__nand2_1 _17601_ (.A(_01736_),
    .B(_01744_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_2 _17602_ (.A(_06340_),
    .B(_09019_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _17603_ (.A(_10265_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor2_1 _17604_ (.A(_01718_),
    .B(_01716_),
    .Y(_01836_));
 sky130_fd_sc_hd__xnor2_1 _17605_ (.A(_01835_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__or3_1 _17606_ (.A(_01714_),
    .B(_08336_),
    .C(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__o21ai_1 _17607_ (.A1(_01714_),
    .A2(_08336_),
    .B1(_01837_),
    .Y(_01839_));
 sky130_fd_sc_hd__and2_1 _17608_ (.A(_01838_),
    .B(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__nor2_1 _17609_ (.A(_08583_),
    .B(_10173_),
    .Y(_01841_));
 sky130_fd_sc_hd__o22a_1 _17610_ (.A1(_08583_),
    .A2(_09630_),
    .B1(_10173_),
    .B2(_08809_),
    .X(_01842_));
 sky130_fd_sc_hd__a21o_1 _17611_ (.A1(_01725_),
    .A2(_01841_),
    .B1(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__nor2_1 _17612_ (.A(_09358_),
    .B(_09633_),
    .Y(_01844_));
 sky130_fd_sc_hd__xor2_1 _17613_ (.A(_01843_),
    .B(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__o2bb2a_1 _17614_ (.A1_N(_01724_),
    .A2_N(_01725_),
    .B1(_01726_),
    .B2(_01727_),
    .X(_01846_));
 sky130_fd_sc_hd__nor2_1 _17615_ (.A(_01845_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__and2_1 _17616_ (.A(_01845_),
    .B(_01846_),
    .X(_01848_));
 sky130_fd_sc_hd__nor2_1 _17617_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__xnor2_1 _17618_ (.A(_01840_),
    .B(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__a21o_1 _17619_ (.A1(_01832_),
    .A2(_01833_),
    .B1(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__nand3_1 _17620_ (.A(_01832_),
    .B(_01833_),
    .C(_01850_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _17621_ (.A(_01851_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__xnor2_1 _17622_ (.A(_01831_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__and2b_1 _17623_ (.A_N(_01741_),
    .B(_01742_),
    .X(_01855_));
 sky130_fd_sc_hd__a31o_1 _17624_ (.A1(_08469_),
    .A2(_09763_),
    .A3(_01740_),
    .B1(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__o21ai_4 _17625_ (.A1(_09751_),
    .A2(_10416_),
    .B1(_10404_),
    .Y(_01857_));
 sky130_fd_sc_hd__or3_1 _17626_ (.A(_09372_),
    .B(_09371_),
    .C(_10414_),
    .X(_01858_));
 sky130_fd_sc_hd__o22a_1 _17627_ (.A1(_09372_),
    .A2(_10414_),
    .B1(_10403_),
    .B2(_09371_),
    .X(_01859_));
 sky130_fd_sc_hd__o21ba_1 _17628_ (.A1(_10403_),
    .A2(_01858_),
    .B1_N(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__and2b_1 _17629_ (.A_N(_10159_),
    .B(_09763_),
    .X(_01861_));
 sky130_fd_sc_hd__xor2_1 _17630_ (.A(_01860_),
    .B(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__xnor2_1 _17631_ (.A(_01857_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__xnor2_1 _17632_ (.A(_01856_),
    .B(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__or2b_1 _17633_ (.A(_10180_),
    .B_N(_01748_),
    .X(_01865_));
 sky130_fd_sc_hd__or2_1 _17634_ (.A(_10179_),
    .B(_01748_),
    .X(_01866_));
 sky130_fd_sc_hd__and2_1 _17635_ (.A(_01865_),
    .B(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__buf_2 _17636_ (.A(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__xnor2_1 _17637_ (.A(_01864_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__a21oi_1 _17638_ (.A1(_01745_),
    .A2(_01752_),
    .B1(_01750_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _17639_ (.A(_01869_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__nand2_1 _17640_ (.A(_01869_),
    .B(_01870_),
    .Y(_01872_));
 sky130_fd_sc_hd__and2b_1 _17641_ (.A_N(_01871_),
    .B(_01872_),
    .X(_01873_));
 sky130_fd_sc_hd__xnor2_1 _17642_ (.A(_01854_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _17643_ (.A(_01753_),
    .B(_01755_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21oi_1 _17644_ (.A1(_01734_),
    .A2(_01756_),
    .B1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__xor2_1 _17645_ (.A(_01874_),
    .B(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__xnor2_1 _17646_ (.A(_01829_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _17647_ (.A(_01757_),
    .B(_01759_),
    .Y(_01879_));
 sky130_fd_sc_hd__a21oi_1 _17648_ (.A1(_01709_),
    .A2(_01760_),
    .B1(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__xor2_1 _17649_ (.A(_01878_),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__xnor2_1 _17650_ (.A(_01795_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21oi_1 _17651_ (.A1(_01676_),
    .A2(_01764_),
    .B1(_01763_),
    .Y(_01883_));
 sky130_fd_sc_hd__nor2_1 _17652_ (.A(_01882_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_1 _17653_ (.A(_01882_),
    .B(_01883_),
    .Y(_01885_));
 sky130_fd_sc_hd__and2b_1 _17654_ (.A_N(_01884_),
    .B(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__xnor2_1 _17655_ (.A(_01674_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__and3_1 _17656_ (.A(_01790_),
    .B(_01769_),
    .C(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__a21oi_1 _17657_ (.A1(_01790_),
    .A2(_01769_),
    .B1(_01887_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor2_2 _17658_ (.A(_01888_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__or2_1 _17659_ (.A(_01771_),
    .B(_01772_),
    .X(_01891_));
 sky130_fd_sc_hd__a21boi_2 _17660_ (.A1(_01773_),
    .A2(_01776_),
    .B1_N(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__xnor2_4 _17661_ (.A(_01890_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _17662_ (.A(_09905_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__o311a_1 _17663_ (.A1(_06164_),
    .A2(_01788_),
    .A3(_01789_),
    .B1(_09917_),
    .C1(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__a21oi_1 _17664_ (.A1(_06206_),
    .A2(_09860_),
    .B1(_01895_),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_1 _17665_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01896_));
 sky130_fd_sc_hd__and2_1 _17666_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .X(_01897_));
 sky130_fd_sc_hd__o21ba_1 _17667_ (.A1(_01785_),
    .A2(_01787_),
    .B1_N(_01786_),
    .X(_01898_));
 sky130_fd_sc_hd__o21ai_1 _17668_ (.A1(_01896_),
    .A2(_01897_),
    .B1(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__o31a_1 _17669_ (.A1(_01896_),
    .A2(_01897_),
    .A3(_01898_),
    .B1(_08193_),
    .X(_01900_));
 sky130_fd_sc_hd__or2b_1 _17670_ (.A(_01828_),
    .B_N(_01796_),
    .X(_01901_));
 sky130_fd_sc_hd__o2bb2a_2 _17671_ (.A1_N(_01805_),
    .A2_N(_01806_),
    .B1(_01803_),
    .B2(_01804_),
    .X(_01902_));
 sky130_fd_sc_hd__a21oi_4 _17672_ (.A1(_01826_),
    .A2(_01901_),
    .B1(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__and3_1 _17673_ (.A(_01826_),
    .B(_01901_),
    .C(_01902_),
    .X(_01904_));
 sky130_fd_sc_hd__nor2_1 _17674_ (.A(_01903_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__a21o_1 _17675_ (.A1(_01807_),
    .A2(_01824_),
    .B1(_01822_),
    .X(_01906_));
 sky130_fd_sc_hd__or2b_1 _17676_ (.A(_01853_),
    .B_N(_01831_),
    .X(_01907_));
 sky130_fd_sc_hd__o22a_1 _17677_ (.A1(_10262_),
    .A2(_09314_),
    .B1(_09441_),
    .B2(_10144_),
    .X(_01908_));
 sky130_fd_sc_hd__or4_1 _17678_ (.A(_10262_),
    .B(_10144_),
    .C(_09314_),
    .D(_09441_),
    .X(_01909_));
 sky130_fd_sc_hd__or2b_1 _17679_ (.A(_01908_),
    .B_N(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__nor2_1 _17680_ (.A(_10012_),
    .B(_09706_),
    .Y(_01911_));
 sky130_fd_sc_hd__xor2_1 _17681_ (.A(_01910_),
    .B(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__o31a_1 _17682_ (.A1(_09466_),
    .A2(_09706_),
    .A3(_01801_),
    .B1(_01800_),
    .X(_01913_));
 sky130_fd_sc_hd__xnor2_1 _17683_ (.A(_01912_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _17684_ (.A(_08779_),
    .B(_09687_),
    .Y(_01915_));
 sky130_fd_sc_hd__xnor2_1 _17685_ (.A(_01914_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__a21bo_1 _17686_ (.A1(_01812_),
    .A2(_01814_),
    .B1_N(_01811_),
    .X(_01917_));
 sky130_fd_sc_hd__nand2_1 _17687_ (.A(_01835_),
    .B(_01836_),
    .Y(_01918_));
 sky130_fd_sc_hd__nand2_1 _17688_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08321_),
    .Y(_01919_));
 sky130_fd_sc_hd__or2_1 _17689_ (.A(_10140_),
    .B(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__or2_1 _17690_ (.A(_08303_),
    .B(_09159_),
    .X(_01921_));
 sky130_fd_sc_hd__or3_1 _17691_ (.A(_01809_),
    .B(_08304_),
    .C(_08336_),
    .X(_01922_));
 sky130_fd_sc_hd__xnor2_1 _17692_ (.A(_01921_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__or2_1 _17693_ (.A(_01920_),
    .B(_01923_),
    .X(_01924_));
 sky130_fd_sc_hd__nand2_1 _17694_ (.A(_01920_),
    .B(_01923_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(_01924_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__a21oi_1 _17696_ (.A1(_01918_),
    .A2(_01838_),
    .B1(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__and3_1 _17697_ (.A(_01918_),
    .B(_01838_),
    .C(_01926_),
    .X(_01928_));
 sky130_fd_sc_hd__nor2_1 _17698_ (.A(_01927_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__xnor2_1 _17699_ (.A(_01917_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__a21oi_1 _17700_ (.A1(_01808_),
    .A2(_01818_),
    .B1(_01816_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _17701_ (.A(_01930_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__and2_1 _17702_ (.A(_01930_),
    .B(_01931_),
    .X(_01933_));
 sky130_fd_sc_hd__nor2_1 _17703_ (.A(_01932_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_01916_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__a21o_1 _17705_ (.A1(_01851_),
    .A2(_01907_),
    .B1(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__nand3_1 _17706_ (.A(_01851_),
    .B(_01907_),
    .C(_01935_),
    .Y(_01937_));
 sky130_fd_sc_hd__nand2_1 _17707_ (.A(_01936_),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__xnor2_1 _17708_ (.A(_01906_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__a21o_1 _17709_ (.A1(_01840_),
    .A2(_01849_),
    .B1(_01847_),
    .X(_01940_));
 sky130_fd_sc_hd__nand2_1 _17710_ (.A(_01857_),
    .B(_01862_),
    .Y(_01941_));
 sky130_fd_sc_hd__or2b_1 _17711_ (.A(_01863_),
    .B_N(_01856_),
    .X(_01942_));
 sky130_fd_sc_hd__or4_1 _17712_ (.A(_10265_),
    .B(_01718_),
    .C(_01834_),
    .D(_10163_),
    .X(_01943_));
 sky130_fd_sc_hd__o22ai_1 _17713_ (.A1(_01718_),
    .A2(_01834_),
    .B1(_10163_),
    .B2(_10265_),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_1 _17714_ (.A(_01943_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__or3_1 _17715_ (.A(_01716_),
    .B(_10386_),
    .C(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__o21ai_1 _17716_ (.A1(_01716_),
    .A2(_10386_),
    .B1(_01945_),
    .Y(_01947_));
 sky130_fd_sc_hd__and2_1 _17717_ (.A(_01946_),
    .B(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__or2_1 _17718_ (.A(_08583_),
    .B(_10173_),
    .X(_01949_));
 sky130_fd_sc_hd__or2b_1 _17719_ (.A(_08809_),
    .B_N(_09763_),
    .X(_01950_));
 sky130_fd_sc_hd__xnor2_1 _17720_ (.A(_01949_),
    .B(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__or3_1 _17721_ (.A(_01729_),
    .B(_09630_),
    .C(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__o21ai_1 _17722_ (.A1(_01729_),
    .A2(_09630_),
    .B1(_01951_),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_1 _17723_ (.A(_01952_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_1 _17724_ (.A(_01725_),
    .B(_01841_),
    .Y(_01955_));
 sky130_fd_sc_hd__o31a_1 _17725_ (.A1(_01729_),
    .A2(_09633_),
    .A3(_01842_),
    .B1(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__nor2_1 _17726_ (.A(_01954_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__and2_1 _17727_ (.A(_01954_),
    .B(_01956_),
    .X(_01958_));
 sky130_fd_sc_hd__nor2_1 _17728_ (.A(_01957_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__xnor2_1 _17729_ (.A(_01948_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__a21o_1 _17730_ (.A1(_01941_),
    .A2(_01942_),
    .B1(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__nand3_1 _17731_ (.A(_01941_),
    .B(_01942_),
    .C(_01960_),
    .Y(_01962_));
 sky130_fd_sc_hd__nand2_1 _17732_ (.A(_01961_),
    .B(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__xnor2_1 _17733_ (.A(_01940_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__a2bb2o_1 _17734_ (.A1_N(_01737_),
    .A2_N(_01858_),
    .B1(_01860_),
    .B2(_01861_),
    .X(_01965_));
 sky130_fd_sc_hd__a21oi_1 _17735_ (.A1(_09372_),
    .A2(_09371_),
    .B1(_10414_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(_01858_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _17737_ (.A(_10159_),
    .B(_01737_),
    .Y(_01968_));
 sky130_fd_sc_hd__xnor2_1 _17738_ (.A(_01967_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__xor2_1 _17739_ (.A(_01857_),
    .B(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_1 _17740_ (.A(_01965_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__or2_1 _17741_ (.A(_01965_),
    .B(_01970_),
    .X(_01972_));
 sky130_fd_sc_hd__and2_1 _17742_ (.A(_01971_),
    .B(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__xnor2_1 _17743_ (.A(_01868_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__inv_2 _17744_ (.A(_01865_),
    .Y(_01975_));
 sky130_fd_sc_hd__a21oi_1 _17745_ (.A1(_01864_),
    .A2(_01868_),
    .B1(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__nor2_1 _17746_ (.A(_01974_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__and2_1 _17747_ (.A(_01974_),
    .B(_01976_),
    .X(_01978_));
 sky130_fd_sc_hd__nor2_1 _17748_ (.A(_01977_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__xnor2_1 _17749_ (.A(_01964_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21oi_1 _17750_ (.A1(_01854_),
    .A2(_01872_),
    .B1(_01871_),
    .Y(_01981_));
 sky130_fd_sc_hd__xor2_1 _17751_ (.A(_01980_),
    .B(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__xnor2_1 _17752_ (.A(_01939_),
    .B(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _17753_ (.A(_01874_),
    .B(_01876_),
    .Y(_01984_));
 sky130_fd_sc_hd__a21oi_2 _17754_ (.A1(_01829_),
    .A2(_01877_),
    .B1(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__xor2_1 _17755_ (.A(_01983_),
    .B(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__xnor2_1 _17756_ (.A(_01905_),
    .B(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2_1 _17757_ (.A(_01878_),
    .B(_01880_),
    .Y(_01988_));
 sky130_fd_sc_hd__a21oi_2 _17758_ (.A1(_01795_),
    .A2(_01881_),
    .B1(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__or2_1 _17759_ (.A(_01987_),
    .B(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__nand2_1 _17760_ (.A(_01987_),
    .B(_01989_),
    .Y(_01991_));
 sky130_fd_sc_hd__and2_1 _17761_ (.A(_01990_),
    .B(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__nand2_1 _17762_ (.A(_01793_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__or2_1 _17763_ (.A(_01793_),
    .B(_01992_),
    .X(_01994_));
 sky130_fd_sc_hd__nand2_1 _17764_ (.A(_01993_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__a21oi_4 _17765_ (.A1(_01674_),
    .A2(_01885_),
    .B1(_01884_),
    .Y(_01996_));
 sky130_fd_sc_hd__or2_1 _17766_ (.A(_01995_),
    .B(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _17767_ (.A(_01995_),
    .B(_01996_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_1 _17768_ (.A(_01997_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__or3b_1 _17769_ (.A(_01888_),
    .B(_01889_),
    .C_N(_01773_),
    .X(_02000_));
 sky130_fd_sc_hd__or2b_1 _17770_ (.A(_02000_),
    .B_N(_01775_),
    .X(_02001_));
 sky130_fd_sc_hd__o31a_2 _17771_ (.A1(_10332_),
    .A2(_01774_),
    .A3(_02000_),
    .B1(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__o21ba_2 _17772_ (.A1(_01891_),
    .A2(_01888_),
    .B1_N(_01889_),
    .X(_02003_));
 sky130_fd_sc_hd__and3_1 _17773_ (.A(_01999_),
    .B(_02002_),
    .C(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__a21o_1 _17774_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_01999_),
    .X(_02005_));
 sky130_fd_sc_hd__or3b_1 _17775_ (.A(_08192_),
    .B(_02004_),
    .C_N(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__a21bo_1 _17776_ (.A1(_01899_),
    .A2(_01900_),
    .B1_N(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _17777_ (.A0(\rbzero.wall_tracer.trackDistX[6] ),
    .A1(_02007_),
    .S(_09917_),
    .X(_02008_));
 sky130_fd_sc_hd__clkbuf_1 _17778_ (.A(_02008_),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _17779_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _17780_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_02010_));
 sky130_fd_sc_hd__or2b_1 _17781_ (.A(_02009_),
    .B_N(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__o21ba_1 _17782_ (.A1(_01896_),
    .A2(_01898_),
    .B1_N(_01897_),
    .X(_02012_));
 sky130_fd_sc_hd__nor2_1 _17783_ (.A(_02011_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__a21o_1 _17784_ (.A1(_02011_),
    .A2(_02012_),
    .B1(_08155_),
    .X(_02014_));
 sky130_fd_sc_hd__or2b_1 _17785_ (.A(_01938_),
    .B_N(_01906_),
    .X(_02015_));
 sky130_fd_sc_hd__o32a_1 _17786_ (.A1(_08779_),
    .A2(_09687_),
    .A3(_01914_),
    .B1(_01913_),
    .B2(_01912_),
    .X(_02016_));
 sky130_fd_sc_hd__a21oi_2 _17787_ (.A1(_01936_),
    .A2(_02015_),
    .B1(_02016_),
    .Y(_02017_));
 sky130_fd_sc_hd__and3_1 _17788_ (.A(_01936_),
    .B(_02015_),
    .C(_02016_),
    .X(_02018_));
 sky130_fd_sc_hd__nor2_1 _17789_ (.A(_02017_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__a21o_1 _17790_ (.A1(_01916_),
    .A2(_01934_),
    .B1(_01932_),
    .X(_02020_));
 sky130_fd_sc_hd__or2b_1 _17791_ (.A(_01963_),
    .B_N(_01940_),
    .X(_02021_));
 sky130_fd_sc_hd__and3_1 _17792_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08496_),
    .C(_08238_),
    .X(_02022_));
 sky130_fd_sc_hd__nand2_1 _17793_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08321_),
    .Y(_02023_));
 sky130_fd_sc_hd__nor2_1 _17794_ (.A(_10140_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _17795_ (.A(_02022_),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__or2_1 _17796_ (.A(_02022_),
    .B(_02024_),
    .X(_02026_));
 sky130_fd_sc_hd__nand2_1 _17797_ (.A(_02025_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _17798_ (.A(_10144_),
    .B(_09706_),
    .Y(_02028_));
 sky130_fd_sc_hd__xor2_1 _17799_ (.A(_02027_),
    .B(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__o31a_1 _17800_ (.A1(_10012_),
    .A2(_09706_),
    .A3(_01908_),
    .B1(_01909_),
    .X(_02030_));
 sky130_fd_sc_hd__xnor2_1 _17801_ (.A(_02029_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__nand2_1 _17802_ (.A(_10012_),
    .B(_09691_),
    .Y(_02032_));
 sky130_fd_sc_hd__xor2_1 _17803_ (.A(_02031_),
    .B(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__o21ai_1 _17804_ (.A1(_01921_),
    .A2(_01922_),
    .B1(_01924_),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _17805_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08340_),
    .Y(_02035_));
 sky130_fd_sc_hd__or3_1 _17806_ (.A(_01716_),
    .B(_01692_),
    .C(_02035_),
    .X(_02036_));
 sky130_fd_sc_hd__o21ai_1 _17807_ (.A1(_01716_),
    .A2(_01692_),
    .B1(_02035_),
    .Y(_02037_));
 sky130_fd_sc_hd__and2_1 _17808_ (.A(_02036_),
    .B(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__nor2_1 _17809_ (.A(_08303_),
    .B(_09213_),
    .Y(_02039_));
 sky130_fd_sc_hd__xnor2_1 _17810_ (.A(_02038_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__a21oi_1 _17811_ (.A1(_01943_),
    .A2(_01946_),
    .B1(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__and3_1 _17812_ (.A(_01943_),
    .B(_01946_),
    .C(_02040_),
    .X(_02042_));
 sky130_fd_sc_hd__nor2_1 _17813_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__xnor2_1 _17814_ (.A(_02034_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__a21oi_1 _17815_ (.A1(_01917_),
    .A2(_01929_),
    .B1(_01927_),
    .Y(_02045_));
 sky130_fd_sc_hd__nor2_1 _17816_ (.A(_02044_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__and2_1 _17817_ (.A(_02044_),
    .B(_02045_),
    .X(_02047_));
 sky130_fd_sc_hd__nor2_1 _17818_ (.A(_02046_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__xnor2_1 _17819_ (.A(_02033_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__a21o_1 _17820_ (.A1(_01961_),
    .A2(_02021_),
    .B1(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__nand3_1 _17821_ (.A(_01961_),
    .B(_02021_),
    .C(_02049_),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _17822_ (.A(_02050_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__xnor2_1 _17823_ (.A(_02020_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__or2_1 _17824_ (.A(_10159_),
    .B(_01967_),
    .X(_02054_));
 sky130_fd_sc_hd__o21ai_1 _17825_ (.A1(_01737_),
    .A2(_02054_),
    .B1(_01858_),
    .Y(_02055_));
 sky130_fd_sc_hd__nor2_1 _17826_ (.A(_10159_),
    .B(_10414_),
    .Y(_02056_));
 sky130_fd_sc_hd__mux2_1 _17827_ (.A0(_10159_),
    .A1(_02056_),
    .S(_01967_),
    .X(_02057_));
 sky130_fd_sc_hd__nand2_1 _17828_ (.A(_01857_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__or2_1 _17829_ (.A(_01857_),
    .B(_02057_),
    .X(_02059_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(_02058_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__xnor2_1 _17831_ (.A(_02055_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__xnor2_1 _17832_ (.A(_01868_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__a21oi_1 _17833_ (.A1(_01868_),
    .A2(_01973_),
    .B1(_01975_),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_1 _17834_ (.A(_02062_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__and2_1 _17835_ (.A(_02062_),
    .B(_02063_),
    .X(_02065_));
 sky130_fd_sc_hd__nor2_1 _17836_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__a21o_1 _17837_ (.A1(_01948_),
    .A2(_01959_),
    .B1(_01957_),
    .X(_02067_));
 sky130_fd_sc_hd__nand2_1 _17838_ (.A(_01857_),
    .B(_01969_),
    .Y(_02068_));
 sky130_fd_sc_hd__or4_1 _17839_ (.A(_10265_),
    .B(_01718_),
    .C(_10163_),
    .D(_09502_),
    .X(_02069_));
 sky130_fd_sc_hd__o22ai_1 _17840_ (.A1(_01718_),
    .A2(_10163_),
    .B1(_09502_),
    .B2(_10265_),
    .Y(_02070_));
 sky130_fd_sc_hd__nand2_1 _17841_ (.A(_02069_),
    .B(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__or3_1 _17842_ (.A(_01834_),
    .B(_10386_),
    .C(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__o21ai_1 _17843_ (.A1(_01834_),
    .A2(_10386_),
    .B1(_02071_),
    .Y(_02073_));
 sky130_fd_sc_hd__and2_1 _17844_ (.A(_02072_),
    .B(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__or2b_1 _17845_ (.A(_08583_),
    .B_N(_09763_),
    .X(_02075_));
 sky130_fd_sc_hd__nor2_1 _17846_ (.A(_08809_),
    .B(_10403_),
    .Y(_02076_));
 sky130_fd_sc_hd__xor2_1 _17847_ (.A(_02075_),
    .B(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__nor2_1 _17848_ (.A(_01729_),
    .B(_10173_),
    .Y(_02078_));
 sky130_fd_sc_hd__xnor2_1 _17849_ (.A(_02077_),
    .B(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__o21ai_1 _17850_ (.A1(_01949_),
    .A2(_01950_),
    .B1(_01952_),
    .Y(_02080_));
 sky130_fd_sc_hd__xor2_1 _17851_ (.A(_02079_),
    .B(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__xnor2_1 _17852_ (.A(_02074_),
    .B(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__a21o_1 _17853_ (.A1(_02068_),
    .A2(_01971_),
    .B1(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__nand3_1 _17854_ (.A(_02068_),
    .B(_01971_),
    .C(_02082_),
    .Y(_02084_));
 sky130_fd_sc_hd__and2_1 _17855_ (.A(_02083_),
    .B(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__nand2_1 _17856_ (.A(_02067_),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__or2_1 _17857_ (.A(_02067_),
    .B(_02085_),
    .X(_02087_));
 sky130_fd_sc_hd__and2_1 _17858_ (.A(_02086_),
    .B(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__xnor2_1 _17859_ (.A(_02066_),
    .B(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__a21oi_1 _17860_ (.A1(_01964_),
    .A2(_01979_),
    .B1(_01977_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _17861_ (.A(_02089_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__and2_1 _17862_ (.A(_02089_),
    .B(_02090_),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_1 _17863_ (.A(_02091_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__xnor2_1 _17864_ (.A(_02053_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__nor2_1 _17865_ (.A(_01980_),
    .B(_01981_),
    .Y(_02095_));
 sky130_fd_sc_hd__a21oi_2 _17866_ (.A1(_01939_),
    .A2(_01982_),
    .B1(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__xor2_1 _17867_ (.A(_02094_),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__xnor2_1 _17868_ (.A(_02019_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_1 _17869_ (.A(_01983_),
    .B(_01985_),
    .Y(_02099_));
 sky130_fd_sc_hd__a21oi_2 _17870_ (.A1(_01905_),
    .A2(_01986_),
    .B1(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_1 _17871_ (.A(_02098_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__and2_1 _17872_ (.A(_02098_),
    .B(_02100_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_1 _17873_ (.A(_02101_),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__xnor2_1 _17874_ (.A(_01903_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__a21o_1 _17875_ (.A1(_01990_),
    .A2(_01993_),
    .B1(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__and3_1 _17876_ (.A(_01990_),
    .B(_01993_),
    .C(_02104_),
    .X(_02106_));
 sky130_fd_sc_hd__inv_2 _17877_ (.A(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand2_1 _17878_ (.A(_02105_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__a21oi_1 _17879_ (.A1(_01997_),
    .A2(_02005_),
    .B1(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__a31o_1 _17880_ (.A1(_01997_),
    .A2(_02005_),
    .A3(_02108_),
    .B1(_08192_),
    .X(_02110_));
 sky130_fd_sc_hd__or2_1 _17881_ (.A(_02109_),
    .B(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__o21ai_1 _17882_ (.A1(_02013_),
    .A2(_02014_),
    .B1(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__mux2_1 _17883_ (.A0(\rbzero.wall_tracer.trackDistX[7] ),
    .A1(_02112_),
    .S(_09917_),
    .X(_02113_));
 sky130_fd_sc_hd__clkbuf_1 _17884_ (.A(_02113_),
    .X(_00546_));
 sky130_fd_sc_hd__or2b_1 _17885_ (.A(_02052_),
    .B_N(_02020_),
    .X(_02114_));
 sky130_fd_sc_hd__o22a_1 _17886_ (.A1(_02029_),
    .A2(_02030_),
    .B1(_02031_),
    .B2(_02032_),
    .X(_02115_));
 sky130_fd_sc_hd__a21o_1 _17887_ (.A1(_02050_),
    .A2(_02114_),
    .B1(_02115_),
    .X(_02116_));
 sky130_fd_sc_hd__nand3_1 _17888_ (.A(_02050_),
    .B(_02114_),
    .C(_02115_),
    .Y(_02117_));
 sky130_fd_sc_hd__and2_1 _17889_ (.A(_02116_),
    .B(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__a21o_1 _17890_ (.A1(_01868_),
    .A2(_02061_),
    .B1(_01975_),
    .X(_02119_));
 sky130_fd_sc_hd__nand2_1 _17891_ (.A(_01858_),
    .B(_02054_),
    .Y(_02120_));
 sky130_fd_sc_hd__xnor2_2 _17892_ (.A(_02060_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__xor2_1 _17893_ (.A(_01868_),
    .B(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__and2_1 _17894_ (.A(_02119_),
    .B(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__nor2_1 _17895_ (.A(_02119_),
    .B(_02122_),
    .Y(_02124_));
 sky130_fd_sc_hd__nor2_1 _17896_ (.A(_02123_),
    .B(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__and2_1 _17897_ (.A(_02079_),
    .B(_02080_),
    .X(_02126_));
 sky130_fd_sc_hd__a21o_1 _17898_ (.A1(_02074_),
    .A2(_02081_),
    .B1(_02126_),
    .X(_02127_));
 sky130_fd_sc_hd__a21bo_1 _17899_ (.A1(_02055_),
    .A2(_02059_),
    .B1_N(_02058_),
    .X(_02128_));
 sky130_fd_sc_hd__nor2_1 _17900_ (.A(_01718_),
    .B(_09502_),
    .Y(_02129_));
 sky130_fd_sc_hd__nor2_1 _17901_ (.A(_10265_),
    .B(_09515_),
    .Y(_02130_));
 sky130_fd_sc_hd__xnor2_1 _17902_ (.A(_02129_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__or3_1 _17903_ (.A(_10386_),
    .B(_10163_),
    .C(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__o21ai_1 _17904_ (.A1(_10386_),
    .A2(_10163_),
    .B1(_02131_),
    .Y(_02133_));
 sky130_fd_sc_hd__and2_1 _17905_ (.A(_02132_),
    .B(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__or3_1 _17906_ (.A(_08809_),
    .B(_08583_),
    .C(_10414_),
    .X(_02135_));
 sky130_fd_sc_hd__o22a_1 _17907_ (.A1(_08809_),
    .A2(_10414_),
    .B1(_10403_),
    .B2(_08583_),
    .X(_02136_));
 sky130_fd_sc_hd__o21ba_1 _17908_ (.A1(_01737_),
    .A2(_02135_),
    .B1_N(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__and2b_1 _17909_ (.A_N(_09358_),
    .B(_09763_),
    .X(_02138_));
 sky130_fd_sc_hd__nand2_1 _17910_ (.A(_02137_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__or2_1 _17911_ (.A(_02137_),
    .B(_02138_),
    .X(_02140_));
 sky130_fd_sc_hd__nand2_1 _17912_ (.A(_02139_),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__or3_1 _17913_ (.A(_01729_),
    .B(_10173_),
    .C(_02077_),
    .X(_02142_));
 sky130_fd_sc_hd__o31a_1 _17914_ (.A1(_08809_),
    .A2(_01737_),
    .A3(_02075_),
    .B1(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__xor2_1 _17915_ (.A(_02141_),
    .B(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__nand2_1 _17916_ (.A(_02134_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__or2_1 _17917_ (.A(_02134_),
    .B(_02144_),
    .X(_02146_));
 sky130_fd_sc_hd__and2_1 _17918_ (.A(_02145_),
    .B(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__xnor2_1 _17919_ (.A(_02128_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__xnor2_1 _17920_ (.A(_02127_),
    .B(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__xnor2_1 _17921_ (.A(_02125_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__a21oi_1 _17922_ (.A1(_02066_),
    .A2(_02088_),
    .B1(_02064_),
    .Y(_02151_));
 sky130_fd_sc_hd__xor2_1 _17923_ (.A(_02150_),
    .B(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__a21o_1 _17924_ (.A1(_02033_),
    .A2(_02048_),
    .B1(_02046_),
    .X(_02153_));
 sky130_fd_sc_hd__or2_2 _17925_ (.A(_08303_),
    .B(_09314_),
    .X(_02154_));
 sky130_fd_sc_hd__or2b_1 _17926_ (.A(_09441_),
    .B_N(_08228_),
    .X(_02155_));
 sky130_fd_sc_hd__xnor2_2 _17927_ (.A(_02154_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__nor2_1 _17928_ (.A(_10262_),
    .B(_09706_),
    .Y(_02157_));
 sky130_fd_sc_hd__xor2_2 _17929_ (.A(_02156_),
    .B(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__o31a_1 _17930_ (.A1(_10144_),
    .A2(_09706_),
    .A3(_02027_),
    .B1(_02025_),
    .X(_02159_));
 sky130_fd_sc_hd__xor2_2 _17931_ (.A(_02158_),
    .B(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__and2_1 _17932_ (.A(_10144_),
    .B(_09691_),
    .X(_02161_));
 sky130_fd_sc_hd__xor2_2 _17933_ (.A(_02160_),
    .B(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__a21bo_1 _17934_ (.A1(_02038_),
    .A2(_02039_),
    .B1_N(_02036_),
    .X(_02163_));
 sky130_fd_sc_hd__nor2_1 _17935_ (.A(_01716_),
    .B(_01810_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _17936_ (.A(_01834_),
    .B(_01692_),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_1 _17937_ (.A(_02164_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__or3_1 _17938_ (.A(_08336_),
    .B(_01919_),
    .C(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__o21ai_1 _17939_ (.A1(_08336_),
    .A2(_01919_),
    .B1(_02166_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _17940_ (.A(_02167_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__a21o_1 _17941_ (.A1(_02069_),
    .A2(_02072_),
    .B1(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__nand3_1 _17942_ (.A(_02069_),
    .B(_02072_),
    .C(_02169_),
    .Y(_02171_));
 sky130_fd_sc_hd__nand2_1 _17943_ (.A(_02170_),
    .B(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__xor2_1 _17944_ (.A(_02163_),
    .B(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__a21oi_1 _17945_ (.A1(_02034_),
    .A2(_02043_),
    .B1(_02041_),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_1 _17946_ (.A(_02173_),
    .B(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__and2_1 _17947_ (.A(_02173_),
    .B(_02174_),
    .X(_02176_));
 sky130_fd_sc_hd__nor2_1 _17948_ (.A(_02175_),
    .B(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__xnor2_1 _17949_ (.A(_02162_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__a21o_1 _17950_ (.A1(_02083_),
    .A2(_02086_),
    .B1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__nand3_1 _17951_ (.A(_02083_),
    .B(_02086_),
    .C(_02178_),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_1 _17952_ (.A(_02179_),
    .B(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__xnor2_1 _17953_ (.A(_02153_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_1 _17954_ (.A(_02152_),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__or2_1 _17955_ (.A(_02152_),
    .B(_02182_),
    .X(_02184_));
 sky130_fd_sc_hd__nand2_1 _17956_ (.A(_02183_),
    .B(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__a21oi_1 _17957_ (.A1(_02053_),
    .A2(_02093_),
    .B1(_02091_),
    .Y(_02186_));
 sky130_fd_sc_hd__xor2_1 _17958_ (.A(_02185_),
    .B(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__nand2_1 _17959_ (.A(_02118_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__or2_1 _17960_ (.A(_02118_),
    .B(_02187_),
    .X(_02189_));
 sky130_fd_sc_hd__nand2_1 _17961_ (.A(_02188_),
    .B(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__nor2_1 _17962_ (.A(_02094_),
    .B(_02096_),
    .Y(_02191_));
 sky130_fd_sc_hd__a21oi_1 _17963_ (.A1(_02019_),
    .A2(_02097_),
    .B1(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__xor2_1 _17964_ (.A(_02190_),
    .B(_02192_),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_1 _17965_ (.A(_02017_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__a21oi_1 _17966_ (.A1(_01903_),
    .A2(_02103_),
    .B1(_02101_),
    .Y(_02195_));
 sky130_fd_sc_hd__or2_1 _17967_ (.A(_02194_),
    .B(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__nand2_1 _17968_ (.A(_02194_),
    .B(_02195_),
    .Y(_02197_));
 sky130_fd_sc_hd__and2_1 _17969_ (.A(_02196_),
    .B(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__inv_2 _17970_ (.A(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__a311o_2 _17971_ (.A1(_01997_),
    .A2(_02005_),
    .A3(_02105_),
    .B1(_02106_),
    .C1(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__a31o_1 _17972_ (.A1(_01997_),
    .A2(_02005_),
    .A3(_02105_),
    .B1(_02106_),
    .X(_02201_));
 sky130_fd_sc_hd__a21oi_1 _17973_ (.A1(_02199_),
    .A2(_02201_),
    .B1(_08195_),
    .Y(_02202_));
 sky130_fd_sc_hd__nand2_1 _17974_ (.A(_02200_),
    .B(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__or2_1 _17975_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .X(_02204_));
 sky130_fd_sc_hd__nand2_1 _17976_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _17977_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__o21ai_1 _17978_ (.A1(_02009_),
    .A2(_02012_),
    .B1(_02010_),
    .Y(_02207_));
 sky130_fd_sc_hd__xnor2_1 _17979_ (.A(_02206_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__a21oi_1 _17980_ (.A1(_08195_),
    .A2(_02208_),
    .B1(_09859_),
    .Y(_02209_));
 sky130_fd_sc_hd__o2bb2a_1 _17981_ (.A1_N(_02203_),
    .A2_N(_02209_),
    .B1(\rbzero.wall_tracer.trackDistX[8] ),
    .B2(_09884_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _17982_ (.A(_02190_),
    .B(_02192_),
    .X(_02210_));
 sky130_fd_sc_hd__nand2_1 _17983_ (.A(_02017_),
    .B(_02193_),
    .Y(_02211_));
 sky130_fd_sc_hd__a21o_1 _17984_ (.A1(_02125_),
    .A2(_02149_),
    .B1(_02123_),
    .X(_02212_));
 sky130_fd_sc_hd__o21ai_1 _17985_ (.A1(_02141_),
    .A2(_02143_),
    .B1(_02145_),
    .Y(_02213_));
 sky130_fd_sc_hd__a21bo_1 _17986_ (.A1(_02059_),
    .A2(_02120_),
    .B1_N(_02058_),
    .X(_02214_));
 sky130_fd_sc_hd__nor2_1 _17987_ (.A(_01718_),
    .B(_09515_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _17988_ (.A(_08495_),
    .B(_09507_),
    .Y(_02216_));
 sky130_fd_sc_hd__xnor2_1 _17989_ (.A(_02215_),
    .B(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__nor2_1 _17990_ (.A(_10386_),
    .B(_09502_),
    .Y(_02218_));
 sky130_fd_sc_hd__xnor2_1 _17991_ (.A(_02217_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__or2_1 _17992_ (.A(_01737_),
    .B(_02135_),
    .X(_02220_));
 sky130_fd_sc_hd__a21oi_1 _17993_ (.A1(_08809_),
    .A2(_08583_),
    .B1(_10414_),
    .Y(_02221_));
 sky130_fd_sc_hd__o211a_1 _17994_ (.A1(_01729_),
    .A2(_01737_),
    .B1(_02135_),
    .C1(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__a211oi_1 _17995_ (.A1(_02135_),
    .A2(_02221_),
    .B1(_01729_),
    .C1(_01737_),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _17996_ (.A(_02222_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__a21oi_1 _17997_ (.A1(_02220_),
    .A2(_02139_),
    .B1(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__and3_1 _17998_ (.A(_02220_),
    .B(_02139_),
    .C(_02224_),
    .X(_02226_));
 sky130_fd_sc_hd__nor2_1 _17999_ (.A(_02225_),
    .B(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__xor2_1 _18000_ (.A(_02219_),
    .B(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__and2_1 _18001_ (.A(_02214_),
    .B(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__nor2_1 _18002_ (.A(_02214_),
    .B(_02228_),
    .Y(_02230_));
 sky130_fd_sc_hd__nor2_1 _18003_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_02213_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__mux2_1 _18005_ (.A0(_01866_),
    .A1(_01865_),
    .S(_02121_),
    .X(_02233_));
 sky130_fd_sc_hd__xnor2_1 _18006_ (.A(_02232_),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__xnor2_1 _18007_ (.A(_02212_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__a21o_1 _18008_ (.A1(_02162_),
    .A2(_02177_),
    .B1(_02175_),
    .X(_02236_));
 sky130_fd_sc_hd__or2b_1 _18009_ (.A(_02148_),
    .B_N(_02127_),
    .X(_02237_));
 sky130_fd_sc_hd__a21bo_1 _18010_ (.A1(_02128_),
    .A2(_02147_),
    .B1_N(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__nand2_1 _18011_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08340_),
    .Y(_02239_));
 sky130_fd_sc_hd__a22o_1 _18012_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_08339_),
    .B1(_08340_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_02240_));
 sky130_fd_sc_hd__o21ai_2 _18013_ (.A1(_02154_),
    .A2(_02239_),
    .B1(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__and3_1 _18014_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_08496_),
    .C(_08228_),
    .X(_02242_));
 sky130_fd_sc_hd__xor2_2 _18015_ (.A(_02241_),
    .B(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__or2_1 _18016_ (.A(_02154_),
    .B(_02155_),
    .X(_02244_));
 sky130_fd_sc_hd__o31a_1 _18017_ (.A1(_10262_),
    .A2(_09706_),
    .A3(_02156_),
    .B1(_02244_),
    .X(_02245_));
 sky130_fd_sc_hd__xor2_2 _18018_ (.A(_02243_),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__and2_1 _18019_ (.A(_10262_),
    .B(_09691_),
    .X(_02247_));
 sky130_fd_sc_hd__xor2_2 _18020_ (.A(_02246_),
    .B(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__or2b_1 _18021_ (.A(_02172_),
    .B_N(_02163_),
    .X(_02249_));
 sky130_fd_sc_hd__a21bo_1 _18022_ (.A1(_02164_),
    .A2(_02165_),
    .B1_N(_02167_),
    .X(_02250_));
 sky130_fd_sc_hd__a21bo_1 _18023_ (.A1(_02129_),
    .A2(_02130_),
    .B1_N(_02132_),
    .X(_02251_));
 sky130_fd_sc_hd__or4_1 _18024_ (.A(_01834_),
    .B(_01692_),
    .C(_10163_),
    .D(_01810_),
    .X(_02252_));
 sky130_fd_sc_hd__o22ai_1 _18025_ (.A1(_01692_),
    .A2(_10163_),
    .B1(_01810_),
    .B2(_01834_),
    .Y(_02253_));
 sky130_fd_sc_hd__and2_1 _18026_ (.A(_02252_),
    .B(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__nor2_1 _18027_ (.A(_01716_),
    .B(_01919_),
    .Y(_02255_));
 sky130_fd_sc_hd__xor2_1 _18028_ (.A(_02254_),
    .B(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__and2_1 _18029_ (.A(_02251_),
    .B(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__or2_1 _18030_ (.A(_02251_),
    .B(_02256_),
    .X(_02258_));
 sky130_fd_sc_hd__and2b_1 _18031_ (.A_N(_02257_),
    .B(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__xnor2_1 _18032_ (.A(_02250_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__a21oi_1 _18033_ (.A1(_02170_),
    .A2(_02249_),
    .B1(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__and3_1 _18034_ (.A(_02170_),
    .B(_02249_),
    .C(_02260_),
    .X(_02262_));
 sky130_fd_sc_hd__nor2_1 _18035_ (.A(_02261_),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__xor2_1 _18036_ (.A(_02248_),
    .B(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__xor2_1 _18037_ (.A(_02238_),
    .B(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__and2_1 _18038_ (.A(_02236_),
    .B(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__nor2_1 _18039_ (.A(_02236_),
    .B(_02265_),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _18040_ (.A(_02266_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__xor2_1 _18041_ (.A(_02235_),
    .B(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__o21a_1 _18042_ (.A1(_02150_),
    .A2(_02151_),
    .B1(_02183_),
    .X(_02270_));
 sky130_fd_sc_hd__xnor2_1 _18043_ (.A(_02269_),
    .B(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hd__or2b_1 _18044_ (.A(_02181_),
    .B_N(_02153_),
    .X(_02272_));
 sky130_fd_sc_hd__o2bb2a_1 _18045_ (.A1_N(_02160_),
    .A2_N(_02161_),
    .B1(_02158_),
    .B2(_02159_),
    .X(_02273_));
 sky130_fd_sc_hd__a21oi_1 _18046_ (.A1(_02179_),
    .A2(_02272_),
    .B1(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__and3_1 _18047_ (.A(_02179_),
    .B(_02272_),
    .C(_02273_),
    .X(_02275_));
 sky130_fd_sc_hd__nor2_1 _18048_ (.A(_02274_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__xor2_1 _18049_ (.A(_02271_),
    .B(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__o21a_1 _18050_ (.A1(_02185_),
    .A2(_02186_),
    .B1(_02188_),
    .X(_02278_));
 sky130_fd_sc_hd__xor2_1 _18051_ (.A(_02277_),
    .B(_02278_),
    .X(_02279_));
 sky130_fd_sc_hd__xor2_1 _18052_ (.A(_02116_),
    .B(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__a21o_1 _18053_ (.A1(_02210_),
    .A2(_02211_),
    .B1(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__inv_2 _18054_ (.A(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__and3_1 _18055_ (.A(_02210_),
    .B(_02211_),
    .C(_02280_),
    .X(_02283_));
 sky130_fd_sc_hd__nor2_1 _18056_ (.A(_02282_),
    .B(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__inv_2 _18057_ (.A(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__a21oi_1 _18058_ (.A1(_02196_),
    .A2(_02200_),
    .B1(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__a31o_1 _18059_ (.A1(_02196_),
    .A2(_02200_),
    .A3(_02285_),
    .B1(_08194_),
    .X(_02287_));
 sky130_fd_sc_hd__or2_1 _18060_ (.A(_02286_),
    .B(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__nand2_1 _18061_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_02289_));
 sky130_fd_sc_hd__or2_1 _18062_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_02290_));
 sky130_fd_sc_hd__nand2_1 _18063_ (.A(_02289_),
    .B(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__a21bo_1 _18064_ (.A1(_02204_),
    .A2(_02207_),
    .B1_N(_02205_),
    .X(_02292_));
 sky130_fd_sc_hd__xnor2_1 _18065_ (.A(_02291_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__a21oi_1 _18066_ (.A1(_08195_),
    .A2(_02293_),
    .B1(_09859_),
    .Y(_02294_));
 sky130_fd_sc_hd__o2bb2a_1 _18067_ (.A1_N(_02288_),
    .A2_N(_02294_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_09884_),
    .X(_00548_));
 sky130_fd_sc_hd__a21o_1 _18068_ (.A1(_02196_),
    .A2(_02281_),
    .B1(_02283_),
    .X(_02295_));
 sky130_fd_sc_hd__or2b_1 _18069_ (.A(_02116_),
    .B_N(_02279_),
    .X(_02296_));
 sky130_fd_sc_hd__o21ai_1 _18070_ (.A1(_02277_),
    .A2(_02278_),
    .B1(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__or2_1 _18071_ (.A(_01866_),
    .B(_02121_),
    .X(_02298_));
 sky130_fd_sc_hd__a22o_1 _18072_ (.A1(_01975_),
    .A2(_02121_),
    .B1(_02298_),
    .B2(_02232_),
    .X(_02299_));
 sky130_fd_sc_hd__xnor2_1 _18073_ (.A(_02214_),
    .B(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__xnor2_1 _18074_ (.A(_02274_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__a21o_1 _18075_ (.A1(_02219_),
    .A2(_02227_),
    .B1(_02225_),
    .X(_02302_));
 sky130_fd_sc_hd__nor2_1 _18076_ (.A(_10386_),
    .B(_09515_),
    .Y(_02303_));
 sky130_fd_sc_hd__xnor2_1 _18077_ (.A(_02302_),
    .B(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__or2_1 _18078_ (.A(_01729_),
    .B(_10414_),
    .X(_02305_));
 sky130_fd_sc_hd__nand2_1 _18079_ (.A(_06340_),
    .B(_09510_),
    .Y(_02306_));
 sky130_fd_sc_hd__o22ai_1 _18080_ (.A1(_01718_),
    .A2(_02306_),
    .B1(_10053_),
    .B2(_10265_),
    .Y(_02307_));
 sky130_fd_sc_hd__o41a_1 _18081_ (.A1(_08495_),
    .A2(_01718_),
    .A3(_02306_),
    .A4(_09773_),
    .B1(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__xnor2_1 _18082_ (.A(_02305_),
    .B(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__a21oi_1 _18083_ (.A1(_02250_),
    .A2(_02259_),
    .B1(_02257_),
    .Y(_02310_));
 sky130_fd_sc_hd__or2_1 _18084_ (.A(_10163_),
    .B(_01810_),
    .X(_02311_));
 sky130_fd_sc_hd__nor2_1 _18085_ (.A(_08228_),
    .B(_09687_),
    .Y(_02312_));
 sky130_fd_sc_hd__xnor2_1 _18086_ (.A(_02311_),
    .B(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__xnor2_1 _18087_ (.A(_02310_),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__a21o_1 _18088_ (.A1(_02248_),
    .A2(_02263_),
    .B1(_02261_),
    .X(_02315_));
 sky130_fd_sc_hd__nor2_1 _18089_ (.A(_01692_),
    .B(_09502_),
    .Y(_02316_));
 sky130_fd_sc_hd__xnor2_1 _18090_ (.A(_02315_),
    .B(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__xnor2_1 _18091_ (.A(_02314_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__xnor2_1 _18092_ (.A(_02309_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _18093_ (.A(_02215_),
    .B(_02216_),
    .Y(_02320_));
 sky130_fd_sc_hd__o31a_1 _18094_ (.A1(_10386_),
    .A2(_09502_),
    .A3(_02217_),
    .B1(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__or2b_1 _18095_ (.A(_02241_),
    .B_N(_02242_),
    .X(_02322_));
 sky130_fd_sc_hd__o21ai_1 _18096_ (.A1(_02154_),
    .A2(_02239_),
    .B1(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__nor2_1 _18097_ (.A(_01716_),
    .B(_02023_),
    .Y(_02324_));
 sky130_fd_sc_hd__nor2_1 _18098_ (.A(_08303_),
    .B(_09706_),
    .Y(_02325_));
 sky130_fd_sc_hd__xnor2_1 _18099_ (.A(_02239_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__xnor2_1 _18100_ (.A(_02324_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__xnor2_1 _18101_ (.A(_02323_),
    .B(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__a21boi_1 _18102_ (.A1(_02253_),
    .A2(_02255_),
    .B1_N(_02252_),
    .Y(_02329_));
 sky130_fd_sc_hd__nor2_1 _18103_ (.A(_01834_),
    .B(_01919_),
    .Y(_02330_));
 sky130_fd_sc_hd__xor2_1 _18104_ (.A(_02329_),
    .B(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__xnor2_1 _18105_ (.A(_02328_),
    .B(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__xnor2_1 _18106_ (.A(_02321_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__a21oi_1 _18107_ (.A1(_02213_),
    .A2(_02231_),
    .B1(_02229_),
    .Y(_02334_));
 sky130_fd_sc_hd__xnor2_1 _18108_ (.A(_02333_),
    .B(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__xnor2_1 _18109_ (.A(_02319_),
    .B(_02335_),
    .Y(_02336_));
 sky130_fd_sc_hd__xnor2_1 _18110_ (.A(_02304_),
    .B(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__xnor2_1 _18111_ (.A(_02301_),
    .B(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__o21ai_1 _18112_ (.A1(_01729_),
    .A2(_01737_),
    .B1(_02221_),
    .Y(_02339_));
 sky130_fd_sc_hd__nand2_1 _18113_ (.A(_02135_),
    .B(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__and2b_1 _18114_ (.A_N(_02235_),
    .B(_02268_),
    .X(_02341_));
 sky130_fd_sc_hd__a21oi_1 _18115_ (.A1(_02212_),
    .A2(_02234_),
    .B1(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__a21oi_1 _18116_ (.A1(_02238_),
    .A2(_02264_),
    .B1(_02266_),
    .Y(_02343_));
 sky130_fd_sc_hd__xnor2_1 _18117_ (.A(_02342_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__xor2_1 _18118_ (.A(_02340_),
    .B(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__xnor2_1 _18119_ (.A(_02338_),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__or2b_1 _18120_ (.A(_02271_),
    .B_N(_02276_),
    .X(_02347_));
 sky130_fd_sc_hd__o21a_1 _18121_ (.A1(_02269_),
    .A2(_02270_),
    .B1(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__a2bb2o_1 _18122_ (.A1_N(_02243_),
    .A2_N(_02245_),
    .B1(_02246_),
    .B2(_02247_),
    .X(_02349_));
 sky130_fd_sc_hd__xnor2_1 _18123_ (.A(_02348_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__xnor2_1 _18124_ (.A(_02346_),
    .B(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__xnor2_1 _18125_ (.A(_02297_),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__o211a_1 _18126_ (.A1(_02200_),
    .A2(_02285_),
    .B1(_02295_),
    .C1(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__a311o_1 _18127_ (.A1(_02196_),
    .A2(_02200_),
    .A3(_02281_),
    .B1(_02283_),
    .C1(_02352_),
    .X(_02354_));
 sky130_fd_sc_hd__or3b_1 _18128_ (.A(_08194_),
    .B(_02353_),
    .C_N(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__a21bo_1 _18129_ (.A1(_02290_),
    .A2(_02292_),
    .B1_N(_02289_),
    .X(_02356_));
 sky130_fd_sc_hd__xor2_1 _18130_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .X(_02357_));
 sky130_fd_sc_hd__xnor2_1 _18131_ (.A(_02356_),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__o21a_1 _18132_ (.A1(_08156_),
    .A2(_02358_),
    .B1(_09883_),
    .X(_02359_));
 sky130_fd_sc_hd__o2bb2a_1 _18133_ (.A1_N(_02355_),
    .A2_N(_02359_),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_09884_),
    .X(_00549_));
 sky130_fd_sc_hd__and2_1 _18134_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_02360_));
 sky130_fd_sc_hd__nor2_1 _18135_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_02361_));
 sky130_fd_sc_hd__a221oi_4 _18136_ (.A1(_06237_),
    .A2(_06331_),
    .B1(_08321_),
    .B2(_06334_),
    .C1(_06341_),
    .Y(_02362_));
 sky130_fd_sc_hd__clkbuf_4 _18137_ (.A(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__o31a_1 _18138_ (.A1(_01779_),
    .A2(_02360_),
    .A3(_02361_),
    .B1(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__clkbuf_4 _18139_ (.A(_02362_),
    .X(_02365_));
 sky130_fd_sc_hd__o2bb2a_1 _18140_ (.A1_N(_09878_),
    .A2_N(_02364_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-11] ),
    .X(_00550_));
 sky130_fd_sc_hd__or2_1 _18141_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_02366_));
 sky130_fd_sc_hd__nand2_1 _18142_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_02367_));
 sky130_fd_sc_hd__and4_1 _18143_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .C(_02366_),
    .D(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__a22oi_1 _18144_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(\rbzero.wall_tracer.stepDistY[-11] ),
    .B1(_02366_),
    .B2(_02367_),
    .Y(_02369_));
 sky130_fd_sc_hd__buf_4 _18145_ (.A(_02362_),
    .X(_02370_));
 sky130_fd_sc_hd__o31a_1 _18146_ (.A1(_01779_),
    .A2(_02368_),
    .A3(_02369_),
    .B1(_02370_),
    .X(_02371_));
 sky130_fd_sc_hd__o2bb2a_1 _18147_ (.A1_N(_09887_),
    .A2_N(_02371_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(_00551_));
 sky130_fd_sc_hd__a21o_1 _18148_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(\rbzero.wall_tracer.stepDistY[-10] ),
    .B1(_02368_),
    .X(_02372_));
 sky130_fd_sc_hd__or2_1 _18149_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_02373_));
 sky130_fd_sc_hd__nand2_1 _18150_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_02374_));
 sky130_fd_sc_hd__and3_1 _18151_ (.A(_02372_),
    .B(_02373_),
    .C(_02374_),
    .X(_02375_));
 sky130_fd_sc_hd__a21oi_1 _18152_ (.A1(_02373_),
    .A2(_02374_),
    .B1(_02372_),
    .Y(_02376_));
 sky130_fd_sc_hd__o31a_1 _18153_ (.A1(_01779_),
    .A2(_02375_),
    .A3(_02376_),
    .B1(_02370_),
    .X(_02377_));
 sky130_fd_sc_hd__o2bb2a_1 _18154_ (.A1_N(_09898_),
    .A2_N(_02377_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(_00552_));
 sky130_fd_sc_hd__or2_1 _18155_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_02378_));
 sky130_fd_sc_hd__nand2_1 _18156_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .Y(_02379_));
 sky130_fd_sc_hd__a21bo_1 _18157_ (.A1(_02372_),
    .A2(_02373_),
    .B1_N(_02374_),
    .X(_02380_));
 sky130_fd_sc_hd__and3_1 _18158_ (.A(_02378_),
    .B(_02379_),
    .C(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__a21oi_1 _18159_ (.A1(_02378_),
    .A2(_02379_),
    .B1(_02380_),
    .Y(_02382_));
 sky130_fd_sc_hd__o31a_1 _18160_ (.A1(_01779_),
    .A2(_02381_),
    .A3(_02382_),
    .B1(_02370_),
    .X(_02383_));
 sky130_fd_sc_hd__o2bb2a_1 _18161_ (.A1_N(_09906_),
    .A2_N(_02383_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-8] ),
    .X(_00553_));
 sky130_fd_sc_hd__nor2_1 _18162_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _18163_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02385_));
 sky130_fd_sc_hd__or2b_1 _18164_ (.A(_02384_),
    .B_N(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__a21boi_1 _18165_ (.A1(_02378_),
    .A2(_02380_),
    .B1_N(_02379_),
    .Y(_02387_));
 sky130_fd_sc_hd__xnor2_1 _18166_ (.A(_02386_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__o21a_1 _18167_ (.A1(_08156_),
    .A2(_02388_),
    .B1(_02363_),
    .X(_02389_));
 sky130_fd_sc_hd__o2bb2a_1 _18168_ (.A1_N(_09915_),
    .A2_N(_02389_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-7] ),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _18169_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_02390_));
 sky130_fd_sc_hd__nand2_1 _18170_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .Y(_02391_));
 sky130_fd_sc_hd__o21ai_1 _18171_ (.A1(_02384_),
    .A2(_02387_),
    .B1(_02385_),
    .Y(_02392_));
 sky130_fd_sc_hd__and3_1 _18172_ (.A(_02390_),
    .B(_02391_),
    .C(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__a21oi_1 _18173_ (.A1(_02390_),
    .A2(_02391_),
    .B1(_02392_),
    .Y(_02394_));
 sky130_fd_sc_hd__o31a_1 _18174_ (.A1(_01779_),
    .A2(_02393_),
    .A3(_02394_),
    .B1(_02370_),
    .X(_02395_));
 sky130_fd_sc_hd__o2bb2a_1 _18175_ (.A1_N(_09924_),
    .A2_N(_02395_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(_00555_));
 sky130_fd_sc_hd__nor2_1 _18176_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02396_));
 sky130_fd_sc_hd__nand2_1 _18177_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02397_));
 sky130_fd_sc_hd__or2b_1 _18178_ (.A(_02396_),
    .B_N(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__a21boi_1 _18179_ (.A1(_02390_),
    .A2(_02392_),
    .B1_N(_02391_),
    .Y(_02399_));
 sky130_fd_sc_hd__nor2_1 _18180_ (.A(_02398_),
    .B(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__a21o_1 _18181_ (.A1(_02398_),
    .A2(_02399_),
    .B1(_06163_),
    .X(_02401_));
 sky130_fd_sc_hd__o21ai_1 _18182_ (.A1(_02400_),
    .A2(_02401_),
    .B1(_09927_),
    .Y(_02402_));
 sky130_fd_sc_hd__mux2_1 _18183_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(_02402_),
    .S(_02362_),
    .X(_02403_));
 sky130_fd_sc_hd__clkbuf_1 _18184_ (.A(_02403_),
    .X(_00556_));
 sky130_fd_sc_hd__or2_1 _18185_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(_02404_));
 sky130_fd_sc_hd__nand2_1 _18186_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02405_));
 sky130_fd_sc_hd__o21ai_1 _18187_ (.A1(_02396_),
    .A2(_02399_),
    .B1(_02397_),
    .Y(_02406_));
 sky130_fd_sc_hd__and3_1 _18188_ (.A(_02404_),
    .B(_02405_),
    .C(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__a21oi_1 _18189_ (.A1(_02404_),
    .A2(_02405_),
    .B1(_02406_),
    .Y(_02408_));
 sky130_fd_sc_hd__o31a_1 _18190_ (.A1(_01779_),
    .A2(_02407_),
    .A3(_02408_),
    .B1(_02370_),
    .X(_02409_));
 sky130_fd_sc_hd__o2bb2a_1 _18191_ (.A1_N(_09934_),
    .A2_N(_02409_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-4] ),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _18192_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_1 _18193_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02411_));
 sky130_fd_sc_hd__or2b_1 _18194_ (.A(_02410_),
    .B_N(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__a21boi_1 _18195_ (.A1(_02404_),
    .A2(_02406_),
    .B1_N(_02405_),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _18196_ (.A(_02412_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__a21o_1 _18197_ (.A1(_02412_),
    .A2(_02413_),
    .B1(_06163_),
    .X(_02415_));
 sky130_fd_sc_hd__o21ai_1 _18198_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_09948_),
    .Y(_02416_));
 sky130_fd_sc_hd__mux2_1 _18199_ (.A0(\rbzero.wall_tracer.trackDistY[-3] ),
    .A1(_02416_),
    .S(_02362_),
    .X(_02417_));
 sky130_fd_sc_hd__clkbuf_1 _18200_ (.A(_02417_),
    .X(_00558_));
 sky130_fd_sc_hd__or2_1 _18201_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_1 _18202_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02419_));
 sky130_fd_sc_hd__o21ai_1 _18203_ (.A1(_02410_),
    .A2(_02413_),
    .B1(_02411_),
    .Y(_02420_));
 sky130_fd_sc_hd__and3_1 _18204_ (.A(_02418_),
    .B(_02419_),
    .C(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__a21oi_1 _18205_ (.A1(_02418_),
    .A2(_02419_),
    .B1(_02420_),
    .Y(_02422_));
 sky130_fd_sc_hd__o31a_1 _18206_ (.A1(_01779_),
    .A2(_02421_),
    .A3(_02422_),
    .B1(_02370_),
    .X(_02423_));
 sky130_fd_sc_hd__o2bb2a_1 _18207_ (.A1_N(_09956_),
    .A2_N(_02423_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_00559_));
 sky130_fd_sc_hd__nor2_1 _18208_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_02424_));
 sky130_fd_sc_hd__and2_1 _18209_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .X(_02425_));
 sky130_fd_sc_hd__or2_1 _18210_ (.A(_02424_),
    .B(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__a21boi_1 _18211_ (.A1(_02418_),
    .A2(_02420_),
    .B1_N(_02419_),
    .Y(_02427_));
 sky130_fd_sc_hd__nor2_1 _18212_ (.A(_02426_),
    .B(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__a21o_1 _18213_ (.A1(_02426_),
    .A2(_02427_),
    .B1(_06163_),
    .X(_02429_));
 sky130_fd_sc_hd__o21ai_1 _18214_ (.A1(_02428_),
    .A2(_02429_),
    .B1(_09964_),
    .Y(_02430_));
 sky130_fd_sc_hd__mux2_1 _18215_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(_02430_),
    .S(_02362_),
    .X(_02431_));
 sky130_fd_sc_hd__clkbuf_1 _18216_ (.A(_02431_),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _18217_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .X(_02432_));
 sky130_fd_sc_hd__nand2_1 _18218_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_02433_));
 sky130_fd_sc_hd__a211oi_1 _18219_ (.A1(_02432_),
    .A2(_02433_),
    .B1(_02425_),
    .C1(_02428_),
    .Y(_02434_));
 sky130_fd_sc_hd__o211a_1 _18220_ (.A1(_02425_),
    .A2(_02428_),
    .B1(_02432_),
    .C1(_02433_),
    .X(_02435_));
 sky130_fd_sc_hd__o31a_1 _18221_ (.A1(_01779_),
    .A2(_02434_),
    .A3(_02435_),
    .B1(_02370_),
    .X(_02436_));
 sky130_fd_sc_hd__o2bb2a_1 _18222_ (.A1_N(_10093_),
    .A2_N(_02436_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[0] ),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_1 _18223_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_02437_));
 sky130_fd_sc_hd__or2_1 _18224_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_02438_));
 sky130_fd_sc_hd__a21o_1 _18225_ (.A1(\rbzero.wall_tracer.trackDistY[0] ),
    .A2(\rbzero.wall_tracer.stepDistY[0] ),
    .B1(_02435_),
    .X(_02439_));
 sky130_fd_sc_hd__and3_1 _18226_ (.A(_02437_),
    .B(_02438_),
    .C(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__a21o_1 _18227_ (.A1(_02437_),
    .A2(_02438_),
    .B1(_02439_),
    .X(_02441_));
 sky130_fd_sc_hd__or3b_1 _18228_ (.A(_06163_),
    .B(_02440_),
    .C_N(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__nand2_1 _18229_ (.A(_10212_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__mux2_1 _18230_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(_02443_),
    .S(_02362_),
    .X(_02444_));
 sky130_fd_sc_hd__clkbuf_1 _18231_ (.A(_02444_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _18232_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_02445_));
 sky130_fd_sc_hd__or2_1 _18233_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_02446_));
 sky130_fd_sc_hd__inv_2 _18234_ (.A(_02437_),
    .Y(_02447_));
 sky130_fd_sc_hd__a211o_1 _18235_ (.A1(_02445_),
    .A2(_02446_),
    .B1(_02447_),
    .C1(_02440_),
    .X(_02448_));
 sky130_fd_sc_hd__o211ai_2 _18236_ (.A1(_02447_),
    .A2(_02440_),
    .B1(_02445_),
    .C1(_02446_),
    .Y(_02449_));
 sky130_fd_sc_hd__a31o_1 _18237_ (.A1(_08194_),
    .A2(_02448_),
    .A3(_02449_),
    .B1(_10335_),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _18238_ (.A0(\rbzero.wall_tracer.trackDistY[2] ),
    .A1(_02450_),
    .S(_02362_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _18239_ (.A(_02451_),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _18240_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_02452_));
 sky130_fd_sc_hd__nor2_1 _18241_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_02453_));
 sky130_fd_sc_hd__o211a_1 _18242_ (.A1(_02452_),
    .A2(_02453_),
    .B1(_02445_),
    .C1(_02449_),
    .X(_02454_));
 sky130_fd_sc_hd__a211oi_2 _18243_ (.A1(_02445_),
    .A2(_02449_),
    .B1(_02452_),
    .C1(_02453_),
    .Y(_02455_));
 sky130_fd_sc_hd__o31a_1 _18244_ (.A1(_01779_),
    .A2(_02454_),
    .A3(_02455_),
    .B1(_02370_),
    .X(_02456_));
 sky130_fd_sc_hd__o2bb2a_1 _18245_ (.A1_N(_01665_),
    .A2_N(_02456_),
    .B1(_02365_),
    .B2(\rbzero.wall_tracer.trackDistY[3] ),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _18246_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .Y(_02457_));
 sky130_fd_sc_hd__or2_1 _18247_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_02458_));
 sky130_fd_sc_hd__o211a_1 _18248_ (.A1(_02452_),
    .A2(_02455_),
    .B1(_02457_),
    .C1(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__a211oi_1 _18249_ (.A1(_02457_),
    .A2(_02458_),
    .B1(_02452_),
    .C1(_02455_),
    .Y(_02460_));
 sky130_fd_sc_hd__o31a_1 _18250_ (.A1(_06164_),
    .A2(_02459_),
    .A3(_02460_),
    .B1(_02370_),
    .X(_02461_));
 sky130_fd_sc_hd__o2bb2a_1 _18251_ (.A1_N(_01778_),
    .A2_N(_02461_),
    .B1(_02363_),
    .B2(\rbzero.wall_tracer.trackDistY[4] ),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _18252_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_02462_));
 sky130_fd_sc_hd__and2_1 _18253_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_02463_));
 sky130_fd_sc_hd__a21oi_1 _18254_ (.A1(\rbzero.wall_tracer.trackDistY[4] ),
    .A2(\rbzero.wall_tracer.stepDistY[4] ),
    .B1(_02459_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor3_1 _18255_ (.A(_02462_),
    .B(_02463_),
    .C(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__o21a_1 _18256_ (.A1(_02462_),
    .A2(_02463_),
    .B1(_02464_),
    .X(_02466_));
 sky130_fd_sc_hd__o31a_1 _18257_ (.A1(_06164_),
    .A2(_02465_),
    .A3(_02466_),
    .B1(_02370_),
    .X(_02467_));
 sky130_fd_sc_hd__o2bb2a_1 _18258_ (.A1_N(_01894_),
    .A2_N(_02467_),
    .B1(_02363_),
    .B2(\rbzero.wall_tracer.trackDistY[5] ),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_1 _18259_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02468_));
 sky130_fd_sc_hd__nand2_1 _18260_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02469_));
 sky130_fd_sc_hd__or2b_1 _18261_ (.A(_02468_),
    .B_N(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__o21ba_1 _18262_ (.A1(_02462_),
    .A2(_02464_),
    .B1_N(_02463_),
    .X(_02471_));
 sky130_fd_sc_hd__nor2_1 _18263_ (.A(_02470_),
    .B(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__a21o_1 _18264_ (.A1(_02470_),
    .A2(_02471_),
    .B1(_06163_),
    .X(_02473_));
 sky130_fd_sc_hd__o21ai_1 _18265_ (.A1(_02472_),
    .A2(_02473_),
    .B1(_02006_),
    .Y(_02474_));
 sky130_fd_sc_hd__mux2_1 _18266_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(_02474_),
    .S(_02362_),
    .X(_02475_));
 sky130_fd_sc_hd__clkbuf_1 _18267_ (.A(_02475_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _18268_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_1 _18269_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02477_));
 sky130_fd_sc_hd__or2b_1 _18270_ (.A(_02476_),
    .B_N(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__o21a_1 _18271_ (.A1(_02468_),
    .A2(_02471_),
    .B1(_02469_),
    .X(_02479_));
 sky130_fd_sc_hd__nor2_1 _18272_ (.A(_02478_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__a21o_1 _18273_ (.A1(_02478_),
    .A2(_02479_),
    .B1(_06163_),
    .X(_02481_));
 sky130_fd_sc_hd__o21ai_1 _18274_ (.A1(_02480_),
    .A2(_02481_),
    .B1(_02111_),
    .Y(_02482_));
 sky130_fd_sc_hd__mux2_1 _18275_ (.A0(\rbzero.wall_tracer.trackDistY[7] ),
    .A1(_02482_),
    .S(_02362_),
    .X(_02483_));
 sky130_fd_sc_hd__clkbuf_1 _18276_ (.A(_02483_),
    .X(_00568_));
 sky130_fd_sc_hd__or2_1 _18277_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .X(_02484_));
 sky130_fd_sc_hd__nand2_1 _18278_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_02485_));
 sky130_fd_sc_hd__nand2_1 _18279_ (.A(_02484_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__o21a_1 _18280_ (.A1(_02476_),
    .A2(_02479_),
    .B1(_02477_),
    .X(_02487_));
 sky130_fd_sc_hd__nor2_1 _18281_ (.A(_02486_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__a21o_1 _18282_ (.A1(_02486_),
    .A2(_02487_),
    .B1(_09905_),
    .X(_02489_));
 sky130_fd_sc_hd__o21a_1 _18283_ (.A1(_02488_),
    .A2(_02489_),
    .B1(_02363_),
    .X(_02490_));
 sky130_fd_sc_hd__o2bb2a_1 _18284_ (.A1_N(_02203_),
    .A2_N(_02490_),
    .B1(_02363_),
    .B2(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_00569_));
 sky130_fd_sc_hd__and2_1 _18285_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_02491_));
 sky130_fd_sc_hd__nor2_1 _18286_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_02492_));
 sky130_fd_sc_hd__nor2_1 _18287_ (.A(_02491_),
    .B(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__nand2_1 _18288_ (.A(_02485_),
    .B(_02487_),
    .Y(_02494_));
 sky130_fd_sc_hd__and2_1 _18289_ (.A(_02484_),
    .B(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__xnor2_1 _18290_ (.A(_02493_),
    .B(_02495_),
    .Y(_02496_));
 sky130_fd_sc_hd__o21a_1 _18291_ (.A1(_08156_),
    .A2(_02496_),
    .B1(_02363_),
    .X(_02497_));
 sky130_fd_sc_hd__o2bb2a_1 _18292_ (.A1_N(_02288_),
    .A2_N(_02497_),
    .B1(_02363_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .X(_00570_));
 sky130_fd_sc_hd__a31o_1 _18293_ (.A1(_02484_),
    .A2(_02493_),
    .A3(_02494_),
    .B1(_02491_),
    .X(_02498_));
 sky130_fd_sc_hd__xor2_1 _18294_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .X(_02499_));
 sky130_fd_sc_hd__xnor2_1 _18295_ (.A(_02498_),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__o21a_1 _18296_ (.A1(_08156_),
    .A2(_02500_),
    .B1(_02363_),
    .X(_02501_));
 sky130_fd_sc_hd__o2bb2a_1 _18297_ (.A1_N(_02355_),
    .A2_N(_02501_),
    .B1(_02363_),
    .B2(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_00571_));
 sky130_fd_sc_hd__clkbuf_8 _18298_ (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .X(_02502_));
 sky130_fd_sc_hd__buf_2 _18299_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02503_));
 sky130_fd_sc_hd__inv_2 _18300_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .Y(_02504_));
 sky130_fd_sc_hd__or4b_4 _18301_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .B(_02504_),
    .C(_04468_),
    .D_N(\rbzero.spi_registers.spi_done ),
    .X(_02505_));
 sky130_fd_sc_hd__nor3b_4 _18302_ (.A(_02503_),
    .B(_02505_),
    .C_N(\rbzero.spi_registers.spi_cmd[0] ),
    .Y(_02506_));
 sky130_fd_sc_hd__clkbuf_4 _18303_ (.A(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _18304_ (.A0(\rbzero.spi_registers.new_texadd[2][0] ),
    .A1(_02502_),
    .S(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__clkbuf_1 _18305_ (.A(_02508_),
    .X(_00572_));
 sky130_fd_sc_hd__buf_4 _18306_ (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _18307_ (.A0(\rbzero.spi_registers.new_texadd[2][1] ),
    .A1(_02509_),
    .S(_02507_),
    .X(_02510_));
 sky130_fd_sc_hd__clkbuf_1 _18308_ (.A(_02510_),
    .X(_00573_));
 sky130_fd_sc_hd__buf_4 _18309_ (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _18310_ (.A0(\rbzero.spi_registers.new_texadd[2][2] ),
    .A1(_02511_),
    .S(_02507_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _18311_ (.A(_02512_),
    .X(_00574_));
 sky130_fd_sc_hd__buf_4 _18312_ (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _18313_ (.A0(\rbzero.spi_registers.new_texadd[2][3] ),
    .A1(_02513_),
    .S(_02507_),
    .X(_02514_));
 sky130_fd_sc_hd__clkbuf_1 _18314_ (.A(_02514_),
    .X(_00575_));
 sky130_fd_sc_hd__buf_4 _18315_ (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _18316_ (.A0(\rbzero.spi_registers.new_texadd[2][4] ),
    .A1(_02515_),
    .S(_02507_),
    .X(_02516_));
 sky130_fd_sc_hd__clkbuf_1 _18317_ (.A(_02516_),
    .X(_00576_));
 sky130_fd_sc_hd__clkbuf_4 _18318_ (.A(\rbzero.spi_registers.spi_buffer[5] ),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _18319_ (.A0(\rbzero.spi_registers.new_texadd[2][5] ),
    .A1(_02517_),
    .S(_02507_),
    .X(_02518_));
 sky130_fd_sc_hd__clkbuf_1 _18320_ (.A(_02518_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _18321_ (.A0(\rbzero.spi_registers.new_texadd[2][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02507_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_1 _18322_ (.A(_02519_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _18323_ (.A0(\rbzero.spi_registers.new_texadd[2][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02507_),
    .X(_02520_));
 sky130_fd_sc_hd__clkbuf_1 _18324_ (.A(_02520_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _18325_ (.A0(\rbzero.spi_registers.new_texadd[2][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02507_),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _18326_ (.A(_02521_),
    .X(_00580_));
 sky130_fd_sc_hd__buf_4 _18327_ (.A(_02506_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _18328_ (.A0(\rbzero.spi_registers.new_texadd[2][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _18329_ (.A(_02523_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _18330_ (.A0(\rbzero.spi_registers.new_texadd[2][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02522_),
    .X(_02524_));
 sky130_fd_sc_hd__clkbuf_1 _18331_ (.A(_02524_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _18332_ (.A0(\rbzero.spi_registers.new_texadd[2][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_02522_),
    .X(_02525_));
 sky130_fd_sc_hd__clkbuf_1 _18333_ (.A(_02525_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _18334_ (.A0(\rbzero.spi_registers.new_texadd[2][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_02522_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_1 _18335_ (.A(_02526_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _18336_ (.A0(\rbzero.spi_registers.new_texadd[2][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_02522_),
    .X(_02527_));
 sky130_fd_sc_hd__clkbuf_1 _18337_ (.A(_02527_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _18338_ (.A0(\rbzero.spi_registers.new_texadd[2][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_02522_),
    .X(_02528_));
 sky130_fd_sc_hd__clkbuf_1 _18339_ (.A(_02528_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _18340_ (.A0(\rbzero.spi_registers.new_texadd[2][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_02522_),
    .X(_02529_));
 sky130_fd_sc_hd__clkbuf_1 _18341_ (.A(_02529_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _18342_ (.A0(\rbzero.spi_registers.new_texadd[2][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_02522_),
    .X(_02530_));
 sky130_fd_sc_hd__clkbuf_1 _18343_ (.A(_02530_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _18344_ (.A0(\rbzero.spi_registers.new_texadd[2][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_02522_),
    .X(_02531_));
 sky130_fd_sc_hd__clkbuf_1 _18345_ (.A(_02531_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _18346_ (.A0(\rbzero.spi_registers.new_texadd[2][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_02522_),
    .X(_02532_));
 sky130_fd_sc_hd__clkbuf_1 _18347_ (.A(_02532_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _18348_ (.A0(\rbzero.spi_registers.new_texadd[2][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_02506_),
    .X(_02533_));
 sky130_fd_sc_hd__clkbuf_1 _18349_ (.A(_02533_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _18350_ (.A0(\rbzero.spi_registers.new_texadd[2][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_02506_),
    .X(_02534_));
 sky130_fd_sc_hd__clkbuf_1 _18351_ (.A(_02534_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _18352_ (.A0(\rbzero.spi_registers.new_texadd[2][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_02506_),
    .X(_02535_));
 sky130_fd_sc_hd__clkbuf_1 _18353_ (.A(_02535_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _18354_ (.A0(\rbzero.spi_registers.new_texadd[2][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_02506_),
    .X(_02536_));
 sky130_fd_sc_hd__clkbuf_1 _18355_ (.A(_02536_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _18356_ (.A0(\rbzero.spi_registers.new_texadd[2][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_02506_),
    .X(_02537_));
 sky130_fd_sc_hd__clkbuf_1 _18357_ (.A(_02537_),
    .X(_00595_));
 sky130_fd_sc_hd__nor2_1 _18358_ (.A(_05153_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2_1 _18359_ (.A(_05153_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02539_));
 sky130_fd_sc_hd__and2b_1 _18360_ (.A_N(_02538_),
    .B(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__or2_1 _18361_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .X(_02541_));
 sky130_fd_sc_hd__nor2_1 _18362_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_1 _18363_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .Y(_02543_));
 sky130_fd_sc_hd__nand2_1 _18364_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_02544_));
 sky130_fd_sc_hd__or2_1 _18365_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_02545_));
 sky130_fd_sc_hd__nand2_1 _18366_ (.A(_02544_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__o21a_1 _18367_ (.A1(_02543_),
    .A2(_02546_),
    .B1(_02544_),
    .X(_02547_));
 sky130_fd_sc_hd__nand2_1 _18368_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02548_));
 sky130_fd_sc_hd__o21ai_1 _18369_ (.A1(_02542_),
    .A2(_02547_),
    .B1(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2_1 _18370_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .Y(_02550_));
 sky130_fd_sc_hd__a21boi_1 _18371_ (.A1(_02541_),
    .A2(_02549_),
    .B1_N(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__xnor2_1 _18372_ (.A(_02540_),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__inv_2 _18373_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _18374_ (.A(_02553_),
    .B(_08128_),
    .Y(_02554_));
 sky130_fd_sc_hd__a221o_1 _18375_ (.A1(\rbzero.wall_tracer.rayAddendX[-5] ),
    .A2(_09822_),
    .B1(_09826_),
    .B2(_02552_),
    .C1(_02554_),
    .X(_00596_));
 sky130_fd_sc_hd__or2_1 _18376_ (.A(_04489_),
    .B(_09819_),
    .X(_02555_));
 sky130_fd_sc_hd__buf_4 _18377_ (.A(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__buf_4 _18378_ (.A(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__nor2_1 _18379_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .Y(_02558_));
 sky130_fd_sc_hd__and2_1 _18380_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_02559_));
 sky130_fd_sc_hd__o21ai_1 _18381_ (.A1(_02538_),
    .A2(_02551_),
    .B1(_02539_),
    .Y(_02560_));
 sky130_fd_sc_hd__or3_1 _18382_ (.A(_02558_),
    .B(_02559_),
    .C(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__o21ai_1 _18383_ (.A1(_02558_),
    .A2(_02559_),
    .B1(_02560_),
    .Y(_02562_));
 sky130_fd_sc_hd__a21oi_1 _18384_ (.A1(_02561_),
    .A2(_02562_),
    .B1(_08201_),
    .Y(_02563_));
 sky130_fd_sc_hd__buf_4 _18385_ (.A(_08200_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _18386_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_02565_));
 sky130_fd_sc_hd__or2_1 _18387_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_02566_));
 sky130_fd_sc_hd__a31o_1 _18388_ (.A1(_02564_),
    .A2(_02565_),
    .A3(_02566_),
    .B1(_09829_),
    .X(_02567_));
 sky130_fd_sc_hd__o22a_1 _18389_ (.A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_02557_),
    .B1(_02563_),
    .B2(_02567_),
    .X(_00597_));
 sky130_fd_sc_hd__nor2_1 _18390_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02568_));
 sky130_fd_sc_hd__and2_1 _18391_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .X(_02569_));
 sky130_fd_sc_hd__or2_1 _18392_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_02570_));
 sky130_fd_sc_hd__a21oi_1 _18393_ (.A1(_02570_),
    .A2(_02560_),
    .B1(_02559_),
    .Y(_02571_));
 sky130_fd_sc_hd__o21ai_1 _18394_ (.A1(_02568_),
    .A2(_02569_),
    .B1(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__o311a_1 _18395_ (.A1(_02568_),
    .A2(_02569_),
    .A3(_02571_),
    .B1(_02572_),
    .C1(_08136_),
    .X(_02573_));
 sky130_fd_sc_hd__or2_1 _18396_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02566_),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_1 _18397_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02566_),
    .Y(_02575_));
 sky130_fd_sc_hd__a31o_1 _18398_ (.A1(_02564_),
    .A2(_02574_),
    .A3(_02575_),
    .B1(_09829_),
    .X(_02576_));
 sky130_fd_sc_hd__o22a_1 _18399_ (.A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A2(_02557_),
    .B1(_02573_),
    .B2(_02576_),
    .X(_00598_));
 sky130_fd_sc_hd__clkbuf_4 _18400_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_02577_));
 sky130_fd_sc_hd__nor2_1 _18401_ (.A(_02577_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_02578_));
 sky130_fd_sc_hd__and2_1 _18402_ (.A(_02577_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02579_));
 sky130_fd_sc_hd__nand2_1 _18403_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02580_));
 sky130_fd_sc_hd__o21ai_1 _18404_ (.A1(_02568_),
    .A2(_02571_),
    .B1(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__or3_1 _18405_ (.A(_02578_),
    .B(_02579_),
    .C(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__o21ai_1 _18406_ (.A1(_02578_),
    .A2(_02579_),
    .B1(_02581_),
    .Y(_02583_));
 sky130_fd_sc_hd__a21oi_1 _18407_ (.A1(_02582_),
    .A2(_02583_),
    .B1(_08201_),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_1 _18408_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_02574_),
    .Y(_02585_));
 sky130_fd_sc_hd__or2_1 _18409_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_02574_),
    .X(_02586_));
 sky130_fd_sc_hd__a31o_1 _18410_ (.A1(_02564_),
    .A2(_02585_),
    .A3(_02586_),
    .B1(_09829_),
    .X(_02587_));
 sky130_fd_sc_hd__o22a_1 _18411_ (.A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A2(_02557_),
    .B1(_02584_),
    .B2(_02587_),
    .X(_00599_));
 sky130_fd_sc_hd__or2_1 _18412_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02588_));
 sky130_fd_sc_hd__nand2_1 _18413_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_02589_));
 sky130_fd_sc_hd__or2_1 _18414_ (.A(_02577_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02590_));
 sky130_fd_sc_hd__a21o_1 _18415_ (.A1(_02590_),
    .A2(_02581_),
    .B1(_02579_),
    .X(_02591_));
 sky130_fd_sc_hd__a21oi_1 _18416_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__a31o_1 _18417_ (.A1(_02588_),
    .A2(_02589_),
    .A3(_02591_),
    .B1(_09828_),
    .X(_02593_));
 sky130_fd_sc_hd__o31a_1 _18418_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(\rbzero.debug_overlay.vplaneX[-7] ),
    .A3(\rbzero.debug_overlay.vplaneX[-8] ),
    .B1(_02553_),
    .X(_02594_));
 sky130_fd_sc_hd__xnor2_1 _18419_ (.A(_05153_),
    .B(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__o2bb2a_1 _18420_ (.A1_N(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A2_N(_09821_),
    .B1(_02595_),
    .B2(_04491_),
    .X(_02596_));
 sky130_fd_sc_hd__o21ai_1 _18421_ (.A1(_02592_),
    .A2(_02593_),
    .B1(_02596_),
    .Y(_00600_));
 sky130_fd_sc_hd__a21bo_1 _18422_ (.A1(_02588_),
    .A2(_02591_),
    .B1_N(_02589_),
    .X(_02597_));
 sky130_fd_sc_hd__clkbuf_4 _18423_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_02598_));
 sky130_fd_sc_hd__nor2_1 _18424_ (.A(_02598_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_02599_));
 sky130_fd_sc_hd__and2_1 _18425_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_02600_));
 sky130_fd_sc_hd__or2_1 _18426_ (.A(_02599_),
    .B(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__xnor2_1 _18427_ (.A(_02597_),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__or2_1 _18428_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_02603_));
 sky130_fd_sc_hd__nand2_1 _18429_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .Y(_02604_));
 sky130_fd_sc_hd__nand2_1 _18430_ (.A(_02603_),
    .B(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__nor2_1 _18431_ (.A(_05153_),
    .B(_02586_),
    .Y(_02606_));
 sky130_fd_sc_hd__a21oi_1 _18432_ (.A1(_05153_),
    .A2(\rbzero.debug_overlay.vplaneX[-9] ),
    .B1(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__xnor2_1 _18433_ (.A(_02605_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__mux2_1 _18434_ (.A0(_02602_),
    .A1(_02608_),
    .S(_08200_),
    .X(_02609_));
 sky130_fd_sc_hd__mux2_1 _18435_ (.A0(\rbzero.wall_tracer.rayAddendX[0] ),
    .A1(_02609_),
    .S(_02556_),
    .X(_02610_));
 sky130_fd_sc_hd__clkbuf_1 _18436_ (.A(_02610_),
    .X(_00601_));
 sky130_fd_sc_hd__buf_4 _18437_ (.A(_09825_),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_1 _18438_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_02612_));
 sky130_fd_sc_hd__or2_1 _18439_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02613_));
 sky130_fd_sc_hd__o21a_1 _18440_ (.A1(_02598_),
    .A2(\rbzero.wall_tracer.rayAddendX[0] ),
    .B1(_02597_),
    .X(_02614_));
 sky130_fd_sc_hd__a211o_1 _18441_ (.A1(_02612_),
    .A2(_02613_),
    .B1(_02614_),
    .C1(_02600_),
    .X(_02615_));
 sky130_fd_sc_hd__o211ai_2 _18442_ (.A1(_02600_),
    .A2(_02614_),
    .B1(_02613_),
    .C1(_02612_),
    .Y(_02616_));
 sky130_fd_sc_hd__clkbuf_4 _18443_ (.A(_08200_),
    .X(_02617_));
 sky130_fd_sc_hd__a21oi_1 _18444_ (.A1(_05153_),
    .A2(\rbzero.debug_overlay.vplaneX[-9] ),
    .B1(_02605_),
    .Y(_02618_));
 sky130_fd_sc_hd__nor2_1 _18445_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_02619_));
 sky130_fd_sc_hd__and2_1 _18446_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_02620_));
 sky130_fd_sc_hd__nor2_1 _18447_ (.A(_02619_),
    .B(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__xnor2_1 _18448_ (.A(_02603_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__o21a_1 _18449_ (.A1(_02606_),
    .A2(_02618_),
    .B1(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__inv_2 _18450_ (.A(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__or3_1 _18451_ (.A(_02606_),
    .B(_02622_),
    .C(_02618_),
    .X(_02625_));
 sky130_fd_sc_hd__a32o_1 _18452_ (.A1(_02617_),
    .A2(_02624_),
    .A3(_02625_),
    .B1(_09822_),
    .B2(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02626_));
 sky130_fd_sc_hd__a31o_1 _18453_ (.A1(_02611_),
    .A2(_02615_),
    .A3(_02616_),
    .B1(_02626_),
    .X(_00602_));
 sky130_fd_sc_hd__buf_2 _18454_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_02627_));
 sky130_fd_sc_hd__buf_2 _18455_ (.A(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__clkbuf_4 _18456_ (.A(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__xnor2_1 _18457_ (.A(_02629_),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_02630_));
 sky130_fd_sc_hd__a21oi_1 _18458_ (.A1(_02612_),
    .A2(_02616_),
    .B1(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__a311oi_1 _18459_ (.A1(_02612_),
    .A2(_02616_),
    .A3(_02630_),
    .B1(_02631_),
    .C1(_08201_),
    .Y(_02632_));
 sky130_fd_sc_hd__xor2_1 _18460_ (.A(_02577_),
    .B(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_02633_));
 sky130_fd_sc_hd__o31ai_1 _18461_ (.A1(_02603_),
    .A2(_02619_),
    .A3(_02620_),
    .B1(_02624_),
    .Y(_02634_));
 sky130_fd_sc_hd__xnor2_1 _18462_ (.A(_02633_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__xnor2_1 _18463_ (.A(_02619_),
    .B(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__a21o_1 _18464_ (.A1(_08201_),
    .A2(_02636_),
    .B1(_09822_),
    .X(_02637_));
 sky130_fd_sc_hd__o22a_1 _18465_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(_02557_),
    .B1(_02632_),
    .B2(_02637_),
    .X(_00603_));
 sky130_fd_sc_hd__and2_1 _18466_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02638_));
 sky130_fd_sc_hd__nor2_1 _18467_ (.A(_02627_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02639_));
 sky130_fd_sc_hd__o21ai_1 _18468_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[1] ),
    .B1(_02627_),
    .Y(_02640_));
 sky130_fd_sc_hd__o21bai_1 _18469_ (.A1(_02627_),
    .A2(\rbzero.wall_tracer.rayAddendX[2] ),
    .B1_N(_02616_),
    .Y(_02641_));
 sky130_fd_sc_hd__o211ai_1 _18470_ (.A1(_02638_),
    .A2(_02639_),
    .B1(_02640_),
    .C1(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__a211o_1 _18471_ (.A1(_02640_),
    .A2(_02641_),
    .B1(_02638_),
    .C1(_02639_),
    .X(_02643_));
 sky130_fd_sc_hd__or2_1 _18472_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05153_),
    .X(_02644_));
 sky130_fd_sc_hd__nand2_1 _18473_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05153_),
    .Y(_02645_));
 sky130_fd_sc_hd__and4bb_1 _18474_ (.A_N(_02577_),
    .B_N(\rbzero.debug_overlay.vplaneX[-6] ),
    .C(_02644_),
    .D(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__a2bb2o_1 _18475_ (.A1_N(_02577_),
    .A2_N(\rbzero.debug_overlay.vplaneX[-6] ),
    .B1(_02644_),
    .B2(_02645_),
    .X(_02647_));
 sky130_fd_sc_hd__and2b_1 _18476_ (.A_N(_02646_),
    .B(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__o21a_1 _18477_ (.A1(_02623_),
    .A2(_02633_),
    .B1(_02619_),
    .X(_02649_));
 sky130_fd_sc_hd__a21o_1 _18478_ (.A1(_02633_),
    .A2(_02634_),
    .B1(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__and2_1 _18479_ (.A(_02648_),
    .B(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__o21ai_1 _18480_ (.A1(_02648_),
    .A2(_02650_),
    .B1(_08200_),
    .Y(_02652_));
 sky130_fd_sc_hd__a2bb2o_1 _18481_ (.A1_N(_02651_),
    .A2_N(_02652_),
    .B1(\rbzero.wall_tracer.rayAddendX[3] ),
    .B2(_09821_),
    .X(_02653_));
 sky130_fd_sc_hd__a31o_1 _18482_ (.A1(_02611_),
    .A2(_02642_),
    .A3(_02643_),
    .B1(_02653_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _18483_ (.A(_02629_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02654_));
 sky130_fd_sc_hd__xor2_1 _18484_ (.A(_02627_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_02655_));
 sky130_fd_sc_hd__a21oi_1 _18485_ (.A1(_02654_),
    .A2(_02643_),
    .B1(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__a31o_1 _18486_ (.A1(_02654_),
    .A2(_02643_),
    .A3(_02655_),
    .B1(_04489_),
    .X(_02657_));
 sky130_fd_sc_hd__xor2_1 _18487_ (.A(_02598_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_02658_));
 sky130_fd_sc_hd__o21ai_1 _18488_ (.A1(_02646_),
    .A2(_02651_),
    .B1(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__or3_1 _18489_ (.A(_02646_),
    .B(_02651_),
    .C(_02658_),
    .X(_02660_));
 sky130_fd_sc_hd__and2_1 _18490_ (.A(_02659_),
    .B(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__xnor2_1 _18491_ (.A(_02644_),
    .B(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__o22a_1 _18492_ (.A1(_02656_),
    .A2(_02657_),
    .B1(_02662_),
    .B2(_04491_),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _18493_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02663_),
    .S(_02556_),
    .X(_02664_));
 sky130_fd_sc_hd__clkbuf_1 _18494_ (.A(_02664_),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _18495_ (.A(_02627_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02665_));
 sky130_fd_sc_hd__or2_1 _18496_ (.A(_02627_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_1 _18497_ (.A(_02665_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__or2b_1 _18498_ (.A(_02643_),
    .B_N(_02655_),
    .X(_02668_));
 sky130_fd_sc_hd__o21ai_1 _18499_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02629_),
    .Y(_02669_));
 sky130_fd_sc_hd__nand3_1 _18500_ (.A(_02667_),
    .B(_02668_),
    .C(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__a21o_1 _18501_ (.A1(_02668_),
    .A2(_02669_),
    .B1(_02667_),
    .X(_02671_));
 sky130_fd_sc_hd__nor2_1 _18502_ (.A(_02627_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .Y(_02672_));
 sky130_fd_sc_hd__and2_1 _18503_ (.A(_02627_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_02673_));
 sky130_fd_sc_hd__o22a_1 _18504_ (.A1(_02598_),
    .A2(\rbzero.debug_overlay.vplaneX[-4] ),
    .B1(_02672_),
    .B2(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__nor4_1 _18505_ (.A(_02598_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .C(_02672_),
    .D(_02673_),
    .Y(_02675_));
 sky130_fd_sc_hd__nor2_1 _18506_ (.A(_02674_),
    .B(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__a2bb2o_1 _18507_ (.A1_N(_02651_),
    .A2_N(_02658_),
    .B1(_02659_),
    .B2(_02644_),
    .X(_02677_));
 sky130_fd_sc_hd__xnor2_1 _18508_ (.A(_02676_),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__a22o_1 _18509_ (.A1(\rbzero.wall_tracer.rayAddendX[5] ),
    .A2(_09821_),
    .B1(_02678_),
    .B2(_02564_),
    .X(_02679_));
 sky130_fd_sc_hd__a31o_1 _18510_ (.A1(_02611_),
    .A2(_02670_),
    .A3(_02671_),
    .B1(_02679_),
    .X(_00606_));
 sky130_fd_sc_hd__xnor2_1 _18511_ (.A(_02628_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_02680_));
 sky130_fd_sc_hd__a21o_1 _18512_ (.A1(_02665_),
    .A2(_02671_),
    .B1(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__nand3_1 _18513_ (.A(_02665_),
    .B(_02671_),
    .C(_02680_),
    .Y(_02682_));
 sky130_fd_sc_hd__or2_1 _18514_ (.A(_02627_),
    .B(_02577_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _18515_ (.A(_02628_),
    .B(_02577_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21o_1 _18516_ (.A1(_02683_),
    .A2(_02684_),
    .B1(_02672_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_1 _18517_ (.A(_02577_),
    .B(_02672_),
    .Y(_02686_));
 sky130_fd_sc_hd__nand2_1 _18518_ (.A(_02685_),
    .B(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__o21bai_1 _18519_ (.A1(_02674_),
    .A2(_02677_),
    .B1_N(_02675_),
    .Y(_02688_));
 sky130_fd_sc_hd__xnor2_1 _18520_ (.A(_02687_),
    .B(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__a22o_1 _18521_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(_09821_),
    .B1(_02689_),
    .B2(_02564_),
    .X(_02690_));
 sky130_fd_sc_hd__a31o_1 _18522_ (.A1(_02611_),
    .A2(_02681_),
    .A3(_02682_),
    .B1(_02690_),
    .X(_00607_));
 sky130_fd_sc_hd__nand2_1 _18523_ (.A(_02628_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_02691_));
 sky130_fd_sc_hd__or2_1 _18524_ (.A(_02628_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02692_));
 sky130_fd_sc_hd__nor3_1 _18525_ (.A(_02667_),
    .B(_02668_),
    .C(_02680_),
    .Y(_02693_));
 sky130_fd_sc_hd__o41a_1 _18526_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .A3(\rbzero.wall_tracer.rayAddendX[4] ),
    .A4(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02628_),
    .X(_02694_));
 sky130_fd_sc_hd__a211o_1 _18527_ (.A1(_02691_),
    .A2(_02692_),
    .B1(_02693_),
    .C1(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__o211ai_2 _18528_ (.A1(_02693_),
    .A2(_02694_),
    .B1(_02691_),
    .C1(_02692_),
    .Y(_02696_));
 sky130_fd_sc_hd__inv_2 _18529_ (.A(_02686_),
    .Y(_02697_));
 sky130_fd_sc_hd__and3_1 _18530_ (.A(_02685_),
    .B(_02686_),
    .C(_02688_),
    .X(_02698_));
 sky130_fd_sc_hd__nor2_1 _18531_ (.A(_02628_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .Y(_02699_));
 sky130_fd_sc_hd__and2_1 _18532_ (.A(_02628_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_02700_));
 sky130_fd_sc_hd__o21ai_1 _18533_ (.A1(_02699_),
    .A2(_02700_),
    .B1(_02683_),
    .Y(_02701_));
 sky130_fd_sc_hd__or3_1 _18534_ (.A(_02683_),
    .B(_02699_),
    .C(_02700_),
    .X(_02702_));
 sky130_fd_sc_hd__o211ai_2 _18535_ (.A1(_02697_),
    .A2(_02698_),
    .B1(_02701_),
    .C1(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__a211o_1 _18536_ (.A1(_02701_),
    .A2(_02702_),
    .B1(_02697_),
    .C1(_02698_),
    .X(_02704_));
 sky130_fd_sc_hd__a32o_1 _18537_ (.A1(_02617_),
    .A2(_02703_),
    .A3(_02704_),
    .B1(_09822_),
    .B2(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02705_));
 sky130_fd_sc_hd__a31o_1 _18538_ (.A1(_02611_),
    .A2(_02695_),
    .A3(_02696_),
    .B1(_02705_),
    .X(_00608_));
 sky130_fd_sc_hd__xnor2_1 _18539_ (.A(_02628_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_02706_));
 sky130_fd_sc_hd__a21oi_1 _18540_ (.A1(_02691_),
    .A2(_02696_),
    .B1(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__a31o_1 _18541_ (.A1(_02691_),
    .A2(_02696_),
    .A3(_02706_),
    .B1(_08200_),
    .X(_02708_));
 sky130_fd_sc_hd__nor2_1 _18542_ (.A(_02707_),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__inv_2 _18543_ (.A(_02598_),
    .Y(_02710_));
 sky130_fd_sc_hd__a21oi_1 _18544_ (.A1(_02598_),
    .A2(\rbzero.debug_overlay.vplaneX[-1] ),
    .B1(_02628_),
    .Y(_02711_));
 sky130_fd_sc_hd__a21oi_1 _18545_ (.A1(_02629_),
    .A2(_02598_),
    .B1(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__a21oi_1 _18546_ (.A1(_02710_),
    .A2(_02699_),
    .B1(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__a21o_1 _18547_ (.A1(_02702_),
    .A2(_02703_),
    .B1(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__nand3_1 _18548_ (.A(_02702_),
    .B(_02703_),
    .C(_02713_),
    .Y(_02715_));
 sky130_fd_sc_hd__a31o_1 _18549_ (.A1(_02564_),
    .A2(_02714_),
    .A3(_02715_),
    .B1(_09829_),
    .X(_02716_));
 sky130_fd_sc_hd__o22a_1 _18550_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(_02557_),
    .B1(_02709_),
    .B2(_02716_),
    .X(_00609_));
 sky130_fd_sc_hd__or2_1 _18551_ (.A(_02629_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_02717_));
 sky130_fd_sc_hd__nand2_1 _18552_ (.A(_02629_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_02718_));
 sky130_fd_sc_hd__nand2_1 _18553_ (.A(_02717_),
    .B(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__o21ai_1 _18554_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[7] ),
    .B1(_02629_),
    .Y(_02720_));
 sky130_fd_sc_hd__o21ai_1 _18555_ (.A1(_02696_),
    .A2(_02706_),
    .B1(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__xnor2_1 _18556_ (.A(_02719_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__inv_2 _18557_ (.A(_02629_),
    .Y(_02723_));
 sky130_fd_sc_hd__a21oi_1 _18558_ (.A1(_02723_),
    .A2(_02710_),
    .B1(_02714_),
    .Y(_02724_));
 sky130_fd_sc_hd__a211o_1 _18559_ (.A1(_02711_),
    .A2(_02714_),
    .B1(_02724_),
    .C1(_08136_),
    .X(_02725_));
 sky130_fd_sc_hd__o221a_1 _18560_ (.A1(\rbzero.wall_tracer.rayAddendX[9] ),
    .A2(_02556_),
    .B1(_09828_),
    .B2(_02722_),
    .C1(_02725_),
    .X(_00610_));
 sky130_fd_sc_hd__a21bo_1 _18561_ (.A1(_02717_),
    .A2(_02721_),
    .B1_N(_02718_),
    .X(_02726_));
 sky130_fd_sc_hd__xnor2_1 _18562_ (.A(_02629_),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_02727_));
 sky130_fd_sc_hd__xnor2_1 _18563_ (.A(_02726_),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__o211a_1 _18564_ (.A1(_02598_),
    .A2(_02714_),
    .B1(_08200_),
    .C1(_02723_),
    .X(_02729_));
 sky130_fd_sc_hd__o22a_1 _18565_ (.A1(_02564_),
    .A2(_02728_),
    .B1(_02729_),
    .B2(_09826_),
    .X(_02730_));
 sky130_fd_sc_hd__a21o_1 _18566_ (.A1(\rbzero.wall_tracer.rayAddendX[10] ),
    .A2(_09823_),
    .B1(_02730_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _18567_ (.A0(\rbzero.debug_overlay.playerY[0] ),
    .A1(_06248_),
    .S(_08193_),
    .X(_02731_));
 sky130_fd_sc_hd__mux2_1 _18568_ (.A0(_02731_),
    .A1(\rbzero.map_rom.d6 ),
    .S(_06346_),
    .X(_02732_));
 sky130_fd_sc_hd__clkbuf_1 _18569_ (.A(_02732_),
    .X(_00612_));
 sky130_fd_sc_hd__or2_1 _18570_ (.A(\rbzero.map_rom.d6 ),
    .B(_06149_),
    .X(_02733_));
 sky130_fd_sc_hd__nor2_1 _18571_ (.A(_06163_),
    .B(_06150_),
    .Y(_02734_));
 sky130_fd_sc_hd__a22o_1 _18572_ (.A1(_04734_),
    .A2(_08155_),
    .B1(_02733_),
    .B2(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__mux2_1 _18573_ (.A0(_02735_),
    .A1(\rbzero.map_rom.c6 ),
    .S(_06346_),
    .X(_02736_));
 sky130_fd_sc_hd__clkbuf_1 _18574_ (.A(_02736_),
    .X(_00613_));
 sky130_fd_sc_hd__or3_1 _18575_ (.A(_06145_),
    .B(_06150_),
    .C(_06152_),
    .X(_02737_));
 sky130_fd_sc_hd__nor2_1 _18576_ (.A(_04736_),
    .B(_08194_),
    .Y(_02738_));
 sky130_fd_sc_hd__a31o_1 _18577_ (.A1(_08194_),
    .A2(_06153_),
    .A3(_02737_),
    .B1(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__mux2_1 _18578_ (.A0(_02739_),
    .A1(_06151_),
    .S(_06346_),
    .X(_02740_));
 sky130_fd_sc_hd__clkbuf_1 _18579_ (.A(_02740_),
    .X(_00614_));
 sky130_fd_sc_hd__nand2_1 _18580_ (.A(_06142_),
    .B(_06155_),
    .Y(_02741_));
 sky130_fd_sc_hd__xnor2_1 _18581_ (.A(_06154_),
    .B(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__mux2_1 _18582_ (.A0(\rbzero.debug_overlay.playerY[3] ),
    .A1(_02742_),
    .S(_08193_),
    .X(_02743_));
 sky130_fd_sc_hd__mux2_1 _18583_ (.A0(_02743_),
    .A1(\rbzero.map_rom.a6 ),
    .S(_06346_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_1 _18584_ (.A(_02744_),
    .X(_00615_));
 sky130_fd_sc_hd__a21oi_1 _18585_ (.A1(_06142_),
    .A2(_06156_),
    .B1(_06140_),
    .Y(_02745_));
 sky130_fd_sc_hd__nand2_1 _18586_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .B(_08155_),
    .Y(_02746_));
 sky130_fd_sc_hd__o31ai_1 _18587_ (.A1(_09905_),
    .A2(_06157_),
    .A3(_02745_),
    .B1(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__mux2_1 _18588_ (.A0(_02747_),
    .A1(\rbzero.map_rom.i_row[4] ),
    .S(_06346_),
    .X(_02748_));
 sky130_fd_sc_hd__clkbuf_1 _18589_ (.A(_02748_),
    .X(_00616_));
 sky130_fd_sc_hd__a21oi_1 _18590_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(_06147_),
    .B1(_06157_),
    .Y(_02749_));
 sky130_fd_sc_hd__xnor2_1 _18591_ (.A(_06139_),
    .B(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__mux2_1 _18592_ (.A0(\rbzero.debug_overlay.playerY[5] ),
    .A1(_02750_),
    .S(_08193_),
    .X(_02751_));
 sky130_fd_sc_hd__mux2_1 _18593_ (.A0(_02751_),
    .A1(\rbzero.wall_tracer.mapY[5] ),
    .S(_06343_),
    .X(_02752_));
 sky130_fd_sc_hd__clkbuf_1 _18594_ (.A(_02752_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _18595_ (.A0(\rbzero.debug_overlay.playerX[0] ),
    .A1(_06244_),
    .S(_08193_),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _18596_ (.A0(_02753_),
    .A1(_06283_),
    .S(_09859_),
    .X(_02754_));
 sky130_fd_sc_hd__clkbuf_1 _18597_ (.A(_02754_),
    .X(_00618_));
 sky130_fd_sc_hd__or2_1 _18598_ (.A(_06283_),
    .B(_09843_),
    .X(_02755_));
 sky130_fd_sc_hd__nor2_1 _18599_ (.A(_04735_),
    .B(_08193_),
    .Y(_02756_));
 sky130_fd_sc_hd__a31o_1 _18600_ (.A1(_08194_),
    .A2(_09844_),
    .A3(_02755_),
    .B1(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__mux2_1 _18601_ (.A0(_02757_),
    .A1(_06262_),
    .S(_09859_),
    .X(_02758_));
 sky130_fd_sc_hd__clkbuf_1 _18602_ (.A(_02758_),
    .X(_00619_));
 sky130_fd_sc_hd__xor2_1 _18603_ (.A(_09845_),
    .B(_09848_),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_1 _18604_ (.A0(\rbzero.debug_overlay.playerX[2] ),
    .A1(_02759_),
    .S(_08193_),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _18605_ (.A0(_02760_),
    .A1(_06239_),
    .S(_09859_),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_1 _18606_ (.A(_02761_),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _18607_ (.A(_09842_),
    .B(_09850_),
    .Y(_02762_));
 sky130_fd_sc_hd__xnor2_1 _18608_ (.A(_09849_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__mux2_1 _18609_ (.A0(\rbzero.debug_overlay.playerX[3] ),
    .A1(_02763_),
    .S(_08193_),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _18610_ (.A0(_02764_),
    .A1(_06259_),
    .S(_09859_),
    .X(_02765_));
 sky130_fd_sc_hd__clkbuf_1 _18611_ (.A(_02765_),
    .X(_00621_));
 sky130_fd_sc_hd__a21oi_2 _18612_ (.A1(_09842_),
    .A2(_09851_),
    .B1(_09841_),
    .Y(_02766_));
 sky130_fd_sc_hd__nand2_1 _18613_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_08155_),
    .Y(_02767_));
 sky130_fd_sc_hd__o31ai_2 _18614_ (.A1(_09905_),
    .A2(_09852_),
    .A3(_02766_),
    .B1(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__mux2_1 _18615_ (.A0(\rbzero.map_rom.i_col[4] ),
    .A1(_02768_),
    .S(_09917_),
    .X(_02769_));
 sky130_fd_sc_hd__clkbuf_1 _18616_ (.A(_02769_),
    .X(_00622_));
 sky130_fd_sc_hd__a21oi_1 _18617_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(_09200_),
    .B1(_09852_),
    .Y(_02770_));
 sky130_fd_sc_hd__xnor2_1 _18618_ (.A(_09840_),
    .B(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__mux2_1 _18619_ (.A0(\rbzero.debug_overlay.playerX[5] ),
    .A1(_02771_),
    .S(_08193_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _18620_ (.A0(\rbzero.wall_tracer.mapX[5] ),
    .A1(_02772_),
    .S(_09882_),
    .X(_02773_));
 sky130_fd_sc_hd__clkbuf_1 _18621_ (.A(_02773_),
    .X(_00623_));
 sky130_fd_sc_hd__nor2_1 _18622_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02774_));
 sky130_fd_sc_hd__and2_1 _18623_ (.A(_05173_),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(_02775_));
 sky130_fd_sc_hd__or2_1 _18624_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .X(_02776_));
 sky130_fd_sc_hd__nor2_1 _18625_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _18626_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_02778_));
 sky130_fd_sc_hd__or2_1 _18627_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_02779_));
 sky130_fd_sc_hd__nand4_1 _18628_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .C(_02778_),
    .D(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__and2_1 _18629_ (.A(_02778_),
    .B(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__nand2_1 _18630_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02782_));
 sky130_fd_sc_hd__o21ai_1 _18631_ (.A1(_02777_),
    .A2(_02781_),
    .B1(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand2_1 _18632_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .Y(_02784_));
 sky130_fd_sc_hd__a21boi_1 _18633_ (.A1(_02776_),
    .A2(_02783_),
    .B1_N(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__o21ai_1 _18634_ (.A1(_02774_),
    .A2(_02775_),
    .B1(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__or3_1 _18635_ (.A(_02774_),
    .B(_02775_),
    .C(_02785_),
    .X(_02787_));
 sky130_fd_sc_hd__a22o_1 _18636_ (.A1(_05172_),
    .A2(_02617_),
    .B1(_09822_),
    .B2(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(_02788_));
 sky130_fd_sc_hd__a31o_1 _18637_ (.A1(_02611_),
    .A2(_02786_),
    .A3(_02787_),
    .B1(_02788_),
    .X(_00624_));
 sky130_fd_sc_hd__nor2_1 _18638_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .Y(_02789_));
 sky130_fd_sc_hd__and2_1 _18639_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02790_));
 sky130_fd_sc_hd__nand2_1 _18640_ (.A(_05173_),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02791_));
 sky130_fd_sc_hd__o21ai_1 _18641_ (.A1(_02774_),
    .A2(_02785_),
    .B1(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__or3_1 _18642_ (.A(_02789_),
    .B(_02790_),
    .C(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__o21ai_1 _18643_ (.A1(_02789_),
    .A2(_02790_),
    .B1(_02792_),
    .Y(_02794_));
 sky130_fd_sc_hd__a21oi_1 _18644_ (.A1(_02793_),
    .A2(_02794_),
    .B1(_08201_),
    .Y(_02795_));
 sky130_fd_sc_hd__nand2_1 _18645_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_05172_),
    .Y(_02796_));
 sky130_fd_sc_hd__or2_1 _18646_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_05172_),
    .X(_02797_));
 sky130_fd_sc_hd__a31o_1 _18647_ (.A1(_02617_),
    .A2(_02796_),
    .A3(_02797_),
    .B1(_09829_),
    .X(_02798_));
 sky130_fd_sc_hd__o22a_1 _18648_ (.A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_02557_),
    .B1(_02795_),
    .B2(_02798_),
    .X(_00625_));
 sky130_fd_sc_hd__nor2_1 _18649_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02799_));
 sky130_fd_sc_hd__and2_1 _18650_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .X(_02800_));
 sky130_fd_sc_hd__or2_1 _18651_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02801_));
 sky130_fd_sc_hd__a21oi_1 _18652_ (.A1(_02801_),
    .A2(_02792_),
    .B1(_02790_),
    .Y(_02802_));
 sky130_fd_sc_hd__o21ai_1 _18653_ (.A1(_02799_),
    .A2(_02800_),
    .B1(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__o311a_1 _18654_ (.A1(_02799_),
    .A2(_02800_),
    .A3(_02802_),
    .B1(_02803_),
    .C1(_08136_),
    .X(_02804_));
 sky130_fd_sc_hd__or2_1 _18655_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02797_),
    .X(_02805_));
 sky130_fd_sc_hd__nand2_1 _18656_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02797_),
    .Y(_02806_));
 sky130_fd_sc_hd__a31o_1 _18657_ (.A1(_02617_),
    .A2(_02805_),
    .A3(_02806_),
    .B1(_09829_),
    .X(_02807_));
 sky130_fd_sc_hd__o22a_1 _18658_ (.A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A2(_02557_),
    .B1(_02804_),
    .B2(_02807_),
    .X(_00626_));
 sky130_fd_sc_hd__nor2_1 _18659_ (.A(_05177_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_02808_));
 sky130_fd_sc_hd__and2_1 _18660_ (.A(_05177_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_02809_));
 sky130_fd_sc_hd__nand2_1 _18661_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02810_));
 sky130_fd_sc_hd__o21ai_1 _18662_ (.A1(_02799_),
    .A2(_02802_),
    .B1(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__or3_1 _18663_ (.A(_02808_),
    .B(_02809_),
    .C(_02811_),
    .X(_02812_));
 sky130_fd_sc_hd__o21ai_1 _18664_ (.A1(_02808_),
    .A2(_02809_),
    .B1(_02811_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21oi_1 _18665_ (.A1(_02812_),
    .A2(_02813_),
    .B1(_08201_),
    .Y(_02814_));
 sky130_fd_sc_hd__nand2_1 _18666_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_02805_),
    .Y(_02815_));
 sky130_fd_sc_hd__or2_1 _18667_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_02805_),
    .X(_02816_));
 sky130_fd_sc_hd__a31o_1 _18668_ (.A1(_02617_),
    .A2(_02815_),
    .A3(_02816_),
    .B1(_09821_),
    .X(_02817_));
 sky130_fd_sc_hd__o22a_1 _18669_ (.A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A2(_02557_),
    .B1(_02814_),
    .B2(_02817_),
    .X(_00627_));
 sky130_fd_sc_hd__or2_1 _18670_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02818_));
 sky130_fd_sc_hd__nand2_1 _18671_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_02819_));
 sky130_fd_sc_hd__or2_1 _18672_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_02820_));
 sky130_fd_sc_hd__a21o_1 _18673_ (.A1(_02820_),
    .A2(_02811_),
    .B1(_02809_),
    .X(_02821_));
 sky130_fd_sc_hd__a21oi_1 _18674_ (.A1(_02818_),
    .A2(_02819_),
    .B1(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__a31o_1 _18675_ (.A1(_02818_),
    .A2(_02819_),
    .A3(_02821_),
    .B1(_09828_),
    .X(_02823_));
 sky130_fd_sc_hd__inv_2 _18676_ (.A(_05172_),
    .Y(_02824_));
 sky130_fd_sc_hd__o31a_1 _18677_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(\rbzero.debug_overlay.vplaneY[-7] ),
    .A3(\rbzero.debug_overlay.vplaneY[-8] ),
    .B1(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__xnor2_1 _18678_ (.A(_05173_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__o2bb2a_1 _18679_ (.A1_N(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A2_N(_09821_),
    .B1(_02826_),
    .B2(_04491_),
    .X(_02827_));
 sky130_fd_sc_hd__o21ai_1 _18680_ (.A1(_02822_),
    .A2(_02823_),
    .B1(_02827_),
    .Y(_00628_));
 sky130_fd_sc_hd__a21bo_1 _18681_ (.A1(_02818_),
    .A2(_02821_),
    .B1_N(_02819_),
    .X(_02828_));
 sky130_fd_sc_hd__clkbuf_4 _18682_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_02829_));
 sky130_fd_sc_hd__nor2_1 _18683_ (.A(_02829_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_02830_));
 sky130_fd_sc_hd__and2_1 _18684_ (.A(_02829_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_02831_));
 sky130_fd_sc_hd__or2_1 _18685_ (.A(_02830_),
    .B(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__xnor2_1 _18686_ (.A(_02828_),
    .B(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__or2_1 _18687_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_02834_));
 sky130_fd_sc_hd__nand2_1 _18688_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_1 _18689_ (.A(_02834_),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__nor2_1 _18690_ (.A(_05173_),
    .B(_02816_),
    .Y(_02837_));
 sky130_fd_sc_hd__a21oi_1 _18691_ (.A1(_05173_),
    .A2(_05172_),
    .B1(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__xnor2_1 _18692_ (.A(_02836_),
    .B(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__mux2_1 _18693_ (.A0(_02833_),
    .A1(_02839_),
    .S(_08200_),
    .X(_02840_));
 sky130_fd_sc_hd__mux2_1 _18694_ (.A0(\rbzero.wall_tracer.rayAddendY[0] ),
    .A1(_02840_),
    .S(_02556_),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _18695_ (.A(_02841_),
    .X(_00629_));
 sky130_fd_sc_hd__nand2_1 _18696_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_02842_));
 sky130_fd_sc_hd__or2_1 _18697_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_02843_));
 sky130_fd_sc_hd__o21a_1 _18698_ (.A1(_02829_),
    .A2(\rbzero.wall_tracer.rayAddendY[0] ),
    .B1(_02828_),
    .X(_02844_));
 sky130_fd_sc_hd__a211o_1 _18699_ (.A1(_02842_),
    .A2(_02843_),
    .B1(_02844_),
    .C1(_02831_),
    .X(_02845_));
 sky130_fd_sc_hd__o211ai_2 _18700_ (.A1(_02831_),
    .A2(_02844_),
    .B1(_02843_),
    .C1(_02842_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21oi_1 _18701_ (.A1(_05173_),
    .A2(_05172_),
    .B1(_02836_),
    .Y(_02847_));
 sky130_fd_sc_hd__nor2_1 _18702_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_02848_));
 sky130_fd_sc_hd__and2_1 _18703_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(_02849_));
 sky130_fd_sc_hd__nor2_1 _18704_ (.A(_02848_),
    .B(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__xnor2_1 _18705_ (.A(_02834_),
    .B(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__o21a_1 _18706_ (.A1(_02837_),
    .A2(_02847_),
    .B1(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__inv_2 _18707_ (.A(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__or3_1 _18708_ (.A(_02837_),
    .B(_02851_),
    .C(_02847_),
    .X(_02854_));
 sky130_fd_sc_hd__a32o_1 _18709_ (.A1(_02617_),
    .A2(_02853_),
    .A3(_02854_),
    .B1(_09822_),
    .B2(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_02855_));
 sky130_fd_sc_hd__a31o_1 _18710_ (.A1(_09826_),
    .A2(_02845_),
    .A3(_02846_),
    .B1(_02855_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_2 _18711_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_02856_));
 sky130_fd_sc_hd__buf_2 _18712_ (.A(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__buf_4 _18713_ (.A(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__xnor2_1 _18714_ (.A(_02858_),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_02859_));
 sky130_fd_sc_hd__a21oi_1 _18715_ (.A1(_02842_),
    .A2(_02846_),
    .B1(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__a311oi_1 _18716_ (.A1(_02842_),
    .A2(_02846_),
    .A3(_02859_),
    .B1(_02860_),
    .C1(_08201_),
    .Y(_02861_));
 sky130_fd_sc_hd__xor2_1 _18717_ (.A(_05177_),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_02862_));
 sky130_fd_sc_hd__o31ai_1 _18718_ (.A1(_02834_),
    .A2(_02848_),
    .A3(_02849_),
    .B1(_02853_),
    .Y(_02863_));
 sky130_fd_sc_hd__xnor2_1 _18719_ (.A(_02862_),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__xnor2_1 _18720_ (.A(_02848_),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__a21o_1 _18721_ (.A1(_02564_),
    .A2(_02865_),
    .B1(_09822_),
    .X(_02866_));
 sky130_fd_sc_hd__o22a_1 _18722_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(_02557_),
    .B1(_02861_),
    .B2(_02866_),
    .X(_00631_));
 sky130_fd_sc_hd__o21ai_1 _18723_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(_02856_),
    .Y(_02867_));
 sky130_fd_sc_hd__o21bai_1 _18724_ (.A1(_02856_),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1_N(_02846_),
    .Y(_02868_));
 sky130_fd_sc_hd__and2_1 _18725_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02869_));
 sky130_fd_sc_hd__nor2_1 _18726_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02870_));
 sky130_fd_sc_hd__a211o_1 _18727_ (.A1(_02867_),
    .A2(_02868_),
    .B1(_02869_),
    .C1(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__o211ai_1 _18728_ (.A1(_02869_),
    .A2(_02870_),
    .B1(_02867_),
    .C1(_02868_),
    .Y(_02872_));
 sky130_fd_sc_hd__nand2_1 _18729_ (.A(_02862_),
    .B(_02863_),
    .Y(_02873_));
 sky130_fd_sc_hd__o21ai_1 _18730_ (.A1(_02852_),
    .A2(_02862_),
    .B1(_02848_),
    .Y(_02874_));
 sky130_fd_sc_hd__or2_1 _18731_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_05173_),
    .X(_02875_));
 sky130_fd_sc_hd__nand2_1 _18732_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_05173_),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _18733_ (.A(_02875_),
    .B(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__or3_1 _18734_ (.A(_05177_),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .C(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__o21ai_1 _18735_ (.A1(_05177_),
    .A2(\rbzero.debug_overlay.vplaneY[-6] ),
    .B1(_02877_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_1 _18736_ (.A(_02878_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__a21o_1 _18737_ (.A1(_02873_),
    .A2(_02874_),
    .B1(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__nand3_1 _18738_ (.A(_02873_),
    .B(_02880_),
    .C(_02874_),
    .Y(_02882_));
 sky130_fd_sc_hd__a32o_1 _18739_ (.A1(_02617_),
    .A2(_02881_),
    .A3(_02882_),
    .B1(_09822_),
    .B2(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02883_));
 sky130_fd_sc_hd__a31o_1 _18740_ (.A1(_09826_),
    .A2(_02871_),
    .A3(_02872_),
    .B1(_02883_),
    .X(_00632_));
 sky130_fd_sc_hd__nand2_1 _18741_ (.A(_02858_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02884_));
 sky130_fd_sc_hd__xor2_1 _18742_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_02885_));
 sky130_fd_sc_hd__a21oi_1 _18743_ (.A1(_02884_),
    .A2(_02871_),
    .B1(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__a31o_1 _18744_ (.A1(_02884_),
    .A2(_02871_),
    .A3(_02885_),
    .B1(_04489_),
    .X(_02887_));
 sky130_fd_sc_hd__or2_1 _18745_ (.A(_02829_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_02888_));
 sky130_fd_sc_hd__nand2_1 _18746_ (.A(_02829_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .Y(_02889_));
 sky130_fd_sc_hd__nand2_1 _18747_ (.A(_02888_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__a21o_1 _18748_ (.A1(_02878_),
    .A2(_02881_),
    .B1(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__nand3_1 _18749_ (.A(_02878_),
    .B(_02881_),
    .C(_02890_),
    .Y(_02892_));
 sky130_fd_sc_hd__and2_1 _18750_ (.A(_02891_),
    .B(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__xnor2_1 _18751_ (.A(_02875_),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__o22a_1 _18752_ (.A1(_02886_),
    .A2(_02887_),
    .B1(_02894_),
    .B2(_04491_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _18753_ (.A0(\rbzero.wall_tracer.rayAddendY[4] ),
    .A1(_02895_),
    .S(_02556_),
    .X(_02896_));
 sky130_fd_sc_hd__clkbuf_1 _18754_ (.A(_02896_),
    .X(_00633_));
 sky130_fd_sc_hd__nand2_1 _18755_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_02897_));
 sky130_fd_sc_hd__or2_1 _18756_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_02898_));
 sky130_fd_sc_hd__nand2_1 _18757_ (.A(_02897_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__or2b_1 _18758_ (.A(_02871_),
    .B_N(_02885_),
    .X(_02900_));
 sky130_fd_sc_hd__o21ai_1 _18759_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02857_),
    .Y(_02901_));
 sky130_fd_sc_hd__nand3_1 _18760_ (.A(_02899_),
    .B(_02900_),
    .C(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__a21o_1 _18761_ (.A1(_02900_),
    .A2(_02901_),
    .B1(_02899_),
    .X(_02903_));
 sky130_fd_sc_hd__nor2_1 _18762_ (.A(_02857_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .Y(_02904_));
 sky130_fd_sc_hd__and2_1 _18763_ (.A(_02857_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_02905_));
 sky130_fd_sc_hd__o21a_1 _18764_ (.A1(_02904_),
    .A2(_02905_),
    .B1(_02888_),
    .X(_02906_));
 sky130_fd_sc_hd__nor3_1 _18765_ (.A(_02888_),
    .B(_02904_),
    .C(_02905_),
    .Y(_02907_));
 sky130_fd_sc_hd__nor2_1 _18766_ (.A(_02906_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__a22o_1 _18767_ (.A1(_02881_),
    .A2(_02890_),
    .B1(_02891_),
    .B2(_02875_),
    .X(_02909_));
 sky130_fd_sc_hd__xnor2_1 _18768_ (.A(_02908_),
    .B(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__a22o_1 _18769_ (.A1(\rbzero.wall_tracer.rayAddendY[5] ),
    .A2(_09821_),
    .B1(_02910_),
    .B2(_02564_),
    .X(_02911_));
 sky130_fd_sc_hd__a31o_1 _18770_ (.A1(_09826_),
    .A2(_02902_),
    .A3(_02903_),
    .B1(_02911_),
    .X(_00634_));
 sky130_fd_sc_hd__xnor2_1 _18771_ (.A(_02856_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_02912_));
 sky130_fd_sc_hd__a21oi_1 _18772_ (.A1(_02897_),
    .A2(_02903_),
    .B1(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__a31o_1 _18773_ (.A1(_02897_),
    .A2(_02903_),
    .A3(_02912_),
    .B1(_04489_),
    .X(_02914_));
 sky130_fd_sc_hd__or2_1 _18774_ (.A(_02857_),
    .B(_05177_),
    .X(_02915_));
 sky130_fd_sc_hd__nand2_1 _18775_ (.A(_02857_),
    .B(_05177_),
    .Y(_02916_));
 sky130_fd_sc_hd__a21o_1 _18776_ (.A1(_02915_),
    .A2(_02916_),
    .B1(_02904_),
    .X(_02917_));
 sky130_fd_sc_hd__nand2_1 _18777_ (.A(_05177_),
    .B(_02904_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand2_1 _18778_ (.A(_02917_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__o21bai_1 _18779_ (.A1(_02906_),
    .A2(_02909_),
    .B1_N(_02907_),
    .Y(_02920_));
 sky130_fd_sc_hd__xnor2_1 _18780_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__a2bb2o_1 _18781_ (.A1_N(_02913_),
    .A2_N(_02914_),
    .B1(_02921_),
    .B2(_08200_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _18782_ (.A0(\rbzero.wall_tracer.rayAddendY[6] ),
    .A1(_02922_),
    .S(_02556_),
    .X(_02923_));
 sky130_fd_sc_hd__clkbuf_1 _18783_ (.A(_02923_),
    .X(_00635_));
 sky130_fd_sc_hd__and2_1 _18784_ (.A(_02857_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_02924_));
 sky130_fd_sc_hd__nor2_1 _18785_ (.A(_02857_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_02925_));
 sky130_fd_sc_hd__inv_2 _18786_ (.A(_02856_),
    .Y(_02926_));
 sky130_fd_sc_hd__inv_2 _18787_ (.A(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_02927_));
 sky130_fd_sc_hd__or3_1 _18788_ (.A(_02899_),
    .B(_02900_),
    .C(_02912_),
    .X(_02928_));
 sky130_fd_sc_hd__o2111a_1 _18789_ (.A1(_02926_),
    .A2(_02927_),
    .B1(_02897_),
    .C1(_02901_),
    .D1(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__o21ai_1 _18790_ (.A1(_02924_),
    .A2(_02925_),
    .B1(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__or3_1 _18791_ (.A(_02924_),
    .B(_02925_),
    .C(_02929_),
    .X(_02931_));
 sky130_fd_sc_hd__inv_2 _18792_ (.A(_02918_),
    .Y(_02932_));
 sky130_fd_sc_hd__and3_1 _18793_ (.A(_02917_),
    .B(_02918_),
    .C(_02920_),
    .X(_02933_));
 sky130_fd_sc_hd__nor2_1 _18794_ (.A(_02857_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .Y(_02934_));
 sky130_fd_sc_hd__and2_1 _18795_ (.A(_02857_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_02935_));
 sky130_fd_sc_hd__o21ai_1 _18796_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02915_),
    .Y(_02936_));
 sky130_fd_sc_hd__or3_1 _18797_ (.A(_02915_),
    .B(_02934_),
    .C(_02935_),
    .X(_02937_));
 sky130_fd_sc_hd__o211ai_2 _18798_ (.A1(_02932_),
    .A2(_02933_),
    .B1(_02936_),
    .C1(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__a211o_1 _18799_ (.A1(_02936_),
    .A2(_02937_),
    .B1(_02932_),
    .C1(_02933_),
    .X(_02939_));
 sky130_fd_sc_hd__a32o_1 _18800_ (.A1(_02617_),
    .A2(_02938_),
    .A3(_02939_),
    .B1(_09822_),
    .B2(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_02940_));
 sky130_fd_sc_hd__a31o_1 _18801_ (.A1(_09826_),
    .A2(_02930_),
    .A3(_02931_),
    .B1(_02940_),
    .X(_00636_));
 sky130_fd_sc_hd__xnor2_1 _18802_ (.A(_02858_),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_02941_));
 sky130_fd_sc_hd__and2b_1 _18803_ (.A_N(_02924_),
    .B(_02931_),
    .X(_02942_));
 sky130_fd_sc_hd__o21ai_1 _18804_ (.A1(_02941_),
    .A2(_02942_),
    .B1(_04491_),
    .Y(_02943_));
 sky130_fd_sc_hd__a21oi_1 _18805_ (.A1(_02941_),
    .A2(_02942_),
    .B1(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__inv_2 _18806_ (.A(_02829_),
    .Y(_02945_));
 sky130_fd_sc_hd__a21oi_1 _18807_ (.A1(_02829_),
    .A2(\rbzero.debug_overlay.vplaneY[-1] ),
    .B1(_02858_),
    .Y(_02946_));
 sky130_fd_sc_hd__a21oi_1 _18808_ (.A1(_02858_),
    .A2(_02829_),
    .B1(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__a21oi_1 _18809_ (.A1(_02945_),
    .A2(_02934_),
    .B1(_02947_),
    .Y(_02948_));
 sky130_fd_sc_hd__a21o_1 _18810_ (.A1(_02937_),
    .A2(_02938_),
    .B1(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__nand3_1 _18811_ (.A(_02937_),
    .B(_02938_),
    .C(_02948_),
    .Y(_02950_));
 sky130_fd_sc_hd__a31o_1 _18812_ (.A1(_02617_),
    .A2(_02949_),
    .A3(_02950_),
    .B1(_09821_),
    .X(_02951_));
 sky130_fd_sc_hd__o22a_1 _18813_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(_02557_),
    .B1(_02944_),
    .B2(_02951_),
    .X(_00637_));
 sky130_fd_sc_hd__or2_1 _18814_ (.A(_02858_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_02952_));
 sky130_fd_sc_hd__nand2_1 _18815_ (.A(_02858_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_02953_));
 sky130_fd_sc_hd__nand2_1 _18816_ (.A(_02952_),
    .B(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__nor2_1 _18817_ (.A(_02931_),
    .B(_02941_),
    .Y(_02955_));
 sky130_fd_sc_hd__a211o_1 _18818_ (.A1(_02858_),
    .A2(\rbzero.wall_tracer.rayAddendY[8] ),
    .B1(_02924_),
    .C1(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__xnor2_1 _18819_ (.A(_02954_),
    .B(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__a21oi_1 _18820_ (.A1(_02926_),
    .A2(_02945_),
    .B1(_02949_),
    .Y(_02958_));
 sky130_fd_sc_hd__a211o_1 _18821_ (.A1(_02946_),
    .A2(_02949_),
    .B1(_02958_),
    .C1(_08136_),
    .X(_02959_));
 sky130_fd_sc_hd__o221a_1 _18822_ (.A1(\rbzero.wall_tracer.rayAddendY[9] ),
    .A2(_02556_),
    .B1(_09828_),
    .B2(_02957_),
    .C1(_02959_),
    .X(_00638_));
 sky130_fd_sc_hd__a21bo_1 _18823_ (.A1(_02952_),
    .A2(_02956_),
    .B1_N(_02953_),
    .X(_02960_));
 sky130_fd_sc_hd__xnor2_1 _18824_ (.A(_02858_),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_02961_));
 sky130_fd_sc_hd__xnor2_1 _18825_ (.A(_02960_),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__o211a_1 _18826_ (.A1(_02829_),
    .A2(_02949_),
    .B1(_08200_),
    .C1(_02926_),
    .X(_02963_));
 sky130_fd_sc_hd__o22a_1 _18827_ (.A1(_02564_),
    .A2(_02962_),
    .B1(_02963_),
    .B2(_09826_),
    .X(_02964_));
 sky130_fd_sc_hd__a21o_1 _18828_ (.A1(\rbzero.wall_tracer.rayAddendY[10] ),
    .A2(_09823_),
    .B1(_02964_),
    .X(_00639_));
 sky130_fd_sc_hd__and2b_1 _18829_ (.A_N(\rbzero.spi_registers.sclk_buffer[2] ),
    .B(\rbzero.spi_registers.sclk_buffer[1] ),
    .X(_02965_));
 sky130_fd_sc_hd__buf_2 _18830_ (.A(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__or2_2 _18831_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02503_),
    .X(_02967_));
 sky130_fd_sc_hd__a21oi_1 _18832_ (.A1(\rbzero.spi_registers.spi_cmd[2] ),
    .A2(_02967_),
    .B1(\rbzero.spi_registers.spi_cmd[3] ),
    .Y(_02968_));
 sky130_fd_sc_hd__and2_1 _18833_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .B(_02504_),
    .X(_02969_));
 sky130_fd_sc_hd__nand2_1 _18834_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(\rbzero.spi_registers.spi_cmd[1] ),
    .Y(_02970_));
 sky130_fd_sc_hd__and3b_1 _18835_ (.A_N(\rbzero.spi_registers.spi_cmd[2] ),
    .B(\rbzero.spi_registers.spi_cmd[3] ),
    .C(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__a21oi_1 _18836_ (.A1(_02503_),
    .A2(_02969_),
    .B1(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__or2b_1 _18837_ (.A(_02968_),
    .B_N(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__or3_1 _18838_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .C(\rbzero.spi_registers.spi_cmd[3] ),
    .X(_02974_));
 sky130_fd_sc_hd__o21a_1 _18839_ (.A1(\rbzero.spi_registers.spi_cmd[2] ),
    .A2(\rbzero.spi_registers.spi_cmd[3] ),
    .B1(\rbzero.spi_registers.spi_counter[2] ),
    .X(_02975_));
 sky130_fd_sc_hd__a21oi_1 _18840_ (.A1(_02970_),
    .A2(_02968_),
    .B1(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__and4bb_1 _18841_ (.A_N(\rbzero.spi_registers.spi_counter[2] ),
    .B_N(\rbzero.spi_registers.spi_counter[1] ),
    .C(_02970_),
    .D(_02968_),
    .X(_02977_));
 sky130_fd_sc_hd__a31o_1 _18842_ (.A1(\rbzero.spi_registers.spi_counter[1] ),
    .A2(_02974_),
    .A3(_02976_),
    .B1(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__or4b_1 _18843_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .C(_02973_),
    .D_N(\rbzero.spi_registers.spi_counter[2] ),
    .X(_02979_));
 sky130_fd_sc_hd__inv_2 _18844_ (.A(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__a31o_1 _18845_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02973_),
    .A3(_02978_),
    .B1(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__or2_1 _18846_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02972_),
    .X(_02982_));
 sky130_fd_sc_hd__or2_1 _18847_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(\rbzero.spi_registers.spi_counter[5] ),
    .X(_02983_));
 sky130_fd_sc_hd__a21oi_1 _18848_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_02972_),
    .B1(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__and2_1 _18849_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02503_),
    .X(_02985_));
 sky130_fd_sc_hd__a211o_1 _18850_ (.A1(_02985_),
    .A2(_02969_),
    .B1(_02968_),
    .C1(_02971_),
    .X(_02986_));
 sky130_fd_sc_hd__xnor2_1 _18851_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__and4_1 _18852_ (.A(_02981_),
    .B(_02982_),
    .C(_02984_),
    .D(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__nor2_2 _18853_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_04468_),
    .Y(_02989_));
 sky130_fd_sc_hd__a21bo_1 _18854_ (.A1(_02966_),
    .A2(_02988_),
    .B1_N(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__xnor2_1 _18855_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .B(_02966_),
    .Y(_02991_));
 sky130_fd_sc_hd__nor2_1 _18856_ (.A(_02990_),
    .B(_02991_),
    .Y(_00640_));
 sky130_fd_sc_hd__a21oi_1 _18857_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02966_),
    .B1(\rbzero.spi_registers.spi_counter[1] ),
    .Y(_02992_));
 sky130_fd_sc_hd__and3_1 _18858_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .C(_02966_),
    .X(_02993_));
 sky130_fd_sc_hd__nor3_1 _18859_ (.A(_02990_),
    .B(_02992_),
    .C(_02993_),
    .Y(_00641_));
 sky130_fd_sc_hd__xnor2_1 _18860_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__nor2_1 _18861_ (.A(_02990_),
    .B(_02994_),
    .Y(_00642_));
 sky130_fd_sc_hd__and4_1 _18862_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(\rbzero.spi_registers.spi_counter[2] ),
    .C(\rbzero.spi_registers.spi_counter[1] ),
    .D(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02995_));
 sky130_fd_sc_hd__a21oi_1 _18863_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(_02993_),
    .B1(\rbzero.spi_registers.spi_counter[3] ),
    .Y(_02996_));
 sky130_fd_sc_hd__a211oi_1 _18864_ (.A1(_02966_),
    .A2(_02995_),
    .B1(_02996_),
    .C1(_02990_),
    .Y(_00643_));
 sky130_fd_sc_hd__and3_1 _18865_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02966_),
    .C(_02995_),
    .X(_02997_));
 sky130_fd_sc_hd__a21oi_1 _18866_ (.A1(_02966_),
    .A2(_02995_),
    .B1(\rbzero.spi_registers.spi_counter[4] ),
    .Y(_02998_));
 sky130_fd_sc_hd__nor3_1 _18867_ (.A(_02990_),
    .B(_02997_),
    .C(_02998_),
    .Y(_00644_));
 sky130_fd_sc_hd__and2_1 _18868_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(_02997_),
    .X(_02999_));
 sky130_fd_sc_hd__o21ai_1 _18869_ (.A1(\rbzero.spi_registers.spi_counter[5] ),
    .A2(_02997_),
    .B1(_02989_),
    .Y(_03000_));
 sky130_fd_sc_hd__nor2_1 _18870_ (.A(_02999_),
    .B(_03000_),
    .Y(_00645_));
 sky130_fd_sc_hd__or2_1 _18871_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(_02999_),
    .X(_03001_));
 sky130_fd_sc_hd__nand2_1 _18872_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(_02999_),
    .Y(_03002_));
 sky130_fd_sc_hd__and3_1 _18873_ (.A(_02989_),
    .B(_03001_),
    .C(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_1 _18874_ (.A(_03003_),
    .X(_00646_));
 sky130_fd_sc_hd__nand2_1 _18875_ (.A(\rbzero.pov.spi_done ),
    .B(_04112_),
    .Y(_03004_));
 sky130_fd_sc_hd__buf_4 _18876_ (.A(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_4 _18877_ (.A(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _18878_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.ready_buffer[0] ),
    .S(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _18879_ (.A(_03007_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18880_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.ready_buffer[1] ),
    .S(_03006_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _18881_ (.A(_03008_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _18882_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.ready_buffer[2] ),
    .S(_03006_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _18883_ (.A(_03009_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18884_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.ready_buffer[3] ),
    .S(_03006_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_1 _18885_ (.A(_03010_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _18886_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.ready_buffer[4] ),
    .S(_03006_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_1 _18887_ (.A(_03011_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _18888_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.ready_buffer[5] ),
    .S(_03006_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _18889_ (.A(_03012_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _18890_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.ready_buffer[6] ),
    .S(_03006_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _18891_ (.A(_03013_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18892_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.ready_buffer[7] ),
    .S(_03006_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_1 _18893_ (.A(_03014_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _18894_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.ready_buffer[8] ),
    .S(_03006_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_1 _18895_ (.A(_03015_),
    .X(_00655_));
 sky130_fd_sc_hd__clkbuf_4 _18896_ (.A(_03005_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _18897_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.ready_buffer[9] ),
    .S(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_1 _18898_ (.A(_03017_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _18899_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.ready_buffer[10] ),
    .S(_03016_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _18900_ (.A(_03018_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _18901_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.ready_buffer[11] ),
    .S(_03016_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _18902_ (.A(_03019_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _18903_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.ready_buffer[12] ),
    .S(_03016_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_1 _18904_ (.A(_03020_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _18905_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.ready_buffer[13] ),
    .S(_03016_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_1 _18906_ (.A(_03021_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _18907_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.ready_buffer[14] ),
    .S(_03016_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_1 _18908_ (.A(_03022_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _18909_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.ready_buffer[15] ),
    .S(_03016_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_1 _18910_ (.A(_03023_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _18911_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.ready_buffer[16] ),
    .S(_03016_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _18912_ (.A(_03024_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _18913_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.ready_buffer[17] ),
    .S(_03016_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_1 _18914_ (.A(_03025_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _18915_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.ready_buffer[18] ),
    .S(_03016_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_1 _18916_ (.A(_03026_),
    .X(_00665_));
 sky130_fd_sc_hd__clkbuf_4 _18917_ (.A(_03005_),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _18918_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.ready_buffer[19] ),
    .S(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _18919_ (.A(_03028_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _18920_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.ready_buffer[20] ),
    .S(_03027_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _18921_ (.A(_03029_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _18922_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.ready_buffer[21] ),
    .S(_03027_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _18923_ (.A(_03030_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _18924_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.ready_buffer[22] ),
    .S(_03027_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _18925_ (.A(_03031_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _18926_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.ready_buffer[23] ),
    .S(_03027_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _18927_ (.A(_03032_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _18928_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.ready_buffer[24] ),
    .S(_03027_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _18929_ (.A(_03033_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _18930_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.ready_buffer[25] ),
    .S(_03027_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _18931_ (.A(_03034_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _18932_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.ready_buffer[26] ),
    .S(_03027_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _18933_ (.A(_03035_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _18934_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.ready_buffer[27] ),
    .S(_03027_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_1 _18935_ (.A(_03036_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _18936_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.ready_buffer[28] ),
    .S(_03027_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_1 _18937_ (.A(_03037_),
    .X(_00675_));
 sky130_fd_sc_hd__clkbuf_4 _18938_ (.A(_03005_),
    .X(_03038_));
 sky130_fd_sc_hd__mux2_1 _18939_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.ready_buffer[29] ),
    .S(_03038_),
    .X(_03039_));
 sky130_fd_sc_hd__clkbuf_1 _18940_ (.A(_03039_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _18941_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.ready_buffer[30] ),
    .S(_03038_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _18942_ (.A(_03040_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _18943_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.ready_buffer[31] ),
    .S(_03038_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _18944_ (.A(_03041_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _18945_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.ready_buffer[32] ),
    .S(_03038_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _18946_ (.A(_03042_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _18947_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.ready_buffer[33] ),
    .S(_03038_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _18948_ (.A(_03043_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _18949_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.ready_buffer[34] ),
    .S(_03038_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_1 _18950_ (.A(_03044_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _18951_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.ready_buffer[35] ),
    .S(_03038_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _18952_ (.A(_03045_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _18953_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.ready_buffer[36] ),
    .S(_03038_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _18954_ (.A(_03046_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _18955_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.ready_buffer[37] ),
    .S(_03038_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_1 _18956_ (.A(_03047_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _18957_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.ready_buffer[38] ),
    .S(_03038_),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _18958_ (.A(_03048_),
    .X(_00685_));
 sky130_fd_sc_hd__buf_4 _18959_ (.A(_03005_),
    .X(_03049_));
 sky130_fd_sc_hd__mux2_1 _18960_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.ready_buffer[39] ),
    .S(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_1 _18961_ (.A(_03050_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _18962_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.ready_buffer[40] ),
    .S(_03049_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _18963_ (.A(_03051_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _18964_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.ready_buffer[41] ),
    .S(_03049_),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _18965_ (.A(_03052_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _18966_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.ready_buffer[42] ),
    .S(_03049_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _18967_ (.A(_03053_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _18968_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.ready_buffer[43] ),
    .S(_03049_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _18969_ (.A(_03054_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _18970_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_03049_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _18971_ (.A(_03055_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _18972_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.ready_buffer[45] ),
    .S(_03049_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _18973_ (.A(_03056_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _18974_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.ready_buffer[46] ),
    .S(_03049_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _18975_ (.A(_03057_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _18976_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.ready_buffer[47] ),
    .S(_03049_),
    .X(_03058_));
 sky130_fd_sc_hd__clkbuf_1 _18977_ (.A(_03058_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _18978_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.ready_buffer[48] ),
    .S(_03049_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_1 _18979_ (.A(_03059_),
    .X(_00695_));
 sky130_fd_sc_hd__clkbuf_4 _18980_ (.A(_03004_),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_1 _18981_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.ready_buffer[49] ),
    .S(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_1 _18982_ (.A(_03061_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _18983_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.ready_buffer[50] ),
    .S(_03060_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_1 _18984_ (.A(_03062_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _18985_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.ready_buffer[51] ),
    .S(_03060_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _18986_ (.A(_03063_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _18987_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.ready_buffer[52] ),
    .S(_03060_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _18988_ (.A(_03064_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _18989_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.ready_buffer[53] ),
    .S(_03060_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _18990_ (.A(_03065_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _18991_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.ready_buffer[54] ),
    .S(_03060_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _18992_ (.A(_03066_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _18993_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.ready_buffer[55] ),
    .S(_03060_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _18994_ (.A(_03067_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _18995_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.ready_buffer[56] ),
    .S(_03060_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _18996_ (.A(_03068_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _18997_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.ready_buffer[57] ),
    .S(_03060_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _18998_ (.A(_03069_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _18999_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.ready_buffer[58] ),
    .S(_03060_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _19000_ (.A(_03070_),
    .X(_00705_));
 sky130_fd_sc_hd__clkbuf_4 _19001_ (.A(_03004_),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _19002_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _19003_ (.A(_03072_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _19004_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.ready_buffer[60] ),
    .S(_03071_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _19005_ (.A(_03073_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _19006_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.ready_buffer[61] ),
    .S(_03071_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_1 _19007_ (.A(_03074_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _19008_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.ready_buffer[62] ),
    .S(_03071_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_1 _19009_ (.A(_03075_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _19010_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.ready_buffer[63] ),
    .S(_03071_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _19011_ (.A(_03076_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _19012_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.ready_buffer[64] ),
    .S(_03071_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_1 _19013_ (.A(_03077_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _19014_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.ready_buffer[65] ),
    .S(_03071_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _19015_ (.A(_03078_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _19016_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.ready_buffer[66] ),
    .S(_03071_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _19017_ (.A(_03079_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _19018_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.ready_buffer[67] ),
    .S(_03071_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _19019_ (.A(_03080_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _19020_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.ready_buffer[68] ),
    .S(_03071_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _19021_ (.A(_03081_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _19022_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.ready_buffer[69] ),
    .S(_03005_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _19023_ (.A(_03082_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _19024_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.ready_buffer[70] ),
    .S(_03005_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _19025_ (.A(_03083_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _19026_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.ready_buffer[71] ),
    .S(_03005_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_1 _19027_ (.A(_03084_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _19028_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.ready_buffer[72] ),
    .S(_03005_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _19029_ (.A(_03085_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _19030_ (.A0(\rbzero.pov.spi_buffer[73] ),
    .A1(\rbzero.pov.ready_buffer[73] ),
    .S(_03005_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _19031_ (.A(_03086_),
    .X(_00720_));
 sky130_fd_sc_hd__or4_1 _19032_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(\rbzero.spi_registers.spi_counter[3] ),
    .C(\rbzero.spi_registers.spi_counter[2] ),
    .D(_02983_),
    .X(_03087_));
 sky130_fd_sc_hd__and3_1 _19033_ (.A(_02989_),
    .B(_02966_),
    .C(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_4 _19034_ (.A(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__buf_4 _19035_ (.A(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__mux2_1 _19036_ (.A0(_02502_),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_03090_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _19037_ (.A(_03091_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _19038_ (.A0(_02509_),
    .A1(_02502_),
    .S(_03090_),
    .X(_03092_));
 sky130_fd_sc_hd__clkbuf_1 _19039_ (.A(_03092_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _19040_ (.A0(_02511_),
    .A1(_02509_),
    .S(_03090_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _19041_ (.A(_03093_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _19042_ (.A0(_02513_),
    .A1(_02511_),
    .S(_03090_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_1 _19043_ (.A(_03094_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _19044_ (.A0(_02515_),
    .A1(_02513_),
    .S(_03090_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_1 _19045_ (.A(_03095_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _19046_ (.A0(_02517_),
    .A1(_02515_),
    .S(_03090_),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _19047_ (.A(_03096_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _19048_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(_02517_),
    .S(_03090_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _19049_ (.A(_03097_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _19050_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03090_),
    .X(_03098_));
 sky130_fd_sc_hd__clkbuf_1 _19051_ (.A(_03098_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _19052_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03090_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _19053_ (.A(_03099_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _19054_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03090_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _19055_ (.A(_03100_),
    .X(_00730_));
 sky130_fd_sc_hd__buf_4 _19056_ (.A(_03089_),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _19057_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _19058_ (.A(_03102_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _19059_ (.A0(\rbzero.spi_registers.spi_buffer[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03101_),
    .X(_03103_));
 sky130_fd_sc_hd__clkbuf_1 _19060_ (.A(_03103_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _19061_ (.A0(\rbzero.spi_registers.spi_buffer[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03101_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _19062_ (.A(_03104_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _19063_ (.A0(\rbzero.spi_registers.spi_buffer[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03101_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _19064_ (.A(_03105_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _19065_ (.A0(\rbzero.spi_registers.spi_buffer[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03101_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _19066_ (.A(_03106_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _19067_ (.A0(\rbzero.spi_registers.spi_buffer[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03101_),
    .X(_03107_));
 sky130_fd_sc_hd__clkbuf_1 _19068_ (.A(_03107_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _19069_ (.A0(\rbzero.spi_registers.spi_buffer[16] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03101_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _19070_ (.A(_03108_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _19071_ (.A0(\rbzero.spi_registers.spi_buffer[17] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03101_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _19072_ (.A(_03109_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _19073_ (.A0(\rbzero.spi_registers.spi_buffer[18] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03101_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _19074_ (.A(_03110_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _19075_ (.A0(\rbzero.spi_registers.spi_buffer[19] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03101_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _19076_ (.A(_03111_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _19077_ (.A0(\rbzero.spi_registers.spi_buffer[20] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03089_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _19078_ (.A(_03112_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _19079_ (.A0(\rbzero.spi_registers.spi_buffer[21] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03089_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_1 _19080_ (.A(_03113_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _19081_ (.A0(\rbzero.spi_registers.spi_buffer[22] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03089_),
    .X(_03114_));
 sky130_fd_sc_hd__clkbuf_1 _19082_ (.A(_03114_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _19083_ (.A0(\rbzero.spi_registers.spi_buffer[23] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03089_),
    .X(_03115_));
 sky130_fd_sc_hd__clkbuf_1 _19084_ (.A(_03115_),
    .X(_00744_));
 sky130_fd_sc_hd__nand2_1 _19085_ (.A(_02989_),
    .B(_02966_),
    .Y(_03116_));
 sky130_fd_sc_hd__nor2_2 _19086_ (.A(_03087_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__mux2_1 _19087_ (.A0(\rbzero.spi_registers.spi_cmd[0] ),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _19088_ (.A(_03118_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _19089_ (.A0(_02503_),
    .A1(\rbzero.spi_registers.spi_cmd[0] ),
    .S(_03117_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _19090_ (.A(_03119_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _19091_ (.A0(\rbzero.spi_registers.spi_cmd[2] ),
    .A1(_02503_),
    .S(_03117_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _19092_ (.A(_03120_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _19093_ (.A0(\rbzero.spi_registers.spi_cmd[3] ),
    .A1(\rbzero.spi_registers.spi_cmd[2] ),
    .S(_03117_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_1 _19094_ (.A(_03121_),
    .X(_00748_));
 sky130_fd_sc_hd__buf_4 _19095_ (.A(_04469_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_1 _19096_ (.A0(net44),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__clkbuf_1 _19097_ (.A(_03123_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _19098_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_08185_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_1 _19099_ (.A(_03124_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _19100_ (.A0(net43),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_03122_),
    .X(_03125_));
 sky130_fd_sc_hd__clkbuf_1 _19101_ (.A(_03125_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _19102_ (.A0(\rbzero.spi_registers.ss_buffer[1] ),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_08185_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _19103_ (.A(_03126_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _19104_ (.A0(net46),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_03122_),
    .X(_03127_));
 sky130_fd_sc_hd__clkbuf_1 _19105_ (.A(_03127_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _19106_ (.A0(\rbzero.spi_registers.sclk_buffer[1] ),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_08185_),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _19107_ (.A(_03128_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _19108_ (.A0(\rbzero.spi_registers.sclk_buffer[1] ),
    .A1(\rbzero.spi_registers.sclk_buffer[2] ),
    .S(_03122_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _19109_ (.A(_03129_),
    .X(_00755_));
 sky130_fd_sc_hd__and3_1 _19110_ (.A(\gpout0.vpos[2] ),
    .B(_04744_),
    .C(\gpout0.vpos[0] ),
    .X(_03130_));
 sky130_fd_sc_hd__nand2_1 _19111_ (.A(_09805_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__nor2_1 _19112_ (.A(_04703_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__and2b_1 _19113_ (.A_N(_05762_),
    .B(_05761_),
    .X(_03133_));
 sky130_fd_sc_hd__and3_1 _19114_ (.A(_05756_),
    .B(_05755_),
    .C(_04729_),
    .X(_03134_));
 sky130_fd_sc_hd__and3_1 _19115_ (.A(_03132_),
    .B(_03133_),
    .C(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__buf_4 _19116_ (.A(_03135_),
    .X(_03136_));
 sky130_fd_sc_hd__nand2_4 _19117_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__and3_1 _19118_ (.A(_04723_),
    .B(_09805_),
    .C(_03130_),
    .X(_03138_));
 sky130_fd_sc_hd__and4_4 _19119_ (.A(_05758_),
    .B(_03133_),
    .C(_03134_),
    .D(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__buf_6 _19120_ (.A(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__and2_2 _19121_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__or2_1 _19122_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_4 _19123_ (.A(_09808_),
    .X(_03143_));
 sky130_fd_sc_hd__o211a_1 _19124_ (.A1(\rbzero.spi_registers.new_other[6] ),
    .A2(_03137_),
    .B1(_03142_),
    .C1(_03143_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _19125_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .B(_03141_),
    .X(_03144_));
 sky130_fd_sc_hd__o211a_1 _19126_ (.A1(\rbzero.spi_registers.new_other[7] ),
    .A2(_03137_),
    .B1(_03144_),
    .C1(_03143_),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _19127_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .B(_03141_),
    .X(_03145_));
 sky130_fd_sc_hd__o211a_1 _19128_ (.A1(\rbzero.spi_registers.new_other[8] ),
    .A2(_03137_),
    .B1(_03145_),
    .C1(_03143_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _19129_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .B(_03141_),
    .X(_03146_));
 sky130_fd_sc_hd__o211a_1 _19130_ (.A1(\rbzero.spi_registers.new_other[9] ),
    .A2(_03137_),
    .B1(_03146_),
    .C1(_03143_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _19131_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_03141_),
    .X(_03147_));
 sky130_fd_sc_hd__o211a_1 _19132_ (.A1(\rbzero.spi_registers.new_other[10] ),
    .A2(_03137_),
    .B1(_03147_),
    .C1(_03143_),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _19133_ (.A(\rbzero.map_overlay.i_othery[0] ),
    .B(_03141_),
    .X(_03148_));
 sky130_fd_sc_hd__o211a_1 _19134_ (.A1(\rbzero.spi_registers.new_other[0] ),
    .A2(_03137_),
    .B1(_03148_),
    .C1(_03143_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _19135_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(_03141_),
    .X(_03149_));
 sky130_fd_sc_hd__buf_4 _19136_ (.A(_04112_),
    .X(_03150_));
 sky130_fd_sc_hd__buf_2 _19137_ (.A(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__o211a_1 _19138_ (.A1(\rbzero.spi_registers.new_other[1] ),
    .A2(_03137_),
    .B1(_03149_),
    .C1(_03151_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _19139_ (.A(\rbzero.map_overlay.i_othery[2] ),
    .B(_03141_),
    .X(_03152_));
 sky130_fd_sc_hd__o211a_1 _19140_ (.A1(\rbzero.spi_registers.new_other[2] ),
    .A2(_03137_),
    .B1(_03152_),
    .C1(_03151_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _19141_ (.A(\rbzero.map_overlay.i_othery[3] ),
    .B(_03141_),
    .X(_03153_));
 sky130_fd_sc_hd__o211a_1 _19142_ (.A1(\rbzero.spi_registers.new_other[3] ),
    .A2(_03137_),
    .B1(_03153_),
    .C1(_03151_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _19143_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .B(_03141_),
    .X(_03154_));
 sky130_fd_sc_hd__o211a_1 _19144_ (.A1(\rbzero.spi_registers.new_other[4] ),
    .A2(_03137_),
    .B1(_03154_),
    .C1(_03151_),
    .X(_00765_));
 sky130_fd_sc_hd__inv_2 _19145_ (.A(\rbzero.spi_registers.got_new_vinf ),
    .Y(_03155_));
 sky130_fd_sc_hd__nand4_4 _19146_ (.A(_05758_),
    .B(_03133_),
    .C(_03134_),
    .D(_03138_),
    .Y(_03156_));
 sky130_fd_sc_hd__buf_2 _19147_ (.A(_03140_),
    .X(_03157_));
 sky130_fd_sc_hd__a21o_1 _19148_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_03157_),
    .B1(\rbzero.row_render.vinf ),
    .X(_03158_));
 sky130_fd_sc_hd__buf_4 _19149_ (.A(_08185_),
    .X(_03159_));
 sky130_fd_sc_hd__o311a_1 _19150_ (.A1(\rbzero.spi_registers.new_vinf ),
    .A2(_03155_),
    .A3(_03156_),
    .B1(_03158_),
    .C1(_03159_),
    .X(_00766_));
 sky130_fd_sc_hd__nand2_2 _19151_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_03136_),
    .Y(_03160_));
 sky130_fd_sc_hd__clkbuf_4 _19152_ (.A(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__and2_1 _19153_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_03139_),
    .X(_03162_));
 sky130_fd_sc_hd__clkbuf_2 _19154_ (.A(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__or2_1 _19155_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__o211a_1 _19156_ (.A1(net517),
    .A2(_03161_),
    .B1(_03164_),
    .C1(_03151_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _19157_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .B(_03163_),
    .X(_03165_));
 sky130_fd_sc_hd__o211a_1 _19158_ (.A1(\rbzero.spi_registers.new_mapd[11] ),
    .A2(_03161_),
    .B1(_03165_),
    .C1(_03151_),
    .X(_00768_));
 sky130_fd_sc_hd__or2_1 _19159_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_03163_),
    .X(_03166_));
 sky130_fd_sc_hd__o211a_1 _19160_ (.A1(\rbzero.spi_registers.new_mapd[12] ),
    .A2(_03161_),
    .B1(_03166_),
    .C1(_03151_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _19161_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_03163_),
    .X(_03167_));
 sky130_fd_sc_hd__o211a_1 _19162_ (.A1(\rbzero.spi_registers.new_mapd[13] ),
    .A2(_03161_),
    .B1(_03167_),
    .C1(_03151_),
    .X(_00770_));
 sky130_fd_sc_hd__or2_1 _19163_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .B(_03163_),
    .X(_03168_));
 sky130_fd_sc_hd__o211a_1 _19164_ (.A1(\rbzero.spi_registers.new_mapd[14] ),
    .A2(_03161_),
    .B1(_03168_),
    .C1(_03151_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _19165_ (.A(\rbzero.map_overlay.i_mapdx[5] ),
    .B(_03163_),
    .X(_03169_));
 sky130_fd_sc_hd__o211a_1 _19166_ (.A1(\rbzero.spi_registers.new_mapd[15] ),
    .A2(_03161_),
    .B1(_03169_),
    .C1(_03151_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _19167_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(_03163_),
    .X(_03170_));
 sky130_fd_sc_hd__buf_2 _19168_ (.A(_03150_),
    .X(_03171_));
 sky130_fd_sc_hd__o211a_1 _19169_ (.A1(net513),
    .A2(_03161_),
    .B1(_03170_),
    .C1(_03171_),
    .X(_00773_));
 sky130_fd_sc_hd__or2_1 _19170_ (.A(\rbzero.map_overlay.i_mapdy[1] ),
    .B(_03163_),
    .X(_03172_));
 sky130_fd_sc_hd__o211a_1 _19171_ (.A1(\rbzero.spi_registers.new_mapd[5] ),
    .A2(_03161_),
    .B1(_03172_),
    .C1(_03171_),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _19172_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(_03163_),
    .X(_03173_));
 sky130_fd_sc_hd__o211a_1 _19173_ (.A1(\rbzero.spi_registers.new_mapd[6] ),
    .A2(_03161_),
    .B1(_03173_),
    .C1(_03171_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _19174_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(_03163_),
    .X(_03174_));
 sky130_fd_sc_hd__o211a_1 _19175_ (.A1(\rbzero.spi_registers.new_mapd[7] ),
    .A2(_03161_),
    .B1(_03174_),
    .C1(_03171_),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _19176_ (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .B(_03162_),
    .X(_03175_));
 sky130_fd_sc_hd__o211a_1 _19177_ (.A1(\rbzero.spi_registers.new_mapd[8] ),
    .A2(_03160_),
    .B1(_03175_),
    .C1(_03171_),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _19178_ (.A(\rbzero.map_overlay.i_mapdy[5] ),
    .B(_03162_),
    .X(_03176_));
 sky130_fd_sc_hd__o211a_1 _19179_ (.A1(\rbzero.spi_registers.new_mapd[9] ),
    .A2(_03160_),
    .B1(_03176_),
    .C1(_03171_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _19180_ (.A(\rbzero.mapdxw[0] ),
    .B(_03162_),
    .X(_03177_));
 sky130_fd_sc_hd__o211a_1 _19181_ (.A1(\rbzero.spi_registers.new_mapd[2] ),
    .A2(_03160_),
    .B1(_03177_),
    .C1(_03171_),
    .X(_00779_));
 sky130_fd_sc_hd__or2_1 _19182_ (.A(\rbzero.mapdxw[1] ),
    .B(_03162_),
    .X(_03178_));
 sky130_fd_sc_hd__o211a_1 _19183_ (.A1(\rbzero.spi_registers.new_mapd[3] ),
    .A2(_03160_),
    .B1(_03178_),
    .C1(_03171_),
    .X(_00780_));
 sky130_fd_sc_hd__or2_1 _19184_ (.A(\rbzero.mapdyw[0] ),
    .B(_03162_),
    .X(_03179_));
 sky130_fd_sc_hd__o211a_1 _19185_ (.A1(\rbzero.spi_registers.new_mapd[0] ),
    .A2(_03160_),
    .B1(_03179_),
    .C1(_03171_),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _19186_ (.A(\rbzero.mapdyw[1] ),
    .B(_03162_),
    .X(_03180_));
 sky130_fd_sc_hd__o211a_1 _19187_ (.A1(\rbzero.spi_registers.new_mapd[1] ),
    .A2(_03160_),
    .B1(_03180_),
    .C1(_03171_),
    .X(_00782_));
 sky130_fd_sc_hd__nand2_2 _19188_ (.A(\rbzero.spi_registers.got_new_texadd[0] ),
    .B(_03136_),
    .Y(_03181_));
 sky130_fd_sc_hd__clkbuf_4 _19189_ (.A(_03181_),
    .X(_03182_));
 sky130_fd_sc_hd__and2_2 _19190_ (.A(\rbzero.spi_registers.got_new_texadd[0] ),
    .B(_03140_),
    .X(_03183_));
 sky130_fd_sc_hd__buf_2 _19191_ (.A(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__or2_1 _19192_ (.A(\rbzero.spi_registers.texadd0[0] ),
    .B(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__buf_2 _19193_ (.A(_03150_),
    .X(_03186_));
 sky130_fd_sc_hd__o211a_1 _19194_ (.A1(\rbzero.spi_registers.new_texadd[0][0] ),
    .A2(_03182_),
    .B1(_03185_),
    .C1(_03186_),
    .X(_00783_));
 sky130_fd_sc_hd__or2_1 _19195_ (.A(\rbzero.spi_registers.texadd0[1] ),
    .B(_03184_),
    .X(_03187_));
 sky130_fd_sc_hd__o211a_1 _19196_ (.A1(\rbzero.spi_registers.new_texadd[0][1] ),
    .A2(_03182_),
    .B1(_03187_),
    .C1(_03186_),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _19197_ (.A(\rbzero.spi_registers.texadd0[2] ),
    .B(_03184_),
    .X(_03188_));
 sky130_fd_sc_hd__o211a_1 _19198_ (.A1(\rbzero.spi_registers.new_texadd[0][2] ),
    .A2(_03182_),
    .B1(_03188_),
    .C1(_03186_),
    .X(_00785_));
 sky130_fd_sc_hd__or2_1 _19199_ (.A(\rbzero.spi_registers.texadd0[3] ),
    .B(_03184_),
    .X(_03189_));
 sky130_fd_sc_hd__o211a_1 _19200_ (.A1(\rbzero.spi_registers.new_texadd[0][3] ),
    .A2(_03182_),
    .B1(_03189_),
    .C1(_03186_),
    .X(_00786_));
 sky130_fd_sc_hd__or2_1 _19201_ (.A(\rbzero.spi_registers.texadd0[4] ),
    .B(_03184_),
    .X(_03190_));
 sky130_fd_sc_hd__o211a_1 _19202_ (.A1(\rbzero.spi_registers.new_texadd[0][4] ),
    .A2(_03182_),
    .B1(_03190_),
    .C1(_03186_),
    .X(_00787_));
 sky130_fd_sc_hd__or2_1 _19203_ (.A(\rbzero.spi_registers.texadd0[5] ),
    .B(_03184_),
    .X(_03191_));
 sky130_fd_sc_hd__o211a_1 _19204_ (.A1(\rbzero.spi_registers.new_texadd[0][5] ),
    .A2(_03182_),
    .B1(_03191_),
    .C1(_03186_),
    .X(_00788_));
 sky130_fd_sc_hd__or2_1 _19205_ (.A(\rbzero.spi_registers.texadd0[6] ),
    .B(_03184_),
    .X(_03192_));
 sky130_fd_sc_hd__o211a_1 _19206_ (.A1(\rbzero.spi_registers.new_texadd[0][6] ),
    .A2(_03182_),
    .B1(_03192_),
    .C1(_03186_),
    .X(_00789_));
 sky130_fd_sc_hd__or2_1 _19207_ (.A(\rbzero.spi_registers.texadd0[7] ),
    .B(_03184_),
    .X(_03193_));
 sky130_fd_sc_hd__o211a_1 _19208_ (.A1(\rbzero.spi_registers.new_texadd[0][7] ),
    .A2(_03182_),
    .B1(_03193_),
    .C1(_03186_),
    .X(_00790_));
 sky130_fd_sc_hd__or2_1 _19209_ (.A(\rbzero.spi_registers.texadd0[8] ),
    .B(_03184_),
    .X(_03194_));
 sky130_fd_sc_hd__o211a_1 _19210_ (.A1(\rbzero.spi_registers.new_texadd[0][8] ),
    .A2(_03182_),
    .B1(_03194_),
    .C1(_03186_),
    .X(_00791_));
 sky130_fd_sc_hd__or2_1 _19211_ (.A(\rbzero.spi_registers.texadd0[9] ),
    .B(_03184_),
    .X(_03195_));
 sky130_fd_sc_hd__o211a_1 _19212_ (.A1(\rbzero.spi_registers.new_texadd[0][9] ),
    .A2(_03182_),
    .B1(_03195_),
    .C1(_03186_),
    .X(_00792_));
 sky130_fd_sc_hd__clkbuf_4 _19213_ (.A(_03181_),
    .X(_03196_));
 sky130_fd_sc_hd__buf_2 _19214_ (.A(_03183_),
    .X(_03197_));
 sky130_fd_sc_hd__or2_1 _19215_ (.A(\rbzero.spi_registers.texadd0[10] ),
    .B(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__buf_2 _19216_ (.A(_03150_),
    .X(_03199_));
 sky130_fd_sc_hd__o211a_1 _19217_ (.A1(\rbzero.spi_registers.new_texadd[0][10] ),
    .A2(_03196_),
    .B1(_03198_),
    .C1(_03199_),
    .X(_00793_));
 sky130_fd_sc_hd__or2_1 _19218_ (.A(\rbzero.spi_registers.texadd0[11] ),
    .B(_03197_),
    .X(_03200_));
 sky130_fd_sc_hd__o211a_1 _19219_ (.A1(\rbzero.spi_registers.new_texadd[0][11] ),
    .A2(_03196_),
    .B1(_03200_),
    .C1(_03199_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _19220_ (.A(\rbzero.spi_registers.texadd0[12] ),
    .B(_03197_),
    .X(_03201_));
 sky130_fd_sc_hd__o211a_1 _19221_ (.A1(\rbzero.spi_registers.new_texadd[0][12] ),
    .A2(_03196_),
    .B1(_03201_),
    .C1(_03199_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _19222_ (.A(\rbzero.spi_registers.texadd0[13] ),
    .B(_03197_),
    .X(_03202_));
 sky130_fd_sc_hd__o211a_1 _19223_ (.A1(\rbzero.spi_registers.new_texadd[0][13] ),
    .A2(_03196_),
    .B1(_03202_),
    .C1(_03199_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _19224_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_03197_),
    .X(_03203_));
 sky130_fd_sc_hd__o211a_1 _19225_ (.A1(\rbzero.spi_registers.new_texadd[0][14] ),
    .A2(_03196_),
    .B1(_03203_),
    .C1(_03199_),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _19226_ (.A(\rbzero.spi_registers.texadd0[15] ),
    .B(_03197_),
    .X(_03204_));
 sky130_fd_sc_hd__o211a_1 _19227_ (.A1(\rbzero.spi_registers.new_texadd[0][15] ),
    .A2(_03196_),
    .B1(_03204_),
    .C1(_03199_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _19228_ (.A(\rbzero.spi_registers.texadd0[16] ),
    .B(_03197_),
    .X(_03205_));
 sky130_fd_sc_hd__o211a_1 _19229_ (.A1(\rbzero.spi_registers.new_texadd[0][16] ),
    .A2(_03196_),
    .B1(_03205_),
    .C1(_03199_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _19230_ (.A(\rbzero.spi_registers.texadd0[17] ),
    .B(_03197_),
    .X(_03206_));
 sky130_fd_sc_hd__o211a_1 _19231_ (.A1(\rbzero.spi_registers.new_texadd[0][17] ),
    .A2(_03196_),
    .B1(_03206_),
    .C1(_03199_),
    .X(_00800_));
 sky130_fd_sc_hd__or2_1 _19232_ (.A(\rbzero.spi_registers.texadd0[18] ),
    .B(_03197_),
    .X(_03207_));
 sky130_fd_sc_hd__o211a_1 _19233_ (.A1(\rbzero.spi_registers.new_texadd[0][18] ),
    .A2(_03196_),
    .B1(_03207_),
    .C1(_03199_),
    .X(_00801_));
 sky130_fd_sc_hd__or2_1 _19234_ (.A(\rbzero.spi_registers.texadd0[19] ),
    .B(_03197_),
    .X(_03208_));
 sky130_fd_sc_hd__o211a_1 _19235_ (.A1(\rbzero.spi_registers.new_texadd[0][19] ),
    .A2(_03196_),
    .B1(_03208_),
    .C1(_03199_),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _19236_ (.A(\rbzero.spi_registers.texadd0[20] ),
    .B(_03183_),
    .X(_03209_));
 sky130_fd_sc_hd__clkbuf_4 _19237_ (.A(_03150_),
    .X(_03210_));
 sky130_fd_sc_hd__o211a_1 _19238_ (.A1(\rbzero.spi_registers.new_texadd[0][20] ),
    .A2(_03181_),
    .B1(_03209_),
    .C1(_03210_),
    .X(_00803_));
 sky130_fd_sc_hd__or2_1 _19239_ (.A(\rbzero.spi_registers.texadd0[21] ),
    .B(_03183_),
    .X(_03211_));
 sky130_fd_sc_hd__o211a_1 _19240_ (.A1(\rbzero.spi_registers.new_texadd[0][21] ),
    .A2(_03181_),
    .B1(_03211_),
    .C1(_03210_),
    .X(_00804_));
 sky130_fd_sc_hd__or2_1 _19241_ (.A(\rbzero.spi_registers.texadd0[22] ),
    .B(_03183_),
    .X(_03212_));
 sky130_fd_sc_hd__o211a_1 _19242_ (.A1(\rbzero.spi_registers.new_texadd[0][22] ),
    .A2(_03181_),
    .B1(_03212_),
    .C1(_03210_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _19243_ (.A(\rbzero.spi_registers.texadd0[23] ),
    .B(_03183_),
    .X(_03213_));
 sky130_fd_sc_hd__o211a_1 _19244_ (.A1(\rbzero.spi_registers.new_texadd[0][23] ),
    .A2(_03181_),
    .B1(_03213_),
    .C1(_03210_),
    .X(_00806_));
 sky130_fd_sc_hd__nand2_2 _19245_ (.A(\rbzero.spi_registers.got_new_texadd[1] ),
    .B(_03136_),
    .Y(_03214_));
 sky130_fd_sc_hd__clkbuf_4 _19246_ (.A(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__and2_1 _19247_ (.A(\rbzero.spi_registers.got_new_texadd[1] ),
    .B(_03139_),
    .X(_03216_));
 sky130_fd_sc_hd__buf_2 _19248_ (.A(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__or2_1 _19249_ (.A(\rbzero.spi_registers.texadd1[0] ),
    .B(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__o211a_1 _19250_ (.A1(\rbzero.spi_registers.new_texadd[1][0] ),
    .A2(_03215_),
    .B1(_03218_),
    .C1(_03210_),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _19251_ (.A(\rbzero.spi_registers.texadd1[1] ),
    .B(_03217_),
    .X(_03219_));
 sky130_fd_sc_hd__o211a_1 _19252_ (.A1(\rbzero.spi_registers.new_texadd[1][1] ),
    .A2(_03215_),
    .B1(_03219_),
    .C1(_03210_),
    .X(_00808_));
 sky130_fd_sc_hd__or2_1 _19253_ (.A(\rbzero.spi_registers.texadd1[2] ),
    .B(_03217_),
    .X(_03220_));
 sky130_fd_sc_hd__o211a_1 _19254_ (.A1(\rbzero.spi_registers.new_texadd[1][2] ),
    .A2(_03215_),
    .B1(_03220_),
    .C1(_03210_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _19255_ (.A(\rbzero.spi_registers.texadd1[3] ),
    .B(_03217_),
    .X(_03221_));
 sky130_fd_sc_hd__o211a_1 _19256_ (.A1(\rbzero.spi_registers.new_texadd[1][3] ),
    .A2(_03215_),
    .B1(_03221_),
    .C1(_03210_),
    .X(_00810_));
 sky130_fd_sc_hd__or2_1 _19257_ (.A(\rbzero.spi_registers.texadd1[4] ),
    .B(_03217_),
    .X(_03222_));
 sky130_fd_sc_hd__o211a_1 _19258_ (.A1(\rbzero.spi_registers.new_texadd[1][4] ),
    .A2(_03215_),
    .B1(_03222_),
    .C1(_03210_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _19259_ (.A(\rbzero.spi_registers.texadd1[5] ),
    .B(_03217_),
    .X(_03223_));
 sky130_fd_sc_hd__o211a_1 _19260_ (.A1(\rbzero.spi_registers.new_texadd[1][5] ),
    .A2(_03215_),
    .B1(_03223_),
    .C1(_03210_),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _19261_ (.A(\rbzero.spi_registers.texadd1[6] ),
    .B(_03217_),
    .X(_03224_));
 sky130_fd_sc_hd__clkbuf_4 _19262_ (.A(_03150_),
    .X(_03225_));
 sky130_fd_sc_hd__o211a_1 _19263_ (.A1(\rbzero.spi_registers.new_texadd[1][6] ),
    .A2(_03215_),
    .B1(_03224_),
    .C1(_03225_),
    .X(_00813_));
 sky130_fd_sc_hd__or2_1 _19264_ (.A(\rbzero.spi_registers.texadd1[7] ),
    .B(_03217_),
    .X(_03226_));
 sky130_fd_sc_hd__o211a_1 _19265_ (.A1(\rbzero.spi_registers.new_texadd[1][7] ),
    .A2(_03215_),
    .B1(_03226_),
    .C1(_03225_),
    .X(_00814_));
 sky130_fd_sc_hd__or2_1 _19266_ (.A(\rbzero.spi_registers.texadd1[8] ),
    .B(_03217_),
    .X(_03227_));
 sky130_fd_sc_hd__o211a_1 _19267_ (.A1(\rbzero.spi_registers.new_texadd[1][8] ),
    .A2(_03215_),
    .B1(_03227_),
    .C1(_03225_),
    .X(_00815_));
 sky130_fd_sc_hd__or2_1 _19268_ (.A(\rbzero.spi_registers.texadd1[9] ),
    .B(_03217_),
    .X(_03228_));
 sky130_fd_sc_hd__o211a_1 _19269_ (.A1(\rbzero.spi_registers.new_texadd[1][9] ),
    .A2(_03215_),
    .B1(_03228_),
    .C1(_03225_),
    .X(_00816_));
 sky130_fd_sc_hd__clkbuf_4 _19270_ (.A(_03214_),
    .X(_03229_));
 sky130_fd_sc_hd__buf_2 _19271_ (.A(_03216_),
    .X(_03230_));
 sky130_fd_sc_hd__or2_1 _19272_ (.A(\rbzero.spi_registers.texadd1[10] ),
    .B(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__o211a_1 _19273_ (.A1(\rbzero.spi_registers.new_texadd[1][10] ),
    .A2(_03229_),
    .B1(_03231_),
    .C1(_03225_),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _19274_ (.A(\rbzero.spi_registers.texadd1[11] ),
    .B(_03230_),
    .X(_03232_));
 sky130_fd_sc_hd__o211a_1 _19275_ (.A1(\rbzero.spi_registers.new_texadd[1][11] ),
    .A2(_03229_),
    .B1(_03232_),
    .C1(_03225_),
    .X(_00818_));
 sky130_fd_sc_hd__or2_1 _19276_ (.A(\rbzero.spi_registers.texadd1[12] ),
    .B(_03230_),
    .X(_03233_));
 sky130_fd_sc_hd__o211a_1 _19277_ (.A1(\rbzero.spi_registers.new_texadd[1][12] ),
    .A2(_03229_),
    .B1(_03233_),
    .C1(_03225_),
    .X(_00819_));
 sky130_fd_sc_hd__or2_1 _19278_ (.A(\rbzero.spi_registers.texadd1[13] ),
    .B(_03230_),
    .X(_03234_));
 sky130_fd_sc_hd__o211a_1 _19279_ (.A1(\rbzero.spi_registers.new_texadd[1][13] ),
    .A2(_03229_),
    .B1(_03234_),
    .C1(_03225_),
    .X(_00820_));
 sky130_fd_sc_hd__or2_1 _19280_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .B(_03230_),
    .X(_03235_));
 sky130_fd_sc_hd__o211a_1 _19281_ (.A1(\rbzero.spi_registers.new_texadd[1][14] ),
    .A2(_03229_),
    .B1(_03235_),
    .C1(_03225_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _19282_ (.A(\rbzero.spi_registers.texadd1[15] ),
    .B(_03230_),
    .X(_03236_));
 sky130_fd_sc_hd__o211a_1 _19283_ (.A1(\rbzero.spi_registers.new_texadd[1][15] ),
    .A2(_03229_),
    .B1(_03236_),
    .C1(_03225_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _19284_ (.A(\rbzero.spi_registers.texadd1[16] ),
    .B(_03230_),
    .X(_03237_));
 sky130_fd_sc_hd__clkbuf_4 _19285_ (.A(_03150_),
    .X(_03238_));
 sky130_fd_sc_hd__o211a_1 _19286_ (.A1(\rbzero.spi_registers.new_texadd[1][16] ),
    .A2(_03229_),
    .B1(_03237_),
    .C1(_03238_),
    .X(_00823_));
 sky130_fd_sc_hd__or2_1 _19287_ (.A(\rbzero.spi_registers.texadd1[17] ),
    .B(_03230_),
    .X(_03239_));
 sky130_fd_sc_hd__o211a_1 _19288_ (.A1(\rbzero.spi_registers.new_texadd[1][17] ),
    .A2(_03229_),
    .B1(_03239_),
    .C1(_03238_),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _19289_ (.A(\rbzero.spi_registers.texadd1[18] ),
    .B(_03230_),
    .X(_03240_));
 sky130_fd_sc_hd__o211a_1 _19290_ (.A1(\rbzero.spi_registers.new_texadd[1][18] ),
    .A2(_03229_),
    .B1(_03240_),
    .C1(_03238_),
    .X(_00825_));
 sky130_fd_sc_hd__or2_1 _19291_ (.A(\rbzero.spi_registers.texadd1[19] ),
    .B(_03230_),
    .X(_03241_));
 sky130_fd_sc_hd__o211a_1 _19292_ (.A1(\rbzero.spi_registers.new_texadd[1][19] ),
    .A2(_03229_),
    .B1(_03241_),
    .C1(_03238_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _19293_ (.A(\rbzero.spi_registers.texadd1[20] ),
    .B(_03216_),
    .X(_03242_));
 sky130_fd_sc_hd__o211a_1 _19294_ (.A1(\rbzero.spi_registers.new_texadd[1][20] ),
    .A2(_03214_),
    .B1(_03242_),
    .C1(_03238_),
    .X(_00827_));
 sky130_fd_sc_hd__or2_1 _19295_ (.A(\rbzero.spi_registers.texadd1[21] ),
    .B(_03216_),
    .X(_03243_));
 sky130_fd_sc_hd__o211a_1 _19296_ (.A1(\rbzero.spi_registers.new_texadd[1][21] ),
    .A2(_03214_),
    .B1(_03243_),
    .C1(_03238_),
    .X(_00828_));
 sky130_fd_sc_hd__or2_1 _19297_ (.A(\rbzero.spi_registers.texadd1[22] ),
    .B(_03216_),
    .X(_03244_));
 sky130_fd_sc_hd__o211a_1 _19298_ (.A1(\rbzero.spi_registers.new_texadd[1][22] ),
    .A2(_03214_),
    .B1(_03244_),
    .C1(_03238_),
    .X(_00829_));
 sky130_fd_sc_hd__or2_1 _19299_ (.A(\rbzero.spi_registers.texadd1[23] ),
    .B(_03216_),
    .X(_03245_));
 sky130_fd_sc_hd__o211a_1 _19300_ (.A1(\rbzero.spi_registers.new_texadd[1][23] ),
    .A2(_03214_),
    .B1(_03245_),
    .C1(_03238_),
    .X(_00830_));
 sky130_fd_sc_hd__nand2_2 _19301_ (.A(\rbzero.spi_registers.got_new_texadd[2] ),
    .B(_03136_),
    .Y(_03246_));
 sky130_fd_sc_hd__clkbuf_4 _19302_ (.A(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__and2_1 _19303_ (.A(\rbzero.spi_registers.got_new_texadd[2] ),
    .B(_03139_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_2 _19304_ (.A(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__or2_1 _19305_ (.A(\rbzero.spi_registers.texadd2[0] ),
    .B(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__o211a_1 _19306_ (.A1(\rbzero.spi_registers.new_texadd[2][0] ),
    .A2(_03247_),
    .B1(_03250_),
    .C1(_03238_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _19307_ (.A(\rbzero.spi_registers.texadd2[1] ),
    .B(_03249_),
    .X(_03251_));
 sky130_fd_sc_hd__o211a_1 _19308_ (.A1(\rbzero.spi_registers.new_texadd[2][1] ),
    .A2(_03247_),
    .B1(_03251_),
    .C1(_03238_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _19309_ (.A(\rbzero.spi_registers.texadd2[2] ),
    .B(_03249_),
    .X(_03252_));
 sky130_fd_sc_hd__clkbuf_4 _19310_ (.A(_03150_),
    .X(_03253_));
 sky130_fd_sc_hd__o211a_1 _19311_ (.A1(\rbzero.spi_registers.new_texadd[2][2] ),
    .A2(_03247_),
    .B1(_03252_),
    .C1(_03253_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_1 _19312_ (.A(\rbzero.spi_registers.texadd2[3] ),
    .B(_03249_),
    .X(_03254_));
 sky130_fd_sc_hd__o211a_1 _19313_ (.A1(\rbzero.spi_registers.new_texadd[2][3] ),
    .A2(_03247_),
    .B1(_03254_),
    .C1(_03253_),
    .X(_00834_));
 sky130_fd_sc_hd__or2_1 _19314_ (.A(\rbzero.spi_registers.texadd2[4] ),
    .B(_03249_),
    .X(_03255_));
 sky130_fd_sc_hd__o211a_1 _19315_ (.A1(\rbzero.spi_registers.new_texadd[2][4] ),
    .A2(_03247_),
    .B1(_03255_),
    .C1(_03253_),
    .X(_00835_));
 sky130_fd_sc_hd__or2_1 _19316_ (.A(\rbzero.spi_registers.texadd2[5] ),
    .B(_03249_),
    .X(_03256_));
 sky130_fd_sc_hd__o211a_1 _19317_ (.A1(\rbzero.spi_registers.new_texadd[2][5] ),
    .A2(_03247_),
    .B1(_03256_),
    .C1(_03253_),
    .X(_00836_));
 sky130_fd_sc_hd__or2_1 _19318_ (.A(\rbzero.spi_registers.texadd2[6] ),
    .B(_03249_),
    .X(_03257_));
 sky130_fd_sc_hd__o211a_1 _19319_ (.A1(\rbzero.spi_registers.new_texadd[2][6] ),
    .A2(_03247_),
    .B1(_03257_),
    .C1(_03253_),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _19320_ (.A(\rbzero.spi_registers.texadd2[7] ),
    .B(_03249_),
    .X(_03258_));
 sky130_fd_sc_hd__o211a_1 _19321_ (.A1(\rbzero.spi_registers.new_texadd[2][7] ),
    .A2(_03247_),
    .B1(_03258_),
    .C1(_03253_),
    .X(_00838_));
 sky130_fd_sc_hd__or2_1 _19322_ (.A(\rbzero.spi_registers.texadd2[8] ),
    .B(_03249_),
    .X(_03259_));
 sky130_fd_sc_hd__o211a_1 _19323_ (.A1(\rbzero.spi_registers.new_texadd[2][8] ),
    .A2(_03247_),
    .B1(_03259_),
    .C1(_03253_),
    .X(_00839_));
 sky130_fd_sc_hd__or2_1 _19324_ (.A(\rbzero.spi_registers.texadd2[9] ),
    .B(_03249_),
    .X(_03260_));
 sky130_fd_sc_hd__o211a_1 _19325_ (.A1(\rbzero.spi_registers.new_texadd[2][9] ),
    .A2(_03247_),
    .B1(_03260_),
    .C1(_03253_),
    .X(_00840_));
 sky130_fd_sc_hd__clkbuf_4 _19326_ (.A(_03246_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_2 _19327_ (.A(_03248_),
    .X(_03262_));
 sky130_fd_sc_hd__or2_1 _19328_ (.A(\rbzero.spi_registers.texadd2[10] ),
    .B(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__o211a_1 _19329_ (.A1(\rbzero.spi_registers.new_texadd[2][10] ),
    .A2(_03261_),
    .B1(_03263_),
    .C1(_03253_),
    .X(_00841_));
 sky130_fd_sc_hd__or2_1 _19330_ (.A(\rbzero.spi_registers.texadd2[11] ),
    .B(_03262_),
    .X(_03264_));
 sky130_fd_sc_hd__o211a_1 _19331_ (.A1(\rbzero.spi_registers.new_texadd[2][11] ),
    .A2(_03261_),
    .B1(_03264_),
    .C1(_03253_),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _19332_ (.A(\rbzero.spi_registers.texadd2[12] ),
    .B(_03262_),
    .X(_03265_));
 sky130_fd_sc_hd__clkbuf_4 _19333_ (.A(_03150_),
    .X(_03266_));
 sky130_fd_sc_hd__o211a_1 _19334_ (.A1(\rbzero.spi_registers.new_texadd[2][12] ),
    .A2(_03261_),
    .B1(_03265_),
    .C1(_03266_),
    .X(_00843_));
 sky130_fd_sc_hd__or2_1 _19335_ (.A(\rbzero.spi_registers.texadd2[13] ),
    .B(_03262_),
    .X(_03267_));
 sky130_fd_sc_hd__o211a_1 _19336_ (.A1(\rbzero.spi_registers.new_texadd[2][13] ),
    .A2(_03261_),
    .B1(_03267_),
    .C1(_03266_),
    .X(_00844_));
 sky130_fd_sc_hd__or2_1 _19337_ (.A(\rbzero.spi_registers.texadd2[14] ),
    .B(_03262_),
    .X(_03268_));
 sky130_fd_sc_hd__o211a_1 _19338_ (.A1(\rbzero.spi_registers.new_texadd[2][14] ),
    .A2(_03261_),
    .B1(_03268_),
    .C1(_03266_),
    .X(_00845_));
 sky130_fd_sc_hd__or2_1 _19339_ (.A(\rbzero.spi_registers.texadd2[15] ),
    .B(_03262_),
    .X(_03269_));
 sky130_fd_sc_hd__o211a_1 _19340_ (.A1(\rbzero.spi_registers.new_texadd[2][15] ),
    .A2(_03261_),
    .B1(_03269_),
    .C1(_03266_),
    .X(_00846_));
 sky130_fd_sc_hd__or2_1 _19341_ (.A(\rbzero.spi_registers.texadd2[16] ),
    .B(_03262_),
    .X(_03270_));
 sky130_fd_sc_hd__o211a_1 _19342_ (.A1(\rbzero.spi_registers.new_texadd[2][16] ),
    .A2(_03261_),
    .B1(_03270_),
    .C1(_03266_),
    .X(_00847_));
 sky130_fd_sc_hd__or2_1 _19343_ (.A(\rbzero.spi_registers.texadd2[17] ),
    .B(_03262_),
    .X(_03271_));
 sky130_fd_sc_hd__o211a_1 _19344_ (.A1(\rbzero.spi_registers.new_texadd[2][17] ),
    .A2(_03261_),
    .B1(_03271_),
    .C1(_03266_),
    .X(_00848_));
 sky130_fd_sc_hd__or2_1 _19345_ (.A(\rbzero.spi_registers.texadd2[18] ),
    .B(_03262_),
    .X(_03272_));
 sky130_fd_sc_hd__o211a_1 _19346_ (.A1(\rbzero.spi_registers.new_texadd[2][18] ),
    .A2(_03261_),
    .B1(_03272_),
    .C1(_03266_),
    .X(_00849_));
 sky130_fd_sc_hd__or2_1 _19347_ (.A(\rbzero.spi_registers.texadd2[19] ),
    .B(_03262_),
    .X(_03273_));
 sky130_fd_sc_hd__o211a_1 _19348_ (.A1(\rbzero.spi_registers.new_texadd[2][19] ),
    .A2(_03261_),
    .B1(_03273_),
    .C1(_03266_),
    .X(_00850_));
 sky130_fd_sc_hd__or2_1 _19349_ (.A(\rbzero.spi_registers.texadd2[20] ),
    .B(_03248_),
    .X(_03274_));
 sky130_fd_sc_hd__o211a_1 _19350_ (.A1(\rbzero.spi_registers.new_texadd[2][20] ),
    .A2(_03246_),
    .B1(_03274_),
    .C1(_03266_),
    .X(_00851_));
 sky130_fd_sc_hd__or2_1 _19351_ (.A(\rbzero.spi_registers.texadd2[21] ),
    .B(_03248_),
    .X(_03275_));
 sky130_fd_sc_hd__o211a_1 _19352_ (.A1(\rbzero.spi_registers.new_texadd[2][21] ),
    .A2(_03246_),
    .B1(_03275_),
    .C1(_03266_),
    .X(_00852_));
 sky130_fd_sc_hd__or2_1 _19353_ (.A(\rbzero.spi_registers.texadd2[22] ),
    .B(_03248_),
    .X(_03276_));
 sky130_fd_sc_hd__clkbuf_4 _19354_ (.A(_09808_),
    .X(_03277_));
 sky130_fd_sc_hd__o211a_1 _19355_ (.A1(\rbzero.spi_registers.new_texadd[2][22] ),
    .A2(_03246_),
    .B1(_03276_),
    .C1(_03277_),
    .X(_00853_));
 sky130_fd_sc_hd__or2_1 _19356_ (.A(\rbzero.spi_registers.texadd2[23] ),
    .B(_03248_),
    .X(_03278_));
 sky130_fd_sc_hd__o211a_1 _19357_ (.A1(\rbzero.spi_registers.new_texadd[2][23] ),
    .A2(_03246_),
    .B1(_03278_),
    .C1(_03277_),
    .X(_00854_));
 sky130_fd_sc_hd__nand2_2 _19358_ (.A(\rbzero.spi_registers.got_new_texadd[3] ),
    .B(_03136_),
    .Y(_03279_));
 sky130_fd_sc_hd__clkbuf_4 _19359_ (.A(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__and2_1 _19360_ (.A(\rbzero.spi_registers.got_new_texadd[3] ),
    .B(_03139_),
    .X(_03281_));
 sky130_fd_sc_hd__buf_2 _19361_ (.A(_03281_),
    .X(_03282_));
 sky130_fd_sc_hd__or2_1 _19362_ (.A(\rbzero.spi_registers.texadd3[0] ),
    .B(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__o211a_1 _19363_ (.A1(\rbzero.spi_registers.new_texadd[3][0] ),
    .A2(_03280_),
    .B1(_03283_),
    .C1(_03277_),
    .X(_00855_));
 sky130_fd_sc_hd__or2_1 _19364_ (.A(\rbzero.spi_registers.texadd3[1] ),
    .B(_03282_),
    .X(_03284_));
 sky130_fd_sc_hd__o211a_1 _19365_ (.A1(\rbzero.spi_registers.new_texadd[3][1] ),
    .A2(_03280_),
    .B1(_03284_),
    .C1(_03277_),
    .X(_00856_));
 sky130_fd_sc_hd__or2_1 _19366_ (.A(\rbzero.spi_registers.texadd3[2] ),
    .B(_03282_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_1 _19367_ (.A1(\rbzero.spi_registers.new_texadd[3][2] ),
    .A2(_03280_),
    .B1(_03285_),
    .C1(_03277_),
    .X(_00857_));
 sky130_fd_sc_hd__or2_1 _19368_ (.A(\rbzero.spi_registers.texadd3[3] ),
    .B(_03282_),
    .X(_03286_));
 sky130_fd_sc_hd__o211a_1 _19369_ (.A1(\rbzero.spi_registers.new_texadd[3][3] ),
    .A2(_03280_),
    .B1(_03286_),
    .C1(_03277_),
    .X(_00858_));
 sky130_fd_sc_hd__or2_1 _19370_ (.A(\rbzero.spi_registers.texadd3[4] ),
    .B(_03282_),
    .X(_03287_));
 sky130_fd_sc_hd__o211a_1 _19371_ (.A1(\rbzero.spi_registers.new_texadd[3][4] ),
    .A2(_03280_),
    .B1(_03287_),
    .C1(_03277_),
    .X(_00859_));
 sky130_fd_sc_hd__or2_1 _19372_ (.A(\rbzero.spi_registers.texadd3[5] ),
    .B(_03282_),
    .X(_03288_));
 sky130_fd_sc_hd__o211a_1 _19373_ (.A1(\rbzero.spi_registers.new_texadd[3][5] ),
    .A2(_03280_),
    .B1(_03288_),
    .C1(_03277_),
    .X(_00860_));
 sky130_fd_sc_hd__or2_1 _19374_ (.A(\rbzero.spi_registers.texadd3[6] ),
    .B(_03282_),
    .X(_03289_));
 sky130_fd_sc_hd__o211a_1 _19375_ (.A1(\rbzero.spi_registers.new_texadd[3][6] ),
    .A2(_03280_),
    .B1(_03289_),
    .C1(_03277_),
    .X(_00861_));
 sky130_fd_sc_hd__or2_1 _19376_ (.A(\rbzero.spi_registers.texadd3[7] ),
    .B(_03282_),
    .X(_03290_));
 sky130_fd_sc_hd__o211a_1 _19377_ (.A1(\rbzero.spi_registers.new_texadd[3][7] ),
    .A2(_03280_),
    .B1(_03290_),
    .C1(_03277_),
    .X(_00862_));
 sky130_fd_sc_hd__or2_1 _19378_ (.A(\rbzero.spi_registers.texadd3[8] ),
    .B(_03282_),
    .X(_03291_));
 sky130_fd_sc_hd__clkbuf_4 _19379_ (.A(_09808_),
    .X(_03292_));
 sky130_fd_sc_hd__o211a_1 _19380_ (.A1(\rbzero.spi_registers.new_texadd[3][8] ),
    .A2(_03280_),
    .B1(_03291_),
    .C1(_03292_),
    .X(_00863_));
 sky130_fd_sc_hd__or2_1 _19381_ (.A(\rbzero.spi_registers.texadd3[9] ),
    .B(_03282_),
    .X(_03293_));
 sky130_fd_sc_hd__o211a_1 _19382_ (.A1(\rbzero.spi_registers.new_texadd[3][9] ),
    .A2(_03280_),
    .B1(_03293_),
    .C1(_03292_),
    .X(_00864_));
 sky130_fd_sc_hd__clkbuf_4 _19383_ (.A(_03279_),
    .X(_03294_));
 sky130_fd_sc_hd__buf_2 _19384_ (.A(_03281_),
    .X(_03295_));
 sky130_fd_sc_hd__or2_1 _19385_ (.A(\rbzero.spi_registers.texadd3[10] ),
    .B(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__o211a_1 _19386_ (.A1(\rbzero.spi_registers.new_texadd[3][10] ),
    .A2(_03294_),
    .B1(_03296_),
    .C1(_03292_),
    .X(_00865_));
 sky130_fd_sc_hd__or2_1 _19387_ (.A(\rbzero.spi_registers.texadd3[11] ),
    .B(_03295_),
    .X(_03297_));
 sky130_fd_sc_hd__o211a_1 _19388_ (.A1(\rbzero.spi_registers.new_texadd[3][11] ),
    .A2(_03294_),
    .B1(_03297_),
    .C1(_03292_),
    .X(_00866_));
 sky130_fd_sc_hd__or2_1 _19389_ (.A(\rbzero.spi_registers.texadd3[12] ),
    .B(_03295_),
    .X(_03298_));
 sky130_fd_sc_hd__o211a_1 _19390_ (.A1(\rbzero.spi_registers.new_texadd[3][12] ),
    .A2(_03294_),
    .B1(_03298_),
    .C1(_03292_),
    .X(_00867_));
 sky130_fd_sc_hd__or2_1 _19391_ (.A(\rbzero.spi_registers.texadd3[13] ),
    .B(_03295_),
    .X(_03299_));
 sky130_fd_sc_hd__o211a_1 _19392_ (.A1(\rbzero.spi_registers.new_texadd[3][13] ),
    .A2(_03294_),
    .B1(_03299_),
    .C1(_03292_),
    .X(_00868_));
 sky130_fd_sc_hd__or2_1 _19393_ (.A(\rbzero.spi_registers.texadd3[14] ),
    .B(_03295_),
    .X(_03300_));
 sky130_fd_sc_hd__o211a_1 _19394_ (.A1(\rbzero.spi_registers.new_texadd[3][14] ),
    .A2(_03294_),
    .B1(_03300_),
    .C1(_03292_),
    .X(_00869_));
 sky130_fd_sc_hd__or2_1 _19395_ (.A(\rbzero.spi_registers.texadd3[15] ),
    .B(_03295_),
    .X(_03301_));
 sky130_fd_sc_hd__o211a_1 _19396_ (.A1(\rbzero.spi_registers.new_texadd[3][15] ),
    .A2(_03294_),
    .B1(_03301_),
    .C1(_03292_),
    .X(_00870_));
 sky130_fd_sc_hd__or2_1 _19397_ (.A(\rbzero.spi_registers.texadd3[16] ),
    .B(_03295_),
    .X(_03302_));
 sky130_fd_sc_hd__o211a_1 _19398_ (.A1(\rbzero.spi_registers.new_texadd[3][16] ),
    .A2(_03294_),
    .B1(_03302_),
    .C1(_03292_),
    .X(_00871_));
 sky130_fd_sc_hd__or2_1 _19399_ (.A(\rbzero.spi_registers.texadd3[17] ),
    .B(_03295_),
    .X(_03303_));
 sky130_fd_sc_hd__o211a_1 _19400_ (.A1(\rbzero.spi_registers.new_texadd[3][17] ),
    .A2(_03294_),
    .B1(_03303_),
    .C1(_03292_),
    .X(_00872_));
 sky130_fd_sc_hd__or2_1 _19401_ (.A(\rbzero.spi_registers.texadd3[18] ),
    .B(_03295_),
    .X(_03304_));
 sky130_fd_sc_hd__buf_4 _19402_ (.A(_09808_),
    .X(_03305_));
 sky130_fd_sc_hd__o211a_1 _19403_ (.A1(\rbzero.spi_registers.new_texadd[3][18] ),
    .A2(_03294_),
    .B1(_03304_),
    .C1(_03305_),
    .X(_00873_));
 sky130_fd_sc_hd__or2_1 _19404_ (.A(\rbzero.spi_registers.texadd3[19] ),
    .B(_03295_),
    .X(_03306_));
 sky130_fd_sc_hd__o211a_1 _19405_ (.A1(\rbzero.spi_registers.new_texadd[3][19] ),
    .A2(_03294_),
    .B1(_03306_),
    .C1(_03305_),
    .X(_00874_));
 sky130_fd_sc_hd__or2_1 _19406_ (.A(\rbzero.spi_registers.texadd3[20] ),
    .B(_03281_),
    .X(_03307_));
 sky130_fd_sc_hd__o211a_1 _19407_ (.A1(\rbzero.spi_registers.new_texadd[3][20] ),
    .A2(_03279_),
    .B1(_03307_),
    .C1(_03305_),
    .X(_00875_));
 sky130_fd_sc_hd__or2_1 _19408_ (.A(\rbzero.spi_registers.texadd3[21] ),
    .B(_03281_),
    .X(_03308_));
 sky130_fd_sc_hd__o211a_1 _19409_ (.A1(\rbzero.spi_registers.new_texadd[3][21] ),
    .A2(_03279_),
    .B1(_03308_),
    .C1(_03305_),
    .X(_00876_));
 sky130_fd_sc_hd__or2_1 _19410_ (.A(\rbzero.spi_registers.texadd3[22] ),
    .B(_03281_),
    .X(_03309_));
 sky130_fd_sc_hd__o211a_1 _19411_ (.A1(\rbzero.spi_registers.new_texadd[3][22] ),
    .A2(_03279_),
    .B1(_03309_),
    .C1(_03305_),
    .X(_00877_));
 sky130_fd_sc_hd__or2_1 _19412_ (.A(\rbzero.spi_registers.texadd3[23] ),
    .B(_03281_),
    .X(_03310_));
 sky130_fd_sc_hd__o211a_1 _19413_ (.A1(\rbzero.spi_registers.new_texadd[3][23] ),
    .A2(_03279_),
    .B1(_03310_),
    .C1(_03305_),
    .X(_00878_));
 sky130_fd_sc_hd__and2_1 _19414_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_03157_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_2 _19415_ (.A(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__nand2_1 _19416_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_03157_),
    .Y(_03313_));
 sky130_fd_sc_hd__or2_1 _19417_ (.A(\rbzero.spi_registers.new_leak[0] ),
    .B(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__o211a_1 _19418_ (.A1(\rbzero.floor_leak[0] ),
    .A2(_03312_),
    .B1(_03314_),
    .C1(_03305_),
    .X(_00879_));
 sky130_fd_sc_hd__or2_1 _19419_ (.A(\rbzero.spi_registers.new_leak[1] ),
    .B(_03313_),
    .X(_03315_));
 sky130_fd_sc_hd__o211a_1 _19420_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_03312_),
    .B1(_03315_),
    .C1(_03305_),
    .X(_00880_));
 sky130_fd_sc_hd__or2_1 _19421_ (.A(\rbzero.spi_registers.new_leak[2] ),
    .B(_03313_),
    .X(_03316_));
 sky130_fd_sc_hd__o211a_1 _19422_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_03312_),
    .B1(_03316_),
    .C1(_03305_),
    .X(_00881_));
 sky130_fd_sc_hd__or2_1 _19423_ (.A(\rbzero.spi_registers.new_leak[3] ),
    .B(_03313_),
    .X(_03317_));
 sky130_fd_sc_hd__o211a_1 _19424_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_03312_),
    .B1(_03317_),
    .C1(_03305_),
    .X(_00882_));
 sky130_fd_sc_hd__or2_1 _19425_ (.A(\rbzero.spi_registers.new_leak[4] ),
    .B(_03313_),
    .X(_03318_));
 sky130_fd_sc_hd__buf_6 _19426_ (.A(_09808_),
    .X(_03319_));
 sky130_fd_sc_hd__o211a_1 _19427_ (.A1(\rbzero.floor_leak[4] ),
    .A2(_03312_),
    .B1(_03318_),
    .C1(_03319_),
    .X(_00883_));
 sky130_fd_sc_hd__or2_1 _19428_ (.A(\rbzero.spi_registers.new_leak[5] ),
    .B(_03313_),
    .X(_03320_));
 sky130_fd_sc_hd__o211a_1 _19429_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_03312_),
    .B1(_03320_),
    .C1(_03319_),
    .X(_00884_));
 sky130_fd_sc_hd__nand2_2 _19430_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_03140_),
    .Y(_03321_));
 sky130_fd_sc_hd__buf_6 _19431_ (.A(_04469_),
    .X(_03322_));
 sky130_fd_sc_hd__a31o_1 _19432_ (.A1(\rbzero.spi_registers.new_sky[0] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_03157_),
    .B1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__a21o_1 _19433_ (.A1(\rbzero.color_sky[0] ),
    .A2(_03321_),
    .B1(_03323_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _19434_ (.A0(\rbzero.spi_registers.new_sky[1] ),
    .A1(\rbzero.color_sky[1] ),
    .S(_03321_),
    .X(_03324_));
 sky130_fd_sc_hd__and2_1 _19435_ (.A(_08190_),
    .B(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _19436_ (.A(_03325_),
    .X(_00886_));
 sky130_fd_sc_hd__a31o_1 _19437_ (.A1(\rbzero.spi_registers.new_sky[2] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_03157_),
    .B1(_03322_),
    .X(_03326_));
 sky130_fd_sc_hd__a21o_1 _19438_ (.A1(\rbzero.color_sky[2] ),
    .A2(_03321_),
    .B1(_03326_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _19439_ (.A0(\rbzero.spi_registers.new_sky[3] ),
    .A1(\rbzero.color_sky[3] ),
    .S(_03321_),
    .X(_03327_));
 sky130_fd_sc_hd__and2_1 _19440_ (.A(_08190_),
    .B(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__clkbuf_1 _19441_ (.A(_03328_),
    .X(_00888_));
 sky130_fd_sc_hd__a31o_1 _19442_ (.A1(\rbzero.spi_registers.new_sky[4] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_03157_),
    .B1(_03322_),
    .X(_03329_));
 sky130_fd_sc_hd__a21o_1 _19443_ (.A1(\rbzero.color_sky[4] ),
    .A2(_03321_),
    .B1(_03329_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _19444_ (.A0(\rbzero.spi_registers.new_sky[5] ),
    .A1(\rbzero.color_sky[5] ),
    .S(_03321_),
    .X(_03330_));
 sky130_fd_sc_hd__and2_1 _19445_ (.A(_08190_),
    .B(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _19446_ (.A(_03331_),
    .X(_00890_));
 sky130_fd_sc_hd__nand2_2 _19447_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_03140_),
    .Y(_03332_));
 sky130_fd_sc_hd__mux2_1 _19448_ (.A0(\rbzero.spi_registers.new_floor[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__and2_1 _19449_ (.A(_08190_),
    .B(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__clkbuf_1 _19450_ (.A(_03334_),
    .X(_00891_));
 sky130_fd_sc_hd__a31o_1 _19451_ (.A1(\rbzero.spi_registers.new_floor[1] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_03157_),
    .B1(_03322_),
    .X(_03335_));
 sky130_fd_sc_hd__a21o_1 _19452_ (.A1(\rbzero.color_floor[1] ),
    .A2(_03332_),
    .B1(_03335_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _19453_ (.A0(\rbzero.spi_registers.new_floor[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_03332_),
    .X(_03336_));
 sky130_fd_sc_hd__and2_1 _19454_ (.A(_08190_),
    .B(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_1 _19455_ (.A(_03337_),
    .X(_00893_));
 sky130_fd_sc_hd__a31o_1 _19456_ (.A1(\rbzero.spi_registers.new_floor[3] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_03157_),
    .B1(_03322_),
    .X(_03338_));
 sky130_fd_sc_hd__a21o_1 _19457_ (.A1(\rbzero.color_floor[3] ),
    .A2(_03332_),
    .B1(_03338_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _19458_ (.A0(\rbzero.spi_registers.new_floor[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_03332_),
    .X(_03339_));
 sky130_fd_sc_hd__and2_1 _19459_ (.A(_08190_),
    .B(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__clkbuf_1 _19460_ (.A(_03340_),
    .X(_00895_));
 sky130_fd_sc_hd__a31o_1 _19461_ (.A1(\rbzero.spi_registers.new_floor[5] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_03157_),
    .B1(_03322_),
    .X(_03341_));
 sky130_fd_sc_hd__a21o_1 _19462_ (.A1(\rbzero.color_floor[5] ),
    .A2(_03332_),
    .B1(_03341_),
    .X(_00896_));
 sky130_fd_sc_hd__and2_1 _19463_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_03140_),
    .X(_03342_));
 sky130_fd_sc_hd__clkbuf_2 _19464_ (.A(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__nand2_1 _19465_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_03157_),
    .Y(_03344_));
 sky130_fd_sc_hd__or2_1 _19466_ (.A(\rbzero.spi_registers.new_vshift[0] ),
    .B(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__o211a_1 _19467_ (.A1(\rbzero.spi_registers.vshift[0] ),
    .A2(_03343_),
    .B1(_03345_),
    .C1(_03319_),
    .X(_00897_));
 sky130_fd_sc_hd__or2_1 _19468_ (.A(\rbzero.spi_registers.new_vshift[1] ),
    .B(_03344_),
    .X(_03346_));
 sky130_fd_sc_hd__o211a_1 _19469_ (.A1(\rbzero.spi_registers.vshift[1] ),
    .A2(_03343_),
    .B1(_03346_),
    .C1(_03319_),
    .X(_00898_));
 sky130_fd_sc_hd__or2_1 _19470_ (.A(\rbzero.spi_registers.new_vshift[2] ),
    .B(_03344_),
    .X(_03347_));
 sky130_fd_sc_hd__o211a_1 _19471_ (.A1(\rbzero.spi_registers.vshift[2] ),
    .A2(_03343_),
    .B1(_03347_),
    .C1(_03319_),
    .X(_00899_));
 sky130_fd_sc_hd__or2_1 _19472_ (.A(\rbzero.spi_registers.new_vshift[3] ),
    .B(_03344_),
    .X(_03348_));
 sky130_fd_sc_hd__o211a_1 _19473_ (.A1(\rbzero.spi_registers.vshift[3] ),
    .A2(_03343_),
    .B1(_03348_),
    .C1(_03319_),
    .X(_00900_));
 sky130_fd_sc_hd__or2_1 _19474_ (.A(\rbzero.spi_registers.new_vshift[4] ),
    .B(_03344_),
    .X(_03349_));
 sky130_fd_sc_hd__o211a_1 _19475_ (.A1(\rbzero.spi_registers.vshift[4] ),
    .A2(_03343_),
    .B1(_03349_),
    .C1(_03319_),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _19476_ (.A(\rbzero.spi_registers.new_vshift[5] ),
    .B(_03344_),
    .X(_03350_));
 sky130_fd_sc_hd__o211a_1 _19477_ (.A1(\rbzero.spi_registers.vshift[5] ),
    .A2(_03343_),
    .B1(_03350_),
    .C1(_03319_),
    .X(_00902_));
 sky130_fd_sc_hd__and4b_1 _19478_ (.A_N(\rbzero.spi_registers.spi_done ),
    .B(_02989_),
    .C(_02966_),
    .D(_02988_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_1 _19479_ (.A(_03351_),
    .X(_00903_));
 sky130_fd_sc_hd__or3b_1 _19480_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .B(\rbzero.spi_registers.spi_cmd[3] ),
    .C_N(\rbzero.spi_registers.spi_done ),
    .X(_03352_));
 sky130_fd_sc_hd__or3_1 _19481_ (.A(_04469_),
    .B(_02967_),
    .C(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__buf_2 _19482_ (.A(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _19483_ (.A0(_02502_),
    .A1(\rbzero.spi_registers.new_sky[0] ),
    .S(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__clkbuf_1 _19484_ (.A(_03355_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _19485_ (.A0(_02509_),
    .A1(\rbzero.spi_registers.new_sky[1] ),
    .S(_03354_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _19486_ (.A(_03356_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _19487_ (.A0(_02511_),
    .A1(\rbzero.spi_registers.new_sky[2] ),
    .S(_03354_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _19488_ (.A(_03357_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _19489_ (.A0(_02513_),
    .A1(\rbzero.spi_registers.new_sky[3] ),
    .S(_03354_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_1 _19490_ (.A(_03358_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _19491_ (.A0(_02515_),
    .A1(\rbzero.spi_registers.new_sky[4] ),
    .S(_03354_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_1 _19492_ (.A(_03359_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _19493_ (.A0(_02517_),
    .A1(\rbzero.spi_registers.new_sky[5] ),
    .S(_03354_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_1 _19494_ (.A(_03360_),
    .X(_00909_));
 sky130_fd_sc_hd__buf_4 _19495_ (.A(_03156_),
    .X(_03361_));
 sky130_fd_sc_hd__inv_2 _19496_ (.A(_03354_),
    .Y(_03362_));
 sky130_fd_sc_hd__a31o_1 _19497_ (.A1(\rbzero.spi_registers.got_new_sky ),
    .A2(_03159_),
    .A3(_03361_),
    .B1(_03362_),
    .X(_00910_));
 sky130_fd_sc_hd__or4b_2 _19498_ (.A(_02503_),
    .B(_04468_),
    .C(_03352_),
    .D_N(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_03363_));
 sky130_fd_sc_hd__buf_2 _19499_ (.A(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_1 _19500_ (.A0(_02502_),
    .A1(\rbzero.spi_registers.new_floor[0] ),
    .S(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_1 _19501_ (.A(_03365_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _19502_ (.A0(_02509_),
    .A1(\rbzero.spi_registers.new_floor[1] ),
    .S(_03364_),
    .X(_03366_));
 sky130_fd_sc_hd__clkbuf_1 _19503_ (.A(_03366_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _19504_ (.A0(_02511_),
    .A1(\rbzero.spi_registers.new_floor[2] ),
    .S(_03364_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_1 _19505_ (.A(_03367_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _19506_ (.A0(_02513_),
    .A1(\rbzero.spi_registers.new_floor[3] ),
    .S(_03364_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_1 _19507_ (.A(_03368_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _19508_ (.A0(_02515_),
    .A1(\rbzero.spi_registers.new_floor[4] ),
    .S(_03364_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_1 _19509_ (.A(_03369_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _19510_ (.A0(_02517_),
    .A1(\rbzero.spi_registers.new_floor[5] ),
    .S(_03364_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _19511_ (.A(_03370_),
    .X(_00916_));
 sky130_fd_sc_hd__inv_2 _19512_ (.A(_03364_),
    .Y(_03371_));
 sky130_fd_sc_hd__a31o_1 _19513_ (.A1(\rbzero.spi_registers.got_new_floor ),
    .A2(_03159_),
    .A3(_03361_),
    .B1(_03371_),
    .X(_00917_));
 sky130_fd_sc_hd__or2b_1 _19514_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B_N(_02503_),
    .X(_03372_));
 sky130_fd_sc_hd__or3_2 _19515_ (.A(_04468_),
    .B(_03352_),
    .C(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__buf_2 _19516_ (.A(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _19517_ (.A0(_02502_),
    .A1(\rbzero.spi_registers.new_leak[0] ),
    .S(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _19518_ (.A(_03375_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _19519_ (.A0(_02509_),
    .A1(\rbzero.spi_registers.new_leak[1] ),
    .S(_03374_),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_1 _19520_ (.A(_03376_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _19521_ (.A0(_02511_),
    .A1(\rbzero.spi_registers.new_leak[2] ),
    .S(_03374_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_1 _19522_ (.A(_03377_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _19523_ (.A0(_02513_),
    .A1(\rbzero.spi_registers.new_leak[3] ),
    .S(_03374_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _19524_ (.A(_03378_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _19525_ (.A0(_02515_),
    .A1(\rbzero.spi_registers.new_leak[4] ),
    .S(_03374_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_1 _19526_ (.A(_03379_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _19527_ (.A0(_02517_),
    .A1(\rbzero.spi_registers.new_leak[5] ),
    .S(_03374_),
    .X(_03380_));
 sky130_fd_sc_hd__clkbuf_1 _19528_ (.A(_03380_),
    .X(_00923_));
 sky130_fd_sc_hd__inv_2 _19529_ (.A(_03374_),
    .Y(_03381_));
 sky130_fd_sc_hd__a31o_1 _19530_ (.A1(\rbzero.spi_registers.got_new_leak ),
    .A2(_03159_),
    .A3(_03361_),
    .B1(_03381_),
    .X(_00924_));
 sky130_fd_sc_hd__or3_1 _19531_ (.A(_04468_),
    .B(_02970_),
    .C(_03352_),
    .X(_03382_));
 sky130_fd_sc_hd__clkbuf_4 _19532_ (.A(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__mux2_1 _19533_ (.A0(_02502_),
    .A1(\rbzero.spi_registers.new_other[0] ),
    .S(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__clkbuf_1 _19534_ (.A(_03384_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _19535_ (.A0(_02509_),
    .A1(\rbzero.spi_registers.new_other[1] ),
    .S(_03383_),
    .X(_03385_));
 sky130_fd_sc_hd__clkbuf_1 _19536_ (.A(_03385_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _19537_ (.A0(_02511_),
    .A1(\rbzero.spi_registers.new_other[2] ),
    .S(_03383_),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_1 _19538_ (.A(_03386_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19539_ (.A0(_02513_),
    .A1(\rbzero.spi_registers.new_other[3] ),
    .S(_03383_),
    .X(_03387_));
 sky130_fd_sc_hd__clkbuf_1 _19540_ (.A(_03387_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _19541_ (.A0(_02515_),
    .A1(\rbzero.spi_registers.new_other[4] ),
    .S(_03383_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_1 _19542_ (.A(_03388_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19543_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(\rbzero.spi_registers.new_other[6] ),
    .S(_03383_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_1 _19544_ (.A(_03389_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _19545_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.new_other[7] ),
    .S(_03383_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _19546_ (.A(_03390_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _19547_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.new_other[8] ),
    .S(_03383_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _19548_ (.A(_03391_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _19549_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.new_other[9] ),
    .S(_03383_),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_1 _19550_ (.A(_03392_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _19551_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.new_other[10] ),
    .S(_03382_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _19552_ (.A(_03393_),
    .X(_00934_));
 sky130_fd_sc_hd__inv_2 _19553_ (.A(_03383_),
    .Y(_03394_));
 sky130_fd_sc_hd__a31o_1 _19554_ (.A1(\rbzero.spi_registers.got_new_other ),
    .A2(_03159_),
    .A3(_03361_),
    .B1(_03394_),
    .X(_00935_));
 sky130_fd_sc_hd__and3_1 _19555_ (.A(\rbzero.spi_registers.spi_done ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .C(_02504_),
    .X(_03395_));
 sky130_fd_sc_hd__nor3b_4 _19556_ (.A(_04469_),
    .B(_02967_),
    .C_N(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__mux2_1 _19557_ (.A0(\rbzero.spi_registers.new_vshift[0] ),
    .A1(_02502_),
    .S(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_1 _19558_ (.A(_03397_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _19559_ (.A0(\rbzero.spi_registers.new_vshift[1] ),
    .A1(_02509_),
    .S(_03396_),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_1 _19560_ (.A(_03398_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _19561_ (.A0(\rbzero.spi_registers.new_vshift[2] ),
    .A1(_02511_),
    .S(_03396_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _19562_ (.A(_03399_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _19563_ (.A0(\rbzero.spi_registers.new_vshift[3] ),
    .A1(_02513_),
    .S(_03396_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_1 _19564_ (.A(_03400_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _19565_ (.A0(\rbzero.spi_registers.new_vshift[4] ),
    .A1(_02515_),
    .S(_03396_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_1 _19566_ (.A(_03401_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _19567_ (.A0(\rbzero.spi_registers.new_vshift[5] ),
    .A1(_02517_),
    .S(_03396_),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_1 _19568_ (.A(_03402_),
    .X(_00941_));
 sky130_fd_sc_hd__a31o_1 _19569_ (.A1(\rbzero.spi_registers.got_new_vshift ),
    .A2(_03159_),
    .A3(_03361_),
    .B1(_03396_),
    .X(_00942_));
 sky130_fd_sc_hd__and4b_1 _19570_ (.A_N(_02503_),
    .B(_04112_),
    .C(_03395_),
    .D(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _19571_ (.A0(\rbzero.spi_registers.new_vinf ),
    .A1(_02502_),
    .S(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _19572_ (.A(_03404_),
    .X(_00943_));
 sky130_fd_sc_hd__a31o_1 _19573_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_08186_),
    .A3(_03361_),
    .B1(_03403_),
    .X(_00944_));
 sky130_fd_sc_hd__and4b_1 _19574_ (.A_N(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02503_),
    .C(_04036_),
    .D(_03395_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_4 _19575_ (.A(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_4 _19576_ (.A(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__mux2_1 _19577_ (.A0(\rbzero.spi_registers.new_mapd[0] ),
    .A1(_02502_),
    .S(_03407_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _19578_ (.A(_03408_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _19579_ (.A0(\rbzero.spi_registers.new_mapd[1] ),
    .A1(_02509_),
    .S(_03407_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _19580_ (.A(_03409_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _19581_ (.A0(\rbzero.spi_registers.new_mapd[2] ),
    .A1(_02511_),
    .S(_03407_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _19582_ (.A(_03410_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _19583_ (.A0(\rbzero.spi_registers.new_mapd[3] ),
    .A1(_02513_),
    .S(_03407_),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _19584_ (.A(_03411_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _19585_ (.A0(\rbzero.spi_registers.new_mapd[4] ),
    .A1(_02515_),
    .S(_03407_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _19586_ (.A(_03412_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _19587_ (.A0(\rbzero.spi_registers.new_mapd[5] ),
    .A1(_02517_),
    .S(_03407_),
    .X(_03413_));
 sky130_fd_sc_hd__clkbuf_1 _19588_ (.A(_03413_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _19589_ (.A0(\rbzero.spi_registers.new_mapd[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03407_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _19590_ (.A(_03414_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _19591_ (.A0(\rbzero.spi_registers.new_mapd[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03407_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _19592_ (.A(_03415_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _19593_ (.A0(\rbzero.spi_registers.new_mapd[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03407_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _19594_ (.A(_03416_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _19595_ (.A0(\rbzero.spi_registers.new_mapd[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03406_),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _19596_ (.A(_03417_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _19597_ (.A0(\rbzero.spi_registers.new_mapd[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03406_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _19598_ (.A(_03418_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _19599_ (.A0(\rbzero.spi_registers.new_mapd[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03406_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _19600_ (.A(_03419_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _19601_ (.A0(\rbzero.spi_registers.new_mapd[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03406_),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_1 _19602_ (.A(_03420_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _19603_ (.A0(\rbzero.spi_registers.new_mapd[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03406_),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _19604_ (.A(_03421_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _19605_ (.A0(\rbzero.spi_registers.new_mapd[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03406_),
    .X(_03422_));
 sky130_fd_sc_hd__clkbuf_1 _19606_ (.A(_03422_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _19607_ (.A0(\rbzero.spi_registers.new_mapd[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03406_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_1 _19608_ (.A(_03423_),
    .X(_00960_));
 sky130_fd_sc_hd__a31o_1 _19609_ (.A1(\rbzero.spi_registers.got_new_mapd ),
    .A2(_08186_),
    .A3(_03361_),
    .B1(_03407_),
    .X(_00961_));
 sky130_fd_sc_hd__and3_1 _19610_ (.A(_04112_),
    .B(_02985_),
    .C(_03395_),
    .X(_03424_));
 sky130_fd_sc_hd__buf_4 _19611_ (.A(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__clkbuf_4 _19612_ (.A(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__a31o_1 _19613_ (.A1(\rbzero.spi_registers.got_new_texadd[0] ),
    .A2(_08186_),
    .A3(_03361_),
    .B1(_03426_),
    .X(_00962_));
 sky130_fd_sc_hd__nor2_4 _19614_ (.A(_02505_),
    .B(_02967_),
    .Y(_03427_));
 sky130_fd_sc_hd__buf_4 _19615_ (.A(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__a31o_1 _19616_ (.A1(\rbzero.spi_registers.got_new_texadd[1] ),
    .A2(_08186_),
    .A3(_03361_),
    .B1(_03428_),
    .X(_00963_));
 sky130_fd_sc_hd__a31o_1 _19617_ (.A1(\rbzero.spi_registers.got_new_texadd[2] ),
    .A2(_08186_),
    .A3(_03361_),
    .B1(_02507_),
    .X(_00964_));
 sky130_fd_sc_hd__nor2_4 _19618_ (.A(_02505_),
    .B(_03372_),
    .Y(_03429_));
 sky130_fd_sc_hd__buf_4 _19619_ (.A(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__a31o_1 _19620_ (.A1(\rbzero.spi_registers.got_new_texadd[3] ),
    .A2(_08186_),
    .A3(_03156_),
    .B1(_03430_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _19621_ (.A0(\rbzero.spi_registers.new_texadd[0][0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03426_),
    .X(_03431_));
 sky130_fd_sc_hd__clkbuf_1 _19622_ (.A(_03431_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _19623_ (.A0(\rbzero.spi_registers.new_texadd[0][1] ),
    .A1(_02509_),
    .S(_03426_),
    .X(_03432_));
 sky130_fd_sc_hd__clkbuf_1 _19624_ (.A(_03432_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _19625_ (.A0(\rbzero.spi_registers.new_texadd[0][2] ),
    .A1(_02511_),
    .S(_03426_),
    .X(_03433_));
 sky130_fd_sc_hd__clkbuf_1 _19626_ (.A(_03433_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _19627_ (.A0(\rbzero.spi_registers.new_texadd[0][3] ),
    .A1(_02513_),
    .S(_03426_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_1 _19628_ (.A(_03434_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _19629_ (.A0(\rbzero.spi_registers.new_texadd[0][4] ),
    .A1(_02515_),
    .S(_03426_),
    .X(_03435_));
 sky130_fd_sc_hd__clkbuf_1 _19630_ (.A(_03435_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _19631_ (.A0(\rbzero.spi_registers.new_texadd[0][5] ),
    .A1(_02517_),
    .S(_03426_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_1 _19632_ (.A(_03436_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _19633_ (.A0(\rbzero.spi_registers.new_texadd[0][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03426_),
    .X(_03437_));
 sky130_fd_sc_hd__clkbuf_1 _19634_ (.A(_03437_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _19635_ (.A0(\rbzero.spi_registers.new_texadd[0][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03426_),
    .X(_03438_));
 sky130_fd_sc_hd__clkbuf_1 _19636_ (.A(_03438_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _19637_ (.A0(\rbzero.spi_registers.new_texadd[0][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03426_),
    .X(_03439_));
 sky130_fd_sc_hd__clkbuf_1 _19638_ (.A(_03439_),
    .X(_00974_));
 sky130_fd_sc_hd__buf_4 _19639_ (.A(_03425_),
    .X(_03440_));
 sky130_fd_sc_hd__mux2_1 _19640_ (.A0(\rbzero.spi_registers.new_texadd[0][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_1 _19641_ (.A(_03441_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _19642_ (.A0(\rbzero.spi_registers.new_texadd[0][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03440_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_1 _19643_ (.A(_03442_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _19644_ (.A0(\rbzero.spi_registers.new_texadd[0][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03440_),
    .X(_03443_));
 sky130_fd_sc_hd__clkbuf_1 _19645_ (.A(_03443_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _19646_ (.A0(\rbzero.spi_registers.new_texadd[0][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03440_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_1 _19647_ (.A(_03444_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _19648_ (.A0(\rbzero.spi_registers.new_texadd[0][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03440_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_1 _19649_ (.A(_03445_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _19650_ (.A0(\rbzero.spi_registers.new_texadd[0][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03440_),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_1 _19651_ (.A(_03446_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _19652_ (.A0(\rbzero.spi_registers.new_texadd[0][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03440_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _19653_ (.A(_03447_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _19654_ (.A0(\rbzero.spi_registers.new_texadd[0][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03440_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_1 _19655_ (.A(_03448_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _19656_ (.A0(\rbzero.spi_registers.new_texadd[0][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03440_),
    .X(_03449_));
 sky130_fd_sc_hd__clkbuf_1 _19657_ (.A(_03449_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _19658_ (.A0(\rbzero.spi_registers.new_texadd[0][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03440_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_1 _19659_ (.A(_03450_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _19660_ (.A0(\rbzero.spi_registers.new_texadd[0][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03425_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_1 _19661_ (.A(_03451_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _19662_ (.A0(\rbzero.spi_registers.new_texadd[0][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03425_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_1 _19663_ (.A(_03452_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _19664_ (.A0(\rbzero.spi_registers.new_texadd[0][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03425_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _19665_ (.A(_03453_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _19666_ (.A0(\rbzero.spi_registers.new_texadd[0][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03425_),
    .X(_03454_));
 sky130_fd_sc_hd__clkbuf_1 _19667_ (.A(_03454_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _19668_ (.A0(\rbzero.spi_registers.new_texadd[0][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03425_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_1 _19669_ (.A(_03455_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _19670_ (.A0(\rbzero.spi_registers.new_texadd[1][0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03428_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_1 _19671_ (.A(_03456_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _19672_ (.A0(\rbzero.spi_registers.new_texadd[1][1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_03428_),
    .X(_03457_));
 sky130_fd_sc_hd__clkbuf_1 _19673_ (.A(_03457_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _19674_ (.A0(\rbzero.spi_registers.new_texadd[1][2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_03428_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_1 _19675_ (.A(_03458_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _19676_ (.A0(\rbzero.spi_registers.new_texadd[1][3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_03428_),
    .X(_03459_));
 sky130_fd_sc_hd__clkbuf_1 _19677_ (.A(_03459_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _19678_ (.A0(\rbzero.spi_registers.new_texadd[1][4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_03428_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _19679_ (.A(_03460_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _19680_ (.A0(\rbzero.spi_registers.new_texadd[1][5] ),
    .A1(_02517_),
    .S(_03428_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_1 _19681_ (.A(_03461_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _19682_ (.A0(\rbzero.spi_registers.new_texadd[1][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03428_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_1 _19683_ (.A(_03462_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _19684_ (.A0(\rbzero.spi_registers.new_texadd[1][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03428_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_1 _19685_ (.A(_03463_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _19686_ (.A0(\rbzero.spi_registers.new_texadd[1][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03428_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_1 _19687_ (.A(_03464_),
    .X(_00998_));
 sky130_fd_sc_hd__buf_4 _19688_ (.A(_03427_),
    .X(_03465_));
 sky130_fd_sc_hd__mux2_1 _19689_ (.A0(\rbzero.spi_registers.new_texadd[1][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _19690_ (.A(_03466_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _19691_ (.A0(\rbzero.spi_registers.new_texadd[1][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03465_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_1 _19692_ (.A(_03467_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _19693_ (.A0(\rbzero.spi_registers.new_texadd[1][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03465_),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_1 _19694_ (.A(_03468_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _19695_ (.A0(\rbzero.spi_registers.new_texadd[1][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03465_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _19696_ (.A(_03469_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _19697_ (.A0(\rbzero.spi_registers.new_texadd[1][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03465_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_1 _19698_ (.A(_03470_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _19699_ (.A0(\rbzero.spi_registers.new_texadd[1][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03465_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_1 _19700_ (.A(_03471_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _19701_ (.A0(\rbzero.spi_registers.new_texadd[1][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03465_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _19702_ (.A(_03472_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _19703_ (.A0(\rbzero.spi_registers.new_texadd[1][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03465_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_1 _19704_ (.A(_03473_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _19705_ (.A0(\rbzero.spi_registers.new_texadd[1][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03465_),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_1 _19706_ (.A(_03474_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _19707_ (.A0(\rbzero.spi_registers.new_texadd[1][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03465_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _19708_ (.A(_03475_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _19709_ (.A0(\rbzero.spi_registers.new_texadd[1][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03427_),
    .X(_03476_));
 sky130_fd_sc_hd__clkbuf_1 _19710_ (.A(_03476_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _19711_ (.A0(\rbzero.spi_registers.new_texadd[1][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03427_),
    .X(_03477_));
 sky130_fd_sc_hd__clkbuf_1 _19712_ (.A(_03477_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _19713_ (.A0(\rbzero.spi_registers.new_texadd[1][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03427_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_1 _19714_ (.A(_03478_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _19715_ (.A0(\rbzero.spi_registers.new_texadd[1][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03427_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_1 _19716_ (.A(_03479_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _19717_ (.A0(\rbzero.spi_registers.new_texadd[1][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03427_),
    .X(_03480_));
 sky130_fd_sc_hd__clkbuf_1 _19718_ (.A(_03480_),
    .X(_01013_));
 sky130_fd_sc_hd__nor2_2 _19719_ (.A(net41),
    .B(net40),
    .Y(_03481_));
 sky130_fd_sc_hd__or2_1 _19720_ (.A(_03156_),
    .B(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_4 _19721_ (.A(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__clkbuf_4 _19722_ (.A(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__o211a_1 _19723_ (.A1(\rbzero.pov.spi_done ),
    .A2(\rbzero.pov.ready ),
    .B1(_03159_),
    .C1(_03484_),
    .X(_01014_));
 sky130_fd_sc_hd__nor2b_2 _19724_ (.A(\rbzero.pov.sclk_buffer[2] ),
    .B_N(\rbzero.pov.sclk_buffer[1] ),
    .Y(_03485_));
 sky130_fd_sc_hd__nor2_2 _19725_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(_04468_),
    .Y(_03486_));
 sky130_fd_sc_hd__o21ai_1 _19726_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03485_),
    .B1(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__a21oi_1 _19727_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03485_),
    .B1(_03487_),
    .Y(_01015_));
 sky130_fd_sc_hd__and3_1 _19728_ (.A(\rbzero.pov.spi_counter[1] ),
    .B(\rbzero.pov.spi_counter[0] ),
    .C(_03485_),
    .X(_03488_));
 sky130_fd_sc_hd__a21o_1 _19729_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03485_),
    .B1(\rbzero.pov.spi_counter[1] ),
    .X(_03489_));
 sky130_fd_sc_hd__and4bb_1 _19730_ (.A_N(\rbzero.pov.spi_counter[5] ),
    .B_N(\rbzero.pov.spi_counter[4] ),
    .C(\rbzero.pov.spi_counter[3] ),
    .D(\rbzero.pov.spi_counter[6] ),
    .X(_03490_));
 sky130_fd_sc_hd__and4bb_1 _19731_ (.A_N(\rbzero.pov.spi_counter[2] ),
    .B_N(\rbzero.pov.spi_counter[1] ),
    .C(\rbzero.pov.spi_counter[0] ),
    .D(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__a21boi_1 _19732_ (.A1(_03485_),
    .A2(_03491_),
    .B1_N(_03486_),
    .Y(_03492_));
 sky130_fd_sc_hd__and3b_1 _19733_ (.A_N(_03488_),
    .B(_03489_),
    .C(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__clkbuf_1 _19734_ (.A(_03493_),
    .X(_01016_));
 sky130_fd_sc_hd__and2_1 _19735_ (.A(\rbzero.pov.spi_counter[2] ),
    .B(_03488_),
    .X(_03494_));
 sky130_fd_sc_hd__o21ai_1 _19736_ (.A1(\rbzero.pov.spi_counter[2] ),
    .A2(_03488_),
    .B1(_03486_),
    .Y(_03495_));
 sky130_fd_sc_hd__nor2_1 _19737_ (.A(_03494_),
    .B(_03495_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _19738_ (.A(\rbzero.pov.spi_counter[3] ),
    .B(_03494_),
    .Y(_03496_));
 sky130_fd_sc_hd__o211a_1 _19739_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_03494_),
    .B1(_03496_),
    .C1(_03492_),
    .X(_01018_));
 sky130_fd_sc_hd__and3_1 _19740_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[3] ),
    .C(_03494_),
    .X(_03497_));
 sky130_fd_sc_hd__a31o_1 _19741_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(\rbzero.pov.spi_counter[2] ),
    .A3(_03488_),
    .B1(\rbzero.pov.spi_counter[4] ),
    .X(_03498_));
 sky130_fd_sc_hd__and3b_1 _19742_ (.A_N(_03497_),
    .B(_03486_),
    .C(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_1 _19743_ (.A(_03499_),
    .X(_01019_));
 sky130_fd_sc_hd__and2_1 _19744_ (.A(\rbzero.pov.spi_counter[5] ),
    .B(_03497_),
    .X(_03500_));
 sky130_fd_sc_hd__o21ai_1 _19745_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_03497_),
    .B1(_03486_),
    .Y(_03501_));
 sky130_fd_sc_hd__nor2_1 _19746_ (.A(_03500_),
    .B(_03501_),
    .Y(_01020_));
 sky130_fd_sc_hd__a21boi_1 _19747_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03500_),
    .B1_N(_03492_),
    .Y(_03502_));
 sky130_fd_sc_hd__o21a_1 _19748_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03500_),
    .B1(_03502_),
    .X(_01021_));
 sky130_fd_sc_hd__buf_1 _19749_ (.A(clknet_1_1__leaf__05825_),
    .X(_03503_));
 sky130_fd_sc_hd__buf_1 _19750_ (.A(clknet_1_1__leaf__03503_),
    .X(_03504_));
 sky130_fd_sc_hd__inv_2 _19752__29 (.A(clknet_1_0__leaf__03504_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _19753__30 (.A(clknet_1_0__leaf__03504_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _19754__31 (.A(clknet_1_1__leaf__03504_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _19755__32 (.A(clknet_1_1__leaf__03504_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _19756__33 (.A(clknet_1_1__leaf__03504_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _19757__34 (.A(clknet_1_1__leaf__03504_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _19758__35 (.A(clknet_1_1__leaf__03504_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _19759__36 (.A(clknet_1_1__leaf__03504_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _19760__37 (.A(clknet_1_0__leaf__03504_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _19762__38 (.A(clknet_1_1__leaf__03505_),
    .Y(net163));
 sky130_fd_sc_hd__buf_1 _19761_ (.A(clknet_1_1__leaf__03503_),
    .X(_03505_));
 sky130_fd_sc_hd__inv_2 _19763__39 (.A(clknet_1_1__leaf__03505_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _19764__40 (.A(clknet_1_1__leaf__03505_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _19765__41 (.A(clknet_1_1__leaf__03505_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _19766__42 (.A(clknet_1_1__leaf__03505_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _19767__43 (.A(clknet_1_1__leaf__03505_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _19768__44 (.A(clknet_1_0__leaf__03505_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _19769__45 (.A(clknet_1_0__leaf__03505_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _19770__46 (.A(clknet_1_0__leaf__03505_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _19771__47 (.A(clknet_1_0__leaf__03505_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _19773__48 (.A(clknet_1_1__leaf__03506_),
    .Y(net173));
 sky130_fd_sc_hd__buf_1 _19772_ (.A(clknet_1_0__leaf__03503_),
    .X(_03506_));
 sky130_fd_sc_hd__inv_2 _19774__49 (.A(clknet_1_1__leaf__03506_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _19775__50 (.A(clknet_1_1__leaf__03506_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _19776__51 (.A(clknet_1_1__leaf__03506_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _19777__52 (.A(clknet_1_1__leaf__03506_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _19778__53 (.A(clknet_1_0__leaf__03506_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _19779__54 (.A(clknet_1_0__leaf__03506_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _19780__55 (.A(clknet_1_0__leaf__03506_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _19781__56 (.A(clknet_1_0__leaf__03506_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _19782__57 (.A(clknet_1_0__leaf__03506_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _19784__58 (.A(clknet_1_0__leaf__03507_),
    .Y(net183));
 sky130_fd_sc_hd__buf_1 _19783_ (.A(clknet_1_0__leaf__03503_),
    .X(_03507_));
 sky130_fd_sc_hd__inv_2 _19785__59 (.A(clknet_1_0__leaf__03507_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _19786__60 (.A(clknet_1_0__leaf__03507_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _19787__61 (.A(clknet_1_0__leaf__03507_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _19788__62 (.A(clknet_1_0__leaf__03507_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _19789__63 (.A(clknet_1_1__leaf__03507_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _19790__64 (.A(clknet_1_1__leaf__03507_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _19791__65 (.A(clknet_1_1__leaf__03507_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _19792__66 (.A(clknet_1_1__leaf__03507_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _19793__67 (.A(clknet_1_1__leaf__03507_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _19795__68 (.A(clknet_1_0__leaf__03508_),
    .Y(net193));
 sky130_fd_sc_hd__buf_1 _19794_ (.A(clknet_1_1__leaf__03503_),
    .X(_03508_));
 sky130_fd_sc_hd__inv_2 _19796__69 (.A(clknet_1_0__leaf__03508_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _19797__70 (.A(clknet_1_0__leaf__03508_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _19798__71 (.A(clknet_1_0__leaf__03508_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _19799__72 (.A(clknet_1_0__leaf__03508_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _19800__73 (.A(clknet_1_1__leaf__03508_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _19801__74 (.A(clknet_1_1__leaf__03508_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _19802__75 (.A(clknet_1_1__leaf__03508_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _19803__76 (.A(clknet_1_1__leaf__03508_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _19804__77 (.A(clknet_1_1__leaf__03508_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _19806__78 (.A(clknet_1_0__leaf__03509_),
    .Y(net203));
 sky130_fd_sc_hd__buf_1 _19805_ (.A(clknet_1_1__leaf__03503_),
    .X(_03509_));
 sky130_fd_sc_hd__inv_2 _19807__79 (.A(clknet_1_0__leaf__03509_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _19808__80 (.A(clknet_1_0__leaf__03509_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _19809__81 (.A(clknet_1_0__leaf__03509_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _19810__82 (.A(clknet_1_0__leaf__03509_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _19811__83 (.A(clknet_1_1__leaf__03509_),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _19812__84 (.A(clknet_1_1__leaf__03509_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _19813__85 (.A(clknet_1_1__leaf__03509_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _19814__86 (.A(clknet_1_1__leaf__03509_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _19815__87 (.A(clknet_1_1__leaf__03509_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _19818__88 (.A(clknet_1_1__leaf__03511_),
    .Y(net213));
 sky130_fd_sc_hd__buf_1 _19816_ (.A(clknet_1_1__leaf__05825_),
    .X(_03510_));
 sky130_fd_sc_hd__buf_1 _19817_ (.A(clknet_1_1__leaf__03510_),
    .X(_03511_));
 sky130_fd_sc_hd__inv_2 _19819__89 (.A(clknet_1_1__leaf__03511_),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _19820__90 (.A(clknet_1_0__leaf__03511_),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _19821__91 (.A(clknet_1_0__leaf__03511_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _20339__92 (.A(clknet_1_0__leaf__03511_),
    .Y(net217));
 sky130_fd_sc_hd__nand2_1 _19822_ (.A(_03486_),
    .B(_03485_),
    .Y(_03512_));
 sky130_fd_sc_hd__buf_4 _19823_ (.A(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_4 _19824_ (.A(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _19825_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.spi_buffer[0] ),
    .S(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _19826_ (.A(_03515_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _19827_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.spi_buffer[1] ),
    .S(_03514_),
    .X(_03516_));
 sky130_fd_sc_hd__clkbuf_1 _19828_ (.A(_03516_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _19829_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.spi_buffer[2] ),
    .S(_03514_),
    .X(_03517_));
 sky130_fd_sc_hd__clkbuf_1 _19830_ (.A(_03517_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _19831_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.spi_buffer[3] ),
    .S(_03514_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_1 _19832_ (.A(_03518_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _19833_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.spi_buffer[4] ),
    .S(_03514_),
    .X(_03519_));
 sky130_fd_sc_hd__clkbuf_1 _19834_ (.A(_03519_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _19835_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.spi_buffer[5] ),
    .S(_03514_),
    .X(_03520_));
 sky130_fd_sc_hd__clkbuf_1 _19836_ (.A(_03520_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _19837_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.spi_buffer[6] ),
    .S(_03514_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_1 _19838_ (.A(_03521_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _19839_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.spi_buffer[7] ),
    .S(_03514_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _19840_ (.A(_03522_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _19841_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.spi_buffer[8] ),
    .S(_03514_),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_1 _19842_ (.A(_03523_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _19843_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.spi_buffer[9] ),
    .S(_03514_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _19844_ (.A(_03524_),
    .X(_01095_));
 sky130_fd_sc_hd__clkbuf_4 _19845_ (.A(_03513_),
    .X(_03525_));
 sky130_fd_sc_hd__mux2_1 _19846_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.spi_buffer[10] ),
    .S(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _19847_ (.A(_03526_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _19848_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.spi_buffer[11] ),
    .S(_03525_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_1 _19849_ (.A(_03527_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _19850_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.spi_buffer[12] ),
    .S(_03525_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _19851_ (.A(_03528_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _19852_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.spi_buffer[13] ),
    .S(_03525_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _19853_ (.A(_03529_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _19854_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.spi_buffer[14] ),
    .S(_03525_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _19855_ (.A(_03530_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _19856_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.spi_buffer[15] ),
    .S(_03525_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_1 _19857_ (.A(_03531_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _19858_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.spi_buffer[16] ),
    .S(_03525_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_1 _19859_ (.A(_03532_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _19860_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.spi_buffer[17] ),
    .S(_03525_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_1 _19861_ (.A(_03533_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _19862_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.spi_buffer[18] ),
    .S(_03525_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _19863_ (.A(_03534_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _19864_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.spi_buffer[19] ),
    .S(_03525_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _19865_ (.A(_03535_),
    .X(_01105_));
 sky130_fd_sc_hd__clkbuf_4 _19866_ (.A(_03513_),
    .X(_03536_));
 sky130_fd_sc_hd__mux2_1 _19867_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.spi_buffer[20] ),
    .S(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__clkbuf_1 _19868_ (.A(_03537_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _19869_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.spi_buffer[21] ),
    .S(_03536_),
    .X(_03538_));
 sky130_fd_sc_hd__clkbuf_1 _19870_ (.A(_03538_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _19871_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.spi_buffer[22] ),
    .S(_03536_),
    .X(_03539_));
 sky130_fd_sc_hd__clkbuf_1 _19872_ (.A(_03539_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _19873_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.spi_buffer[23] ),
    .S(_03536_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _19874_ (.A(_03540_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _19875_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.spi_buffer[24] ),
    .S(_03536_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_1 _19876_ (.A(_03541_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _19877_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.spi_buffer[25] ),
    .S(_03536_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_1 _19878_ (.A(_03542_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _19879_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.spi_buffer[26] ),
    .S(_03536_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _19880_ (.A(_03543_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _19881_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.spi_buffer[27] ),
    .S(_03536_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _19882_ (.A(_03544_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _19883_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.spi_buffer[28] ),
    .S(_03536_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _19884_ (.A(_03545_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _19885_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.spi_buffer[29] ),
    .S(_03536_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _19886_ (.A(_03546_),
    .X(_01115_));
 sky130_fd_sc_hd__clkbuf_4 _19887_ (.A(_03513_),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_1 _19888_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.spi_buffer[30] ),
    .S(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_1 _19889_ (.A(_03548_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _19890_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.spi_buffer[31] ),
    .S(_03547_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _19891_ (.A(_03549_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _19892_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.spi_buffer[32] ),
    .S(_03547_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _19893_ (.A(_03550_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _19894_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.spi_buffer[33] ),
    .S(_03547_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _19895_ (.A(_03551_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _19896_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.spi_buffer[34] ),
    .S(_03547_),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_1 _19897_ (.A(_03552_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _19898_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.spi_buffer[35] ),
    .S(_03547_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _19899_ (.A(_03553_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _19900_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.spi_buffer[36] ),
    .S(_03547_),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _19901_ (.A(_03554_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _19902_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.spi_buffer[37] ),
    .S(_03547_),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_1 _19903_ (.A(_03555_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _19904_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.spi_buffer[38] ),
    .S(_03547_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _19905_ (.A(_03556_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _19906_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.spi_buffer[39] ),
    .S(_03547_),
    .X(_03557_));
 sky130_fd_sc_hd__clkbuf_1 _19907_ (.A(_03557_),
    .X(_01125_));
 sky130_fd_sc_hd__clkbuf_4 _19908_ (.A(_03513_),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _19909_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.spi_buffer[40] ),
    .S(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__clkbuf_1 _19910_ (.A(_03559_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _19911_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.spi_buffer[41] ),
    .S(_03558_),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _19912_ (.A(_03560_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _19913_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.spi_buffer[42] ),
    .S(_03558_),
    .X(_03561_));
 sky130_fd_sc_hd__clkbuf_1 _19914_ (.A(_03561_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.spi_buffer[43] ),
    .S(_03558_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_1 _19916_ (.A(_03562_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _19917_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.spi_buffer[44] ),
    .S(_03558_),
    .X(_03563_));
 sky130_fd_sc_hd__clkbuf_1 _19918_ (.A(_03563_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _19919_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.spi_buffer[45] ),
    .S(_03558_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _19920_ (.A(_03564_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _19921_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.spi_buffer[46] ),
    .S(_03558_),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _19922_ (.A(_03565_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _19923_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.spi_buffer[47] ),
    .S(_03558_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _19924_ (.A(_03566_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _19925_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.spi_buffer[48] ),
    .S(_03558_),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _19926_ (.A(_03567_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _19927_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.spi_buffer[49] ),
    .S(_03558_),
    .X(_03568_));
 sky130_fd_sc_hd__clkbuf_1 _19928_ (.A(_03568_),
    .X(_01135_));
 sky130_fd_sc_hd__clkbuf_4 _19929_ (.A(_03513_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _19930_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.spi_buffer[50] ),
    .S(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _19931_ (.A(_03570_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _19932_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.spi_buffer[51] ),
    .S(_03569_),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_1 _19933_ (.A(_03571_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _19934_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.spi_buffer[52] ),
    .S(_03569_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _19935_ (.A(_03572_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _19936_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.spi_buffer[53] ),
    .S(_03569_),
    .X(_03573_));
 sky130_fd_sc_hd__clkbuf_1 _19937_ (.A(_03573_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _19938_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.spi_buffer[54] ),
    .S(_03569_),
    .X(_03574_));
 sky130_fd_sc_hd__clkbuf_1 _19939_ (.A(_03574_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _19940_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.spi_buffer[55] ),
    .S(_03569_),
    .X(_03575_));
 sky130_fd_sc_hd__clkbuf_1 _19941_ (.A(_03575_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _19942_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.spi_buffer[56] ),
    .S(_03569_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_1 _19943_ (.A(_03576_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _19944_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.spi_buffer[57] ),
    .S(_03569_),
    .X(_03577_));
 sky130_fd_sc_hd__clkbuf_1 _19945_ (.A(_03577_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _19946_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.spi_buffer[58] ),
    .S(_03569_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_1 _19947_ (.A(_03578_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _19948_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.spi_buffer[59] ),
    .S(_03569_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_1 _19949_ (.A(_03579_),
    .X(_01145_));
 sky130_fd_sc_hd__clkbuf_4 _19950_ (.A(_03512_),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_1 _19951_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.spi_buffer[60] ),
    .S(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__clkbuf_1 _19952_ (.A(_03581_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _19953_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.spi_buffer[61] ),
    .S(_03580_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _19954_ (.A(_03582_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _19955_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.spi_buffer[62] ),
    .S(_03580_),
    .X(_03583_));
 sky130_fd_sc_hd__clkbuf_1 _19956_ (.A(_03583_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _19957_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.spi_buffer[63] ),
    .S(_03580_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _19958_ (.A(_03584_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _19959_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.spi_buffer[64] ),
    .S(_03580_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_1 _19960_ (.A(_03585_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _19961_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.spi_buffer[65] ),
    .S(_03580_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _19962_ (.A(_03586_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _19963_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.spi_buffer[66] ),
    .S(_03580_),
    .X(_03587_));
 sky130_fd_sc_hd__clkbuf_1 _19964_ (.A(_03587_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _19965_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.spi_buffer[67] ),
    .S(_03580_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _19966_ (.A(_03588_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _19967_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.spi_buffer[68] ),
    .S(_03580_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _19968_ (.A(_03589_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _19969_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.spi_buffer[69] ),
    .S(_03580_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _19970_ (.A(_03590_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _19971_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.spi_buffer[70] ),
    .S(_03513_),
    .X(_03591_));
 sky130_fd_sc_hd__clkbuf_1 _19972_ (.A(_03591_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _19973_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.spi_buffer[71] ),
    .S(_03513_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _19974_ (.A(_03592_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _19975_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.spi_buffer[72] ),
    .S(_03513_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _19976_ (.A(_03593_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _19977_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.spi_buffer[73] ),
    .S(_03513_),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_1 _19978_ (.A(_03594_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _19979_ (.A0(_05734_),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_03122_),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_1 _19980_ (.A(_03595_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _19981_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_08185_),
    .X(_03596_));
 sky130_fd_sc_hd__clkbuf_1 _19982_ (.A(_03596_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _19983_ (.A0(net54),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_03122_),
    .X(_03597_));
 sky130_fd_sc_hd__clkbuf_1 _19984_ (.A(_03597_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _19985_ (.A0(\rbzero.pov.ss_buffer[1] ),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_08185_),
    .X(_03598_));
 sky130_fd_sc_hd__clkbuf_1 _19986_ (.A(_03598_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _19987_ (.A0(net56),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_03122_),
    .X(_03599_));
 sky130_fd_sc_hd__clkbuf_1 _19988_ (.A(_03599_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _19989_ (.A0(\rbzero.pov.sclk_buffer[1] ),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_08185_),
    .X(_03600_));
 sky130_fd_sc_hd__clkbuf_1 _19990_ (.A(_03600_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _19991_ (.A0(\rbzero.pov.sclk_buffer[2] ),
    .A1(\rbzero.pov.sclk_buffer[1] ),
    .S(_08185_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _19992_ (.A(_03601_),
    .X(_01166_));
 sky130_fd_sc_hd__and2_2 _19993_ (.A(\rbzero.pov.ready ),
    .B(_03482_),
    .X(_03602_));
 sky130_fd_sc_hd__o21ai_4 _19994_ (.A1(net40),
    .A2(_03602_),
    .B1(_03140_),
    .Y(_03603_));
 sky130_fd_sc_hd__clkbuf_4 _19995_ (.A(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__inv_2 _19996_ (.A(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_03605_));
 sky130_fd_sc_hd__clkbuf_4 _19997_ (.A(_03483_),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_1 _19998_ (.A0(_03605_),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__nand2_1 _19999_ (.A(_03605_),
    .B(_03604_),
    .Y(_03608_));
 sky130_fd_sc_hd__o211a_1 _20000_ (.A1(_03604_),
    .A2(_03607_),
    .B1(_03608_),
    .C1(_03319_),
    .X(_01167_));
 sky130_fd_sc_hd__inv_2 _20001_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .Y(_03609_));
 sky130_fd_sc_hd__o21a_1 _20002_ (.A1(net40),
    .A2(_03602_),
    .B1(_03140_),
    .X(_03610_));
 sky130_fd_sc_hd__nand2_1 _20003_ (.A(\rbzero.pov.ready_buffer[60] ),
    .B(_03483_),
    .Y(_03611_));
 sky130_fd_sc_hd__o211a_1 _20004_ (.A1(_08261_),
    .A2(_03606_),
    .B1(_03610_),
    .C1(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__buf_4 _20005_ (.A(_04469_),
    .X(_03613_));
 sky130_fd_sc_hd__a211oi_1 _20006_ (.A1(_03609_),
    .A2(_03604_),
    .B1(_03612_),
    .C1(_03613_),
    .Y(_01168_));
 sky130_fd_sc_hd__buf_2 _20007_ (.A(_03610_),
    .X(_03614_));
 sky130_fd_sc_hd__nor2_1 _20008_ (.A(_08247_),
    .B(_03606_),
    .Y(_03615_));
 sky130_fd_sc_hd__a211o_1 _20009_ (.A1(\rbzero.pov.ready_buffer[61] ),
    .A2(_03484_),
    .B1(_03603_),
    .C1(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__o211a_1 _20010_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_03614_),
    .B1(_03616_),
    .C1(_03319_),
    .X(_01169_));
 sky130_fd_sc_hd__nor2_1 _20011_ (.A(_03156_),
    .B(_03481_),
    .Y(_03617_));
 sky130_fd_sc_hd__clkbuf_4 _20012_ (.A(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _20013_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(_08283_),
    .S(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__nand2_1 _20014_ (.A(_08284_),
    .B(_03604_),
    .Y(_03620_));
 sky130_fd_sc_hd__clkbuf_4 _20015_ (.A(_09808_),
    .X(_03621_));
 sky130_fd_sc_hd__o211a_1 _20016_ (.A1(_03604_),
    .A2(_03619_),
    .B1(_03620_),
    .C1(_03621_),
    .X(_01170_));
 sky130_fd_sc_hd__nor2_1 _20017_ (.A(_08389_),
    .B(_03606_),
    .Y(_03622_));
 sky130_fd_sc_hd__a211o_1 _20018_ (.A1(\rbzero.pov.ready_buffer[63] ),
    .A2(_03484_),
    .B1(_03603_),
    .C1(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__o211a_1 _20019_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_03614_),
    .B1(_03623_),
    .C1(_03621_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _20020_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(_08405_),
    .S(_03618_),
    .X(_03624_));
 sky130_fd_sc_hd__nand2_1 _20021_ (.A(_08406_),
    .B(_03603_),
    .Y(_03625_));
 sky130_fd_sc_hd__o211a_1 _20022_ (.A1(_03604_),
    .A2(_03624_),
    .B1(_03625_),
    .C1(_03621_),
    .X(_01172_));
 sky130_fd_sc_hd__nor2_1 _20023_ (.A(_08420_),
    .B(_03606_),
    .Y(_03626_));
 sky130_fd_sc_hd__a211o_1 _20024_ (.A1(\rbzero.pov.ready_buffer[65] ),
    .A2(_03484_),
    .B1(_03603_),
    .C1(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__o211a_1 _20025_ (.A1(\rbzero.debug_overlay.playerX[-3] ),
    .A2(_03614_),
    .B1(_03627_),
    .C1(_03621_),
    .X(_01173_));
 sky130_fd_sc_hd__nor2_1 _20026_ (.A(_08530_),
    .B(_03606_),
    .Y(_03628_));
 sky130_fd_sc_hd__a211o_1 _20027_ (.A1(\rbzero.pov.ready_buffer[66] ),
    .A2(_03484_),
    .B1(_03603_),
    .C1(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__o211a_1 _20028_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_03614_),
    .B1(_03629_),
    .C1(_03621_),
    .X(_01174_));
 sky130_fd_sc_hd__buf_4 _20029_ (.A(_03617_),
    .X(_03630_));
 sky130_fd_sc_hd__nand2_1 _20030_ (.A(_08539_),
    .B(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__o211a_1 _20031_ (.A1(\rbzero.pov.ready_buffer[67] ),
    .A2(_03618_),
    .B1(_03610_),
    .C1(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__a211o_1 _20032_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_03604_),
    .B1(_03632_),
    .C1(_09813_),
    .X(_01175_));
 sky130_fd_sc_hd__and2_1 _20033_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_08513_),
    .X(_03633_));
 sky130_fd_sc_hd__or2_1 _20034_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_08513_),
    .X(_03634_));
 sky130_fd_sc_hd__or3b_1 _20035_ (.A(_03633_),
    .B(_03483_),
    .C_N(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__o211a_1 _20036_ (.A1(\rbzero.pov.ready_buffer[68] ),
    .A2(_03618_),
    .B1(_03610_),
    .C1(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__a211o_1 _20037_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03604_),
    .B1(_03636_),
    .C1(_09813_),
    .X(_01176_));
 sky130_fd_sc_hd__nor2_1 _20038_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03634_),
    .Y(_03637_));
 sky130_fd_sc_hd__and2_1 _20039_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03634_),
    .X(_03638_));
 sky130_fd_sc_hd__or2_1 _20040_ (.A(\rbzero.pov.ready_buffer[69] ),
    .B(_03630_),
    .X(_03639_));
 sky130_fd_sc_hd__o311a_1 _20041_ (.A1(_03484_),
    .A2(_03637_),
    .A3(_03638_),
    .B1(_03614_),
    .C1(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__a211o_1 _20042_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03604_),
    .B1(_03640_),
    .C1(_09813_),
    .X(_01177_));
 sky130_fd_sc_hd__or3_1 _20043_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .B(\rbzero.debug_overlay.playerX[1] ),
    .C(_03634_),
    .X(_03641_));
 sky130_fd_sc_hd__o21ai_1 _20044_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03634_),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .Y(_03642_));
 sky130_fd_sc_hd__a21oi_1 _20045_ (.A1(_03641_),
    .A2(_03642_),
    .B1(_03606_),
    .Y(_03643_));
 sky130_fd_sc_hd__a211o_1 _20046_ (.A1(\rbzero.pov.ready_buffer[70] ),
    .A2(_03484_),
    .B1(_03603_),
    .C1(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__o211a_1 _20047_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_03614_),
    .B1(_03644_),
    .C1(_03621_),
    .X(_01178_));
 sky130_fd_sc_hd__nor2_1 _20048_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_03641_),
    .Y(_03645_));
 sky130_fd_sc_hd__a21o_1 _20049_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03641_),
    .B1(_03483_),
    .X(_03646_));
 sky130_fd_sc_hd__o221a_1 _20050_ (.A1(\rbzero.pov.ready_buffer[71] ),
    .A2(_03618_),
    .B1(_03645_),
    .B2(_03646_),
    .C1(_03614_),
    .X(_03647_));
 sky130_fd_sc_hd__a211o_1 _20051_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03604_),
    .B1(_03647_),
    .C1(_09813_),
    .X(_01179_));
 sky130_fd_sc_hd__nor2_1 _20052_ (.A(_03481_),
    .B(_03645_),
    .Y(_03648_));
 sky130_fd_sc_hd__o21a_1 _20053_ (.A1(_03603_),
    .A2(_03648_),
    .B1(\rbzero.debug_overlay.playerX[4] ),
    .X(_03649_));
 sky130_fd_sc_hd__a21o_1 _20054_ (.A1(_04739_),
    .A2(_03645_),
    .B1(_03481_),
    .X(_03650_));
 sky130_fd_sc_hd__o211a_1 _20055_ (.A1(\rbzero.pov.ready_buffer[72] ),
    .A2(_03618_),
    .B1(_03614_),
    .C1(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__o21a_1 _20056_ (.A1(_03649_),
    .A2(_03651_),
    .B1(_03143_),
    .X(_01180_));
 sky130_fd_sc_hd__inv_2 _20057_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .Y(_03652_));
 sky130_fd_sc_hd__a21oi_1 _20058_ (.A1(_03614_),
    .A2(_03650_),
    .B1(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__a31o_1 _20059_ (.A1(_03652_),
    .A2(_04739_),
    .A3(_03645_),
    .B1(_03483_),
    .X(_03654_));
 sky130_fd_sc_hd__o211a_1 _20060_ (.A1(\rbzero.pov.ready_buffer[73] ),
    .A2(_03618_),
    .B1(_03614_),
    .C1(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__o21a_1 _20061_ (.A1(_03653_),
    .A2(_03655_),
    .B1(_03143_),
    .X(_01181_));
 sky130_fd_sc_hd__o21ai_4 _20062_ (.A1(net41),
    .A2(_03602_),
    .B1(_03140_),
    .Y(_03656_));
 sky130_fd_sc_hd__clkbuf_4 _20063_ (.A(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _20064_ (.A0(_08308_),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_03606_),
    .X(_03658_));
 sky130_fd_sc_hd__nand2_1 _20065_ (.A(_08308_),
    .B(_03657_),
    .Y(_03659_));
 sky130_fd_sc_hd__o211a_1 _20066_ (.A1(_03657_),
    .A2(_03658_),
    .B1(_03659_),
    .C1(_03621_),
    .X(_01182_));
 sky130_fd_sc_hd__o21a_1 _20067_ (.A1(net41),
    .A2(_03602_),
    .B1(_03139_),
    .X(_03660_));
 sky130_fd_sc_hd__clkbuf_4 _20068_ (.A(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__nor2_1 _20069_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand2_1 _20070_ (.A(\rbzero.pov.ready_buffer[45] ),
    .B(_03483_),
    .Y(_03663_));
 sky130_fd_sc_hd__o211a_1 _20071_ (.A1(_08263_),
    .A2(_03484_),
    .B1(_03661_),
    .C1(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__nor3_1 _20072_ (.A(_03613_),
    .B(_03662_),
    .C(_03664_),
    .Y(_01183_));
 sky130_fd_sc_hd__or2_1 _20073_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(_03660_),
    .X(_03665_));
 sky130_fd_sc_hd__a21oi_1 _20074_ (.A1(_08254_),
    .A2(_08255_),
    .B1(_03483_),
    .Y(_03666_));
 sky130_fd_sc_hd__a211o_1 _20075_ (.A1(\rbzero.pov.ready_buffer[46] ),
    .A2(_03483_),
    .B1(_03656_),
    .C1(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__and3_1 _20076_ (.A(_09810_),
    .B(_03665_),
    .C(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_1 _20077_ (.A(_03668_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _20078_ (.A0(\rbzero.pov.ready_buffer[47] ),
    .A1(_08278_),
    .S(_03630_),
    .X(_03669_));
 sky130_fd_sc_hd__nand2_1 _20079_ (.A(_08275_),
    .B(_03657_),
    .Y(_03670_));
 sky130_fd_sc_hd__o211a_1 _20080_ (.A1(_03657_),
    .A2(_03669_),
    .B1(_03670_),
    .C1(_03621_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _20081_ (.A0(\rbzero.pov.ready_buffer[48] ),
    .A1(_08391_),
    .S(_03630_),
    .X(_03671_));
 sky130_fd_sc_hd__nand2_1 _20082_ (.A(_09302_),
    .B(_03657_),
    .Y(_03672_));
 sky130_fd_sc_hd__o211a_1 _20083_ (.A1(_03657_),
    .A2(_03671_),
    .B1(_03672_),
    .C1(_03621_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _20084_ (.A0(\rbzero.pov.ready_buffer[49] ),
    .A1(_08399_),
    .S(_03630_),
    .X(_03673_));
 sky130_fd_sc_hd__nand2_1 _20085_ (.A(_09423_),
    .B(_03656_),
    .Y(_03674_));
 sky130_fd_sc_hd__o211a_1 _20086_ (.A1(_03657_),
    .A2(_03673_),
    .B1(_03674_),
    .C1(_03621_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _20087_ (.A0(\rbzero.pov.ready_buffer[50] ),
    .A1(_08424_),
    .S(_03630_),
    .X(_03675_));
 sky130_fd_sc_hd__nand2_1 _20088_ (.A(_04752_),
    .B(_03656_),
    .Y(_03676_));
 sky130_fd_sc_hd__clkbuf_4 _20089_ (.A(_09808_),
    .X(_03677_));
 sky130_fd_sc_hd__o211a_1 _20090_ (.A1(_03657_),
    .A2(_03675_),
    .B1(_03676_),
    .C1(_03677_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _20091_ (.A0(\rbzero.pov.ready_buffer[51] ),
    .A1(_08532_),
    .S(_03630_),
    .X(_03678_));
 sky130_fd_sc_hd__nand2_1 _20092_ (.A(_04746_),
    .B(_03656_),
    .Y(_03679_));
 sky130_fd_sc_hd__o211a_1 _20093_ (.A1(_03657_),
    .A2(_03678_),
    .B1(_03679_),
    .C1(_03677_),
    .X(_01189_));
 sky130_fd_sc_hd__and2_1 _20094_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(_03656_),
    .X(_03680_));
 sky130_fd_sc_hd__nand2_1 _20095_ (.A(_08542_),
    .B(_03617_),
    .Y(_03681_));
 sky130_fd_sc_hd__o211a_1 _20096_ (.A1(\rbzero.pov.ready_buffer[52] ),
    .A2(_03630_),
    .B1(_03660_),
    .C1(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__or3_1 _20097_ (.A(_03122_),
    .B(_03680_),
    .C(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _20098_ (.A(_03683_),
    .X(_01190_));
 sky130_fd_sc_hd__or2_1 _20099_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08514_),
    .X(_03684_));
 sky130_fd_sc_hd__nand2_1 _20100_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08514_),
    .Y(_03685_));
 sky130_fd_sc_hd__a21oi_1 _20101_ (.A1(_03684_),
    .A2(_03685_),
    .B1(_03606_),
    .Y(_03686_));
 sky130_fd_sc_hd__a211o_1 _20102_ (.A1(\rbzero.pov.ready_buffer[53] ),
    .A2(_03484_),
    .B1(_03656_),
    .C1(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__o211a_1 _20103_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_03661_),
    .B1(_03687_),
    .C1(_03677_),
    .X(_01191_));
 sky130_fd_sc_hd__o21ai_1 _20104_ (.A1(_04734_),
    .A2(_03684_),
    .B1(_03630_),
    .Y(_03688_));
 sky130_fd_sc_hd__a21o_1 _20105_ (.A1(_04734_),
    .A2(_03684_),
    .B1(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__o211a_1 _20106_ (.A1(\rbzero.pov.ready_buffer[54] ),
    .A2(_03618_),
    .B1(_03661_),
    .C1(_03689_),
    .X(_03690_));
 sky130_fd_sc_hd__a211o_1 _20107_ (.A1(_04734_),
    .A2(_03657_),
    .B1(_03690_),
    .C1(_09813_),
    .X(_01192_));
 sky130_fd_sc_hd__or3_1 _20108_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(_04734_),
    .C(_03684_),
    .X(_03691_));
 sky130_fd_sc_hd__o21ai_1 _20109_ (.A1(_04734_),
    .A2(_03684_),
    .B1(\rbzero.debug_overlay.playerY[2] ),
    .Y(_03692_));
 sky130_fd_sc_hd__a21oi_1 _20110_ (.A1(_03691_),
    .A2(_03692_),
    .B1(_03606_),
    .Y(_03693_));
 sky130_fd_sc_hd__a211o_1 _20111_ (.A1(\rbzero.pov.ready_buffer[55] ),
    .A2(_03484_),
    .B1(_03656_),
    .C1(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__o211a_1 _20112_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_03661_),
    .B1(_03694_),
    .C1(_03677_),
    .X(_01193_));
 sky130_fd_sc_hd__nor2_1 _20113_ (.A(_06238_),
    .B(_03661_),
    .Y(_03695_));
 sky130_fd_sc_hd__nor2_1 _20114_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .B(_03691_),
    .Y(_03696_));
 sky130_fd_sc_hd__a21o_1 _20115_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03691_),
    .B1(_03482_),
    .X(_03697_));
 sky130_fd_sc_hd__o221a_1 _20116_ (.A1(\rbzero.pov.ready_buffer[56] ),
    .A2(_03630_),
    .B1(_03696_),
    .B2(_03697_),
    .C1(_03660_),
    .X(_03698_));
 sky130_fd_sc_hd__or3_1 _20117_ (.A(_03122_),
    .B(_03695_),
    .C(_03698_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_1 _20118_ (.A(_03699_),
    .X(_01194_));
 sky130_fd_sc_hd__o21a_1 _20119_ (.A1(_03481_),
    .A2(_03696_),
    .B1(_03661_),
    .X(_03700_));
 sky130_fd_sc_hd__nor2_1 _20120_ (.A(_04725_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__a21o_1 _20121_ (.A1(_04725_),
    .A2(_03696_),
    .B1(_03481_),
    .X(_03702_));
 sky130_fd_sc_hd__o211a_1 _20122_ (.A1(\rbzero.pov.ready_buffer[57] ),
    .A2(_03618_),
    .B1(_03661_),
    .C1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__o21a_1 _20123_ (.A1(_03701_),
    .A2(_03703_),
    .B1(_03143_),
    .X(_01195_));
 sky130_fd_sc_hd__a21oi_1 _20124_ (.A1(_03661_),
    .A2(_03702_),
    .B1(_06245_),
    .Y(_03704_));
 sky130_fd_sc_hd__a31o_1 _20125_ (.A1(_06245_),
    .A2(_04725_),
    .A3(_03696_),
    .B1(_03483_),
    .X(_03705_));
 sky130_fd_sc_hd__o211a_1 _20126_ (.A1(\rbzero.pov.ready_buffer[58] ),
    .A2(_03618_),
    .B1(_03661_),
    .C1(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__o21a_1 _20127_ (.A1(_03704_),
    .A2(_03706_),
    .B1(_03143_),
    .X(_01196_));
 sky130_fd_sc_hd__nand2_4 _20128_ (.A(_03140_),
    .B(_03602_),
    .Y(_03707_));
 sky130_fd_sc_hd__clkbuf_4 _20129_ (.A(_03707_),
    .X(_03708_));
 sky130_fd_sc_hd__and3_1 _20130_ (.A(\rbzero.pov.ready ),
    .B(_03139_),
    .C(_03481_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_4 _20131_ (.A(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_4 _20132_ (.A(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_2 _20133_ (.A(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__or2_1 _20134_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__o211a_1 _20135_ (.A1(\rbzero.pov.ready_buffer[33] ),
    .A2(_03708_),
    .B1(_03713_),
    .C1(_03677_),
    .X(_01197_));
 sky130_fd_sc_hd__or2_1 _20136_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(_03712_),
    .X(_03714_));
 sky130_fd_sc_hd__o211a_1 _20137_ (.A1(\rbzero.pov.ready_buffer[34] ),
    .A2(_03708_),
    .B1(_03714_),
    .C1(_03677_),
    .X(_01198_));
 sky130_fd_sc_hd__or2_1 _20138_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(_03712_),
    .X(_03715_));
 sky130_fd_sc_hd__o211a_1 _20139_ (.A1(\rbzero.pov.ready_buffer[35] ),
    .A2(_03708_),
    .B1(_03715_),
    .C1(_03677_),
    .X(_01199_));
 sky130_fd_sc_hd__or2_1 _20140_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(_03712_),
    .X(_03716_));
 sky130_fd_sc_hd__o211a_1 _20141_ (.A1(\rbzero.pov.ready_buffer[36] ),
    .A2(_03708_),
    .B1(_03716_),
    .C1(_03677_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _20142_ (.A0(\rbzero.debug_overlay.facingX[-5] ),
    .A1(\rbzero.pov.ready_buffer[37] ),
    .S(_03711_),
    .X(_03717_));
 sky130_fd_sc_hd__or2_1 _20143_ (.A(_03322_),
    .B(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_1 _20144_ (.A(_03718_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _20145_ (.A0(\rbzero.debug_overlay.facingX[-4] ),
    .A1(\rbzero.pov.ready_buffer[38] ),
    .S(_03711_),
    .X(_03719_));
 sky130_fd_sc_hd__or2_1 _20146_ (.A(_03322_),
    .B(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _20147_ (.A(_03720_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _20148_ (.A0(\rbzero.debug_overlay.facingX[-3] ),
    .A1(\rbzero.pov.ready_buffer[39] ),
    .S(_03711_),
    .X(_03721_));
 sky130_fd_sc_hd__or2_1 _20149_ (.A(_03322_),
    .B(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_1 _20150_ (.A(_03722_),
    .X(_01203_));
 sky130_fd_sc_hd__or2_1 _20151_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(_03712_),
    .X(_03723_));
 sky130_fd_sc_hd__o211a_1 _20152_ (.A1(\rbzero.pov.ready_buffer[40] ),
    .A2(_03708_),
    .B1(_03723_),
    .C1(_03677_),
    .X(_01204_));
 sky130_fd_sc_hd__buf_2 _20153_ (.A(_04469_),
    .X(_03724_));
 sky130_fd_sc_hd__buf_4 _20154_ (.A(_03710_),
    .X(_03725_));
 sky130_fd_sc_hd__mux2_1 _20155_ (.A0(\rbzero.debug_overlay.facingX[-1] ),
    .A1(\rbzero.pov.ready_buffer[41] ),
    .S(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__or2_1 _20156_ (.A(_03724_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _20157_ (.A(_03727_),
    .X(_01205_));
 sky130_fd_sc_hd__or2_1 _20158_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(_03712_),
    .X(_03728_));
 sky130_fd_sc_hd__o211a_1 _20159_ (.A1(\rbzero.pov.ready_buffer[42] ),
    .A2(_03708_),
    .B1(_03728_),
    .C1(_03677_),
    .X(_01206_));
 sky130_fd_sc_hd__or2_1 _20160_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(_03712_),
    .X(_03729_));
 sky130_fd_sc_hd__clkbuf_4 _20161_ (.A(_09808_),
    .X(_03730_));
 sky130_fd_sc_hd__o211a_1 _20162_ (.A1(\rbzero.pov.ready_buffer[43] ),
    .A2(_03708_),
    .B1(_03729_),
    .C1(_03730_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _20163_ (.A0(\rbzero.debug_overlay.facingY[-9] ),
    .A1(\rbzero.pov.ready_buffer[22] ),
    .S(_03725_),
    .X(_03731_));
 sky130_fd_sc_hd__or2_1 _20164_ (.A(_03724_),
    .B(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__clkbuf_1 _20165_ (.A(_03732_),
    .X(_01208_));
 sky130_fd_sc_hd__or2_1 _20166_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_03712_),
    .X(_03733_));
 sky130_fd_sc_hd__o211a_1 _20167_ (.A1(\rbzero.pov.ready_buffer[23] ),
    .A2(_03708_),
    .B1(_03733_),
    .C1(_03730_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _20168_ (.A0(\rbzero.debug_overlay.facingY[-7] ),
    .A1(\rbzero.pov.ready_buffer[24] ),
    .S(_03725_),
    .X(_03734_));
 sky130_fd_sc_hd__or2_1 _20169_ (.A(_03724_),
    .B(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__clkbuf_1 _20170_ (.A(_03735_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _20171_ (.A0(\rbzero.debug_overlay.facingY[-6] ),
    .A1(\rbzero.pov.ready_buffer[25] ),
    .S(_03725_),
    .X(_03736_));
 sky130_fd_sc_hd__or2_1 _20172_ (.A(_03724_),
    .B(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__clkbuf_1 _20173_ (.A(_03737_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _20174_ (.A0(\rbzero.debug_overlay.facingY[-5] ),
    .A1(\rbzero.pov.ready_buffer[26] ),
    .S(_03725_),
    .X(_03738_));
 sky130_fd_sc_hd__or2_1 _20175_ (.A(_03724_),
    .B(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__clkbuf_1 _20176_ (.A(_03739_),
    .X(_01212_));
 sky130_fd_sc_hd__or2_1 _20177_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(_03712_),
    .X(_03740_));
 sky130_fd_sc_hd__o211a_1 _20178_ (.A1(\rbzero.pov.ready_buffer[27] ),
    .A2(_03708_),
    .B1(_03740_),
    .C1(_03730_),
    .X(_01213_));
 sky130_fd_sc_hd__or2_1 _20179_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(_03712_),
    .X(_03741_));
 sky130_fd_sc_hd__o211a_1 _20180_ (.A1(\rbzero.pov.ready_buffer[28] ),
    .A2(_03708_),
    .B1(_03741_),
    .C1(_03730_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _20181_ (.A0(\rbzero.debug_overlay.facingY[-2] ),
    .A1(\rbzero.pov.ready_buffer[29] ),
    .S(_03725_),
    .X(_03742_));
 sky130_fd_sc_hd__or2_1 _20182_ (.A(_03724_),
    .B(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__clkbuf_1 _20183_ (.A(_03743_),
    .X(_01215_));
 sky130_fd_sc_hd__buf_2 _20184_ (.A(_03707_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_2 _20185_ (.A(_03711_),
    .X(_03745_));
 sky130_fd_sc_hd__or2_1 _20186_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__o211a_1 _20187_ (.A1(\rbzero.pov.ready_buffer[30] ),
    .A2(_03744_),
    .B1(_03746_),
    .C1(_03730_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _20188_ (.A0(\rbzero.debug_overlay.facingY[0] ),
    .A1(\rbzero.pov.ready_buffer[31] ),
    .S(_03725_),
    .X(_03747_));
 sky130_fd_sc_hd__or2_1 _20189_ (.A(_03724_),
    .B(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__clkbuf_1 _20190_ (.A(_03748_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _20191_ (.A0(\rbzero.debug_overlay.facingY[10] ),
    .A1(\rbzero.pov.ready_buffer[32] ),
    .S(_03725_),
    .X(_03749_));
 sky130_fd_sc_hd__or2_1 _20192_ (.A(_03724_),
    .B(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__clkbuf_1 _20193_ (.A(_03750_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _20194_ (.A0(\rbzero.debug_overlay.vplaneX[-9] ),
    .A1(\rbzero.pov.ready_buffer[11] ),
    .S(_03725_),
    .X(_03751_));
 sky130_fd_sc_hd__or2_1 _20195_ (.A(_03724_),
    .B(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _20196_ (.A(_03752_),
    .X(_01219_));
 sky130_fd_sc_hd__or2_1 _20197_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(_03745_),
    .X(_03753_));
 sky130_fd_sc_hd__o211a_1 _20198_ (.A1(\rbzero.pov.ready_buffer[12] ),
    .A2(_03744_),
    .B1(_03753_),
    .C1(_03730_),
    .X(_01220_));
 sky130_fd_sc_hd__or2_1 _20199_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_03745_),
    .X(_03754_));
 sky130_fd_sc_hd__o211a_1 _20200_ (.A1(\rbzero.pov.ready_buffer[13] ),
    .A2(_03744_),
    .B1(_03754_),
    .C1(_03730_),
    .X(_01221_));
 sky130_fd_sc_hd__or2_1 _20201_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_03745_),
    .X(_03755_));
 sky130_fd_sc_hd__o211a_1 _20202_ (.A1(\rbzero.pov.ready_buffer[14] ),
    .A2(_03744_),
    .B1(_03755_),
    .C1(_03730_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _20203_ (.A0(_05153_),
    .A1(\rbzero.pov.ready_buffer[15] ),
    .S(_03725_),
    .X(_03756_));
 sky130_fd_sc_hd__or2_1 _20204_ (.A(_03724_),
    .B(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _20205_ (.A(_03757_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _20206_ (.A0(\rbzero.debug_overlay.vplaneX[-4] ),
    .A1(\rbzero.pov.ready_buffer[16] ),
    .S(_03710_),
    .X(_03758_));
 sky130_fd_sc_hd__or2_1 _20207_ (.A(_04470_),
    .B(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_1 _20208_ (.A(_03759_),
    .X(_01224_));
 sky130_fd_sc_hd__or2_1 _20209_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(_03745_),
    .X(_03760_));
 sky130_fd_sc_hd__o211a_1 _20210_ (.A1(\rbzero.pov.ready_buffer[17] ),
    .A2(_03744_),
    .B1(_03760_),
    .C1(_03730_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _20211_ (.A0(_02577_),
    .A1(\rbzero.pov.ready_buffer[18] ),
    .S(_03710_),
    .X(_03761_));
 sky130_fd_sc_hd__or2_1 _20212_ (.A(_04470_),
    .B(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _20213_ (.A(_03762_),
    .X(_01226_));
 sky130_fd_sc_hd__or2_1 _20214_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_03745_),
    .X(_03763_));
 sky130_fd_sc_hd__o211a_1 _20215_ (.A1(\rbzero.pov.ready_buffer[19] ),
    .A2(_03744_),
    .B1(_03763_),
    .C1(_03730_),
    .X(_01227_));
 sky130_fd_sc_hd__or2_1 _20216_ (.A(_02598_),
    .B(_03745_),
    .X(_03764_));
 sky130_fd_sc_hd__buf_4 _20217_ (.A(_09808_),
    .X(_03765_));
 sky130_fd_sc_hd__o211a_1 _20218_ (.A1(\rbzero.pov.ready_buffer[20] ),
    .A2(_03744_),
    .B1(_03764_),
    .C1(_03765_),
    .X(_01228_));
 sky130_fd_sc_hd__or2_1 _20219_ (.A(_02629_),
    .B(_03745_),
    .X(_03766_));
 sky130_fd_sc_hd__o211a_1 _20220_ (.A1(\rbzero.pov.ready_buffer[21] ),
    .A2(_03744_),
    .B1(_03766_),
    .C1(_03765_),
    .X(_01229_));
 sky130_fd_sc_hd__or2_1 _20221_ (.A(_05172_),
    .B(_03745_),
    .X(_03767_));
 sky130_fd_sc_hd__o211a_1 _20222_ (.A1(\rbzero.pov.ready_buffer[0] ),
    .A2(_03744_),
    .B1(_03767_),
    .C1(_03765_),
    .X(_01230_));
 sky130_fd_sc_hd__or2_1 _20223_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_03745_),
    .X(_03768_));
 sky130_fd_sc_hd__o211a_1 _20224_ (.A1(\rbzero.pov.ready_buffer[1] ),
    .A2(_03744_),
    .B1(_03768_),
    .C1(_03765_),
    .X(_01231_));
 sky130_fd_sc_hd__or2_1 _20225_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03711_),
    .X(_03769_));
 sky130_fd_sc_hd__o211a_1 _20226_ (.A1(\rbzero.pov.ready_buffer[2] ),
    .A2(_03707_),
    .B1(_03769_),
    .C1(_03765_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _20227_ (.A0(\rbzero.debug_overlay.vplaneY[-6] ),
    .A1(\rbzero.pov.ready_buffer[3] ),
    .S(_03710_),
    .X(_03770_));
 sky130_fd_sc_hd__or2_1 _20228_ (.A(_04470_),
    .B(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__clkbuf_1 _20229_ (.A(_03771_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _20230_ (.A0(_05173_),
    .A1(\rbzero.pov.ready_buffer[4] ),
    .S(_03710_),
    .X(_03772_));
 sky130_fd_sc_hd__or2_1 _20231_ (.A(_04470_),
    .B(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__clkbuf_1 _20232_ (.A(_03773_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _20233_ (.A0(\rbzero.debug_overlay.vplaneY[-4] ),
    .A1(\rbzero.pov.ready_buffer[5] ),
    .S(_03710_),
    .X(_03774_));
 sky130_fd_sc_hd__or2_1 _20234_ (.A(_04470_),
    .B(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__clkbuf_1 _20235_ (.A(_03775_),
    .X(_01235_));
 sky130_fd_sc_hd__or2_1 _20236_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(_03711_),
    .X(_03776_));
 sky130_fd_sc_hd__o211a_1 _20237_ (.A1(\rbzero.pov.ready_buffer[6] ),
    .A2(_03707_),
    .B1(_03776_),
    .C1(_03765_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _20238_ (.A0(_05177_),
    .A1(\rbzero.pov.ready_buffer[7] ),
    .S(_03710_),
    .X(_03777_));
 sky130_fd_sc_hd__or2_1 _20239_ (.A(_04470_),
    .B(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__clkbuf_1 _20240_ (.A(_03778_),
    .X(_01237_));
 sky130_fd_sc_hd__or2_1 _20241_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_03711_),
    .X(_03779_));
 sky130_fd_sc_hd__o211a_1 _20242_ (.A1(\rbzero.pov.ready_buffer[8] ),
    .A2(_03707_),
    .B1(_03779_),
    .C1(_03765_),
    .X(_01238_));
 sky130_fd_sc_hd__or2_1 _20243_ (.A(_02829_),
    .B(_03711_),
    .X(_03780_));
 sky130_fd_sc_hd__o211a_1 _20244_ (.A1(\rbzero.pov.ready_buffer[9] ),
    .A2(_03707_),
    .B1(_03780_),
    .C1(_03765_),
    .X(_01239_));
 sky130_fd_sc_hd__or2_1 _20245_ (.A(_02858_),
    .B(_03711_),
    .X(_03781_));
 sky130_fd_sc_hd__o211a_1 _20246_ (.A1(\rbzero.pov.ready_buffer[10] ),
    .A2(_03707_),
    .B1(_03781_),
    .C1(_03765_),
    .X(_01240_));
 sky130_fd_sc_hd__a31o_1 _20247_ (.A1(_03486_),
    .A2(_03485_),
    .A3(_03491_),
    .B1(\rbzero.pov.spi_done ),
    .X(_03782_));
 sky130_fd_sc_hd__and2_1 _20248_ (.A(_03006_),
    .B(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_1 _20249_ (.A(_03783_),
    .X(_01241_));
 sky130_fd_sc_hd__nand3b_1 _20250_ (.A_N(_05758_),
    .B(_05099_),
    .C(_03133_),
    .Y(_03784_));
 sky130_fd_sc_hd__or4bb_1 _20251_ (.A(_04744_),
    .B(_05760_),
    .C_N(_05753_),
    .D_N(_05752_),
    .X(_03785_));
 sky130_fd_sc_hd__or4b_1 _20252_ (.A(_05752_),
    .B(_04745_),
    .C(_05760_),
    .D_N(_05753_),
    .X(_03786_));
 sky130_fd_sc_hd__o21ai_1 _20253_ (.A1(_03784_),
    .A2(_03786_),
    .B1(_04488_),
    .Y(_03787_));
 sky130_fd_sc_hd__o211a_1 _20254_ (.A1(_03784_),
    .A2(_03785_),
    .B1(_03787_),
    .C1(_03765_),
    .X(_01242_));
 sky130_fd_sc_hd__clkinv_2 _20255_ (.A(_04510_),
    .Y(_03788_));
 sky130_fd_sc_hd__and4_1 _20256_ (.A(_04476_),
    .B(_04643_),
    .C(_04035_),
    .D(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__or4b_1 _20257_ (.A(_04501_),
    .B(_04481_),
    .C(_05105_),
    .D_N(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__a41o_1 _20258_ (.A1(_04032_),
    .A2(_04481_),
    .A3(_05105_),
    .A4(_03789_),
    .B1(_04470_),
    .X(_03791_));
 sky130_fd_sc_hd__a21oi_1 _20259_ (.A1(_05713_),
    .A2(_03790_),
    .B1(_03791_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_1 _20260_ (.A(_05762_),
    .B(_04700_),
    .Y(_03792_));
 sky130_fd_sc_hd__or4_1 _20261_ (.A(_05761_),
    .B(_04758_),
    .C(_03785_),
    .D(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__and2_1 _20262_ (.A(_09805_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__nand2_1 _20263_ (.A(_05760_),
    .B(_09805_),
    .Y(_03795_));
 sky130_fd_sc_hd__o211a_1 _20264_ (.A1(_05760_),
    .A2(_03794_),
    .B1(_03795_),
    .C1(_03159_),
    .X(_01244_));
 sky130_fd_sc_hd__nor2_1 _20265_ (.A(_04745_),
    .B(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__a211oi_1 _20266_ (.A1(_04745_),
    .A2(_03795_),
    .B1(_03796_),
    .C1(_03322_),
    .Y(_01245_));
 sky130_fd_sc_hd__a21o_1 _20267_ (.A1(_04112_),
    .A2(_03793_),
    .B1(_09816_),
    .X(_03797_));
 sky130_fd_sc_hd__o211a_1 _20268_ (.A1(_05752_),
    .A2(_03796_),
    .B1(_03797_),
    .C1(_03131_),
    .X(_01246_));
 sky130_fd_sc_hd__clkbuf_4 _20269_ (.A(_09816_),
    .X(_03798_));
 sky130_fd_sc_hd__a21oi_1 _20270_ (.A1(_05753_),
    .A2(_03130_),
    .B1(_04469_),
    .Y(_03799_));
 sky130_fd_sc_hd__o21a_1 _20271_ (.A1(_05753_),
    .A2(_03130_),
    .B1(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__a22o_1 _20272_ (.A1(_05753_),
    .A2(_03798_),
    .B1(_03794_),
    .B2(_03800_),
    .X(_01247_));
 sky130_fd_sc_hd__and3_1 _20273_ (.A(_05753_),
    .B(_05752_),
    .C(_03796_),
    .X(_03801_));
 sky130_fd_sc_hd__o221a_1 _20274_ (.A1(_04703_),
    .A2(_03131_),
    .B1(_03801_),
    .B2(_05758_),
    .C1(_03159_),
    .X(_01248_));
 sky130_fd_sc_hd__and3_1 _20275_ (.A(_04704_),
    .B(_05758_),
    .C(_03138_),
    .X(_03802_));
 sky130_fd_sc_hd__inv_2 _20276_ (.A(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__o211a_1 _20277_ (.A1(_04704_),
    .A2(_03132_),
    .B1(_03803_),
    .C1(_03159_),
    .X(_01249_));
 sky130_fd_sc_hd__o21ai_1 _20278_ (.A1(_05755_),
    .A2(_03802_),
    .B1(_08186_),
    .Y(_03804_));
 sky130_fd_sc_hd__nor2_1 _20279_ (.A(_04770_),
    .B(_03803_),
    .Y(_03805_));
 sky130_fd_sc_hd__nor2_1 _20280_ (.A(_03804_),
    .B(_03805_),
    .Y(_01250_));
 sky130_fd_sc_hd__and3_1 _20281_ (.A(_04704_),
    .B(_05758_),
    .C(_03801_),
    .X(_03806_));
 sky130_fd_sc_hd__a31o_1 _20282_ (.A1(_05756_),
    .A2(_05755_),
    .A3(_03806_),
    .B1(_04470_),
    .X(_03807_));
 sky130_fd_sc_hd__o21ba_1 _20283_ (.A1(_05756_),
    .A2(_03805_),
    .B1_N(_03807_),
    .X(_01251_));
 sky130_fd_sc_hd__and4_1 _20284_ (.A(_05761_),
    .B(_05756_),
    .C(_05755_),
    .D(_03806_),
    .X(_03808_));
 sky130_fd_sc_hd__a31o_1 _20285_ (.A1(_05756_),
    .A2(_05755_),
    .A3(_03802_),
    .B1(_05761_),
    .X(_03809_));
 sky130_fd_sc_hd__and3b_1 _20286_ (.A_N(_03808_),
    .B(_08185_),
    .C(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _20287_ (.A(_03810_),
    .X(_01252_));
 sky130_fd_sc_hd__a21boi_1 _20288_ (.A1(_05762_),
    .A2(_03808_),
    .B1_N(_03797_),
    .Y(_03811_));
 sky130_fd_sc_hd__o21a_1 _20289_ (.A1(_05762_),
    .A2(_03808_),
    .B1(_03811_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _20290_ (.A0(\rbzero.spi_registers.new_texadd[3][0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03430_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_1 _20291_ (.A(_03812_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _20292_ (.A0(\rbzero.spi_registers.new_texadd[3][1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_03430_),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_1 _20293_ (.A(_03813_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _20294_ (.A0(\rbzero.spi_registers.new_texadd[3][2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_03430_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_1 _20295_ (.A(_03814_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _20296_ (.A0(\rbzero.spi_registers.new_texadd[3][3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_03430_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _20297_ (.A(_03815_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _20298_ (.A0(\rbzero.spi_registers.new_texadd[3][4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_03430_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _20299_ (.A(_03816_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _20300_ (.A0(\rbzero.spi_registers.new_texadd[3][5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_03430_),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_1 _20301_ (.A(_03817_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _20302_ (.A0(\rbzero.spi_registers.new_texadd[3][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03430_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _20303_ (.A(_03818_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _20304_ (.A0(\rbzero.spi_registers.new_texadd[3][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03430_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_1 _20305_ (.A(_03819_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _20306_ (.A0(\rbzero.spi_registers.new_texadd[3][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03430_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_1 _20307_ (.A(_03820_),
    .X(_01262_));
 sky130_fd_sc_hd__buf_4 _20308_ (.A(_03429_),
    .X(_03821_));
 sky130_fd_sc_hd__mux2_1 _20309_ (.A0(\rbzero.spi_registers.new_texadd[3][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _20310_ (.A(_03822_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _20311_ (.A0(\rbzero.spi_registers.new_texadd[3][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03821_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_1 _20312_ (.A(_03823_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _20313_ (.A0(\rbzero.spi_registers.new_texadd[3][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03821_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _20314_ (.A(_03824_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _20315_ (.A0(\rbzero.spi_registers.new_texadd[3][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03821_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_1 _20316_ (.A(_03825_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _20317_ (.A0(\rbzero.spi_registers.new_texadd[3][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03821_),
    .X(_03826_));
 sky130_fd_sc_hd__clkbuf_1 _20318_ (.A(_03826_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _20319_ (.A0(\rbzero.spi_registers.new_texadd[3][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03821_),
    .X(_03827_));
 sky130_fd_sc_hd__clkbuf_1 _20320_ (.A(_03827_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _20321_ (.A0(\rbzero.spi_registers.new_texadd[3][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03821_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_1 _20322_ (.A(_03828_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _20323_ (.A0(\rbzero.spi_registers.new_texadd[3][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03821_),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_1 _20324_ (.A(_03829_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _20325_ (.A0(\rbzero.spi_registers.new_texadd[3][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03821_),
    .X(_03830_));
 sky130_fd_sc_hd__clkbuf_1 _20326_ (.A(_03830_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _20327_ (.A0(\rbzero.spi_registers.new_texadd[3][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03821_),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _20328_ (.A(_03831_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _20329_ (.A0(\rbzero.spi_registers.new_texadd[3][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03429_),
    .X(_03832_));
 sky130_fd_sc_hd__clkbuf_1 _20330_ (.A(_03832_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _20331_ (.A0(\rbzero.spi_registers.new_texadd[3][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03429_),
    .X(_03833_));
 sky130_fd_sc_hd__clkbuf_1 _20332_ (.A(_03833_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _20333_ (.A0(\rbzero.spi_registers.new_texadd[3][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03429_),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _20334_ (.A(_03834_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _20335_ (.A0(\rbzero.spi_registers.new_texadd[3][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03429_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_1 _20336_ (.A(_03835_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _20337_ (.A0(\rbzero.spi_registers.new_texadd[3][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03429_),
    .X(_03836_));
 sky130_fd_sc_hd__clkbuf_1 _20338_ (.A(_03836_),
    .X(_01277_));
 sky130_fd_sc_hd__inv_2 _20340__93 (.A(clknet_1_0__leaf__03511_),
    .Y(net218));
 sky130_fd_sc_hd__inv_2 _20341__94 (.A(clknet_1_0__leaf__03511_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _20342__95 (.A(clknet_1_0__leaf__03511_),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _20343__96 (.A(clknet_1_1__leaf__03511_),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _20344__97 (.A(clknet_1_1__leaf__03511_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _20346__98 (.A(clknet_1_0__leaf__03837_),
    .Y(net223));
 sky130_fd_sc_hd__buf_1 _20345_ (.A(clknet_1_1__leaf__03510_),
    .X(_03837_));
 sky130_fd_sc_hd__inv_2 _20347__99 (.A(clknet_1_0__leaf__03837_),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _20348__100 (.A(clknet_1_1__leaf__03837_),
    .Y(net225));
 sky130_fd_sc_hd__inv_2 _20349__101 (.A(clknet_1_1__leaf__03837_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _20350__102 (.A(clknet_1_1__leaf__03837_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _20351__103 (.A(clknet_1_1__leaf__03837_),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _20352__104 (.A(clknet_1_1__leaf__03837_),
    .Y(net229));
 sky130_fd_sc_hd__inv_2 _20353__105 (.A(clknet_1_0__leaf__03837_),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _20354__106 (.A(clknet_1_0__leaf__03837_),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _20355__107 (.A(clknet_1_0__leaf__03837_),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _20357__108 (.A(clknet_1_0__leaf__03838_),
    .Y(net233));
 sky130_fd_sc_hd__buf_1 _20356_ (.A(clknet_1_1__leaf__03510_),
    .X(_03838_));
 sky130_fd_sc_hd__inv_2 _20358__109 (.A(clknet_1_0__leaf__03838_),
    .Y(net234));
 sky130_fd_sc_hd__inv_2 _20359__110 (.A(clknet_1_0__leaf__03838_),
    .Y(net235));
 sky130_fd_sc_hd__inv_2 _20360__111 (.A(clknet_1_0__leaf__03838_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _20361__112 (.A(clknet_1_0__leaf__03838_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _20362__113 (.A(clknet_1_0__leaf__03838_),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _20363__114 (.A(clknet_1_1__leaf__03838_),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _20364__115 (.A(clknet_1_1__leaf__03838_),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _20365__116 (.A(clknet_1_1__leaf__03838_),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _20366__117 (.A(clknet_1_1__leaf__03838_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _20368__118 (.A(clknet_1_1__leaf__03839_),
    .Y(net243));
 sky130_fd_sc_hd__buf_1 _20367_ (.A(clknet_1_1__leaf__03510_),
    .X(_03839_));
 sky130_fd_sc_hd__inv_2 _20369__119 (.A(clknet_1_1__leaf__03839_),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _20370__120 (.A(clknet_1_1__leaf__03839_),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _20371__121 (.A(clknet_1_1__leaf__03839_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _20372__122 (.A(clknet_1_1__leaf__03839_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _20373__123 (.A(clknet_1_0__leaf__03839_),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _20374__124 (.A(clknet_1_0__leaf__03839_),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _20375__125 (.A(clknet_1_0__leaf__03839_),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _20376__126 (.A(clknet_1_0__leaf__03839_),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _20377__127 (.A(clknet_1_0__leaf__03839_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _20379__128 (.A(clknet_1_1__leaf__03840_),
    .Y(net253));
 sky130_fd_sc_hd__buf_1 _20378_ (.A(clknet_1_1__leaf__03510_),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _20380__129 (.A(clknet_1_1__leaf__03840_),
    .Y(net254));
 sky130_fd_sc_hd__inv_2 _20381__130 (.A(clknet_1_1__leaf__03840_),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _20382__131 (.A(clknet_1_1__leaf__03840_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _20383__132 (.A(clknet_1_1__leaf__03840_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _20384__133 (.A(clknet_1_0__leaf__03840_),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _20385__134 (.A(clknet_1_0__leaf__03840_),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _20386__135 (.A(clknet_1_0__leaf__03840_),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _20387__136 (.A(clknet_1_0__leaf__03840_),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _20388__137 (.A(clknet_1_0__leaf__03840_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _20390__138 (.A(clknet_1_1__leaf__03841_),
    .Y(net263));
 sky130_fd_sc_hd__buf_1 _20389_ (.A(clknet_1_1__leaf__03510_),
    .X(_03841_));
 sky130_fd_sc_hd__inv_2 _20391__139 (.A(clknet_1_1__leaf__03841_),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _20392__140 (.A(clknet_1_0__leaf__03841_),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _20393__141 (.A(clknet_1_0__leaf__03841_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _20394__142 (.A(clknet_1_0__leaf__03841_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _20395__143 (.A(clknet_1_0__leaf__03841_),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _20396__144 (.A(clknet_1_0__leaf__03841_),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _20397__145 (.A(clknet_1_1__leaf__03841_),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _20398__146 (.A(clknet_1_1__leaf__03841_),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _20399__147 (.A(clknet_1_1__leaf__03841_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _20401__148 (.A(clknet_1_1__leaf__03842_),
    .Y(net273));
 sky130_fd_sc_hd__buf_1 _20400_ (.A(clknet_1_0__leaf__03510_),
    .X(_03842_));
 sky130_fd_sc_hd__inv_2 _20402__149 (.A(clknet_1_1__leaf__03842_),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _20403__150 (.A(clknet_1_1__leaf__03842_),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _20404__151 (.A(clknet_1_1__leaf__03842_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _20405__152 (.A(clknet_1_0__leaf__03842_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _20406__153 (.A(clknet_1_0__leaf__03842_),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _20407__154 (.A(clknet_1_0__leaf__03842_),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _20408__155 (.A(clknet_1_0__leaf__03842_),
    .Y(net280));
 sky130_fd_sc_hd__inv_2 _20409__156 (.A(clknet_1_1__leaf__03842_),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _20410__157 (.A(clknet_1_1__leaf__03842_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _20412__158 (.A(clknet_1_1__leaf__03843_),
    .Y(net283));
 sky130_fd_sc_hd__buf_1 _20411_ (.A(clknet_1_0__leaf__03510_),
    .X(_03843_));
 sky130_fd_sc_hd__inv_2 _20413__159 (.A(clknet_1_1__leaf__03843_),
    .Y(net284));
 sky130_fd_sc_hd__inv_2 _20414__160 (.A(clknet_1_1__leaf__03843_),
    .Y(net285));
 sky130_fd_sc_hd__inv_2 _20415__161 (.A(clknet_1_1__leaf__03843_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _20416__162 (.A(clknet_1_0__leaf__03843_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _20417__163 (.A(clknet_1_0__leaf__03843_),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _20418__164 (.A(clknet_1_0__leaf__03843_),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _20419__165 (.A(clknet_1_0__leaf__03843_),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _20420__166 (.A(clknet_1_0__leaf__03843_),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _20421__167 (.A(clknet_1_0__leaf__03843_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _20423__168 (.A(clknet_1_0__leaf__03844_),
    .Y(net293));
 sky130_fd_sc_hd__buf_1 _20422_ (.A(clknet_1_0__leaf__03510_),
    .X(_03844_));
 sky130_fd_sc_hd__inv_2 _20424__169 (.A(clknet_1_1__leaf__03844_),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _20425__170 (.A(clknet_1_1__leaf__03844_),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _20426__171 (.A(clknet_1_1__leaf__03844_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _20427__172 (.A(clknet_1_1__leaf__03844_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _20428__173 (.A(clknet_1_1__leaf__03844_),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _20429__174 (.A(clknet_1_1__leaf__03844_),
    .Y(net299));
 sky130_fd_sc_hd__inv_2 _20430__175 (.A(clknet_1_0__leaf__03844_),
    .Y(net300));
 sky130_fd_sc_hd__inv_2 _20431__176 (.A(clknet_1_0__leaf__03844_),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _20432__177 (.A(clknet_1_0__leaf__03844_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _20434__178 (.A(clknet_1_1__leaf__03845_),
    .Y(net303));
 sky130_fd_sc_hd__buf_1 _20433_ (.A(clknet_1_0__leaf__03510_),
    .X(_03845_));
 sky130_fd_sc_hd__inv_2 _20435__179 (.A(clknet_1_1__leaf__03845_),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _20436__180 (.A(clknet_1_1__leaf__03845_),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _20437__181 (.A(clknet_1_1__leaf__03845_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _20438__182 (.A(clknet_1_1__leaf__03845_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _20439__183 (.A(clknet_1_0__leaf__03845_),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _20440__184 (.A(clknet_1_0__leaf__03845_),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _20441__185 (.A(clknet_1_0__leaf__03845_),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 _20442__186 (.A(clknet_1_0__leaf__03845_),
    .Y(net311));
 sky130_fd_sc_hd__inv_2 _20443__187 (.A(clknet_1_0__leaf__03845_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _20446__188 (.A(clknet_1_1__leaf__03847_),
    .Y(net313));
 sky130_fd_sc_hd__buf_1 _20444_ (.A(clknet_1_1__leaf__05825_),
    .X(_03846_));
 sky130_fd_sc_hd__buf_1 _20445_ (.A(clknet_1_1__leaf__03846_),
    .X(_03847_));
 sky130_fd_sc_hd__inv_2 _20447__189 (.A(clknet_1_1__leaf__03847_),
    .Y(net314));
 sky130_fd_sc_hd__inv_2 _20448__190 (.A(clknet_1_1__leaf__03847_),
    .Y(net315));
 sky130_fd_sc_hd__inv_2 _20449__191 (.A(clknet_1_1__leaf__03847_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _20450__192 (.A(clknet_1_1__leaf__03847_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _20451__193 (.A(clknet_1_1__leaf__03847_),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _20452__194 (.A(clknet_1_0__leaf__03847_),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 _20453__195 (.A(clknet_1_0__leaf__03847_),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _20454__196 (.A(clknet_1_0__leaf__03847_),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _20455__197 (.A(clknet_1_0__leaf__03847_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _20457__198 (.A(clknet_1_1__leaf__03848_),
    .Y(net323));
 sky130_fd_sc_hd__buf_1 _20456_ (.A(clknet_1_1__leaf__03846_),
    .X(_03848_));
 sky130_fd_sc_hd__inv_2 _20458__199 (.A(clknet_1_1__leaf__03848_),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _20459__200 (.A(clknet_1_1__leaf__03848_),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _20460__201 (.A(clknet_1_1__leaf__03848_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _20461__202 (.A(clknet_1_1__leaf__03848_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _20462__203 (.A(clknet_1_1__leaf__03848_),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _20463__204 (.A(clknet_1_0__leaf__03848_),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _20464__205 (.A(clknet_1_0__leaf__03848_),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _20465__206 (.A(clknet_1_0__leaf__03848_),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _20466__207 (.A(clknet_1_0__leaf__03848_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _20468__208 (.A(clknet_1_1__leaf__03849_),
    .Y(net333));
 sky130_fd_sc_hd__buf_1 _20467_ (.A(clknet_1_1__leaf__03846_),
    .X(_03849_));
 sky130_fd_sc_hd__inv_2 _20469__209 (.A(clknet_1_1__leaf__03849_),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _20470__210 (.A(clknet_1_1__leaf__03849_),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _20471__211 (.A(clknet_1_1__leaf__03849_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _20472__212 (.A(clknet_1_0__leaf__03849_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _20473__213 (.A(clknet_1_0__leaf__03849_),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _20474__214 (.A(clknet_1_0__leaf__03849_),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _20475__215 (.A(clknet_1_0__leaf__03849_),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _20476__216 (.A(clknet_1_0__leaf__03849_),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _20477__217 (.A(clknet_1_0__leaf__03849_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _20479__218 (.A(clknet_1_1__leaf__03850_),
    .Y(net343));
 sky130_fd_sc_hd__buf_1 _20478_ (.A(clknet_1_1__leaf__03846_),
    .X(_03850_));
 sky130_fd_sc_hd__inv_2 _20480__219 (.A(clknet_1_1__leaf__03850_),
    .Y(net344));
 sky130_fd_sc_hd__inv_2 _20481__220 (.A(clknet_1_0__leaf__03850_),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _20482__221 (.A(clknet_1_1__leaf__03850_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _20483__222 (.A(clknet_1_1__leaf__03850_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _20484__223 (.A(clknet_1_1__leaf__03850_),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _20485__224 (.A(clknet_1_0__leaf__03850_),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _20486__225 (.A(clknet_1_0__leaf__03850_),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _20487__226 (.A(clknet_1_0__leaf__03850_),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _20488__227 (.A(clknet_1_0__leaf__03850_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _20490__228 (.A(clknet_1_1__leaf__03851_),
    .Y(net353));
 sky130_fd_sc_hd__buf_1 _20489_ (.A(clknet_1_0__leaf__03846_),
    .X(_03851_));
 sky130_fd_sc_hd__inv_2 _20491__229 (.A(clknet_1_1__leaf__03851_),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _20492__230 (.A(clknet_1_1__leaf__03851_),
    .Y(net355));
 sky130_fd_sc_hd__inv_2 _20493__231 (.A(clknet_1_1__leaf__03851_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _20494__232 (.A(clknet_1_1__leaf__03851_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _20495__233 (.A(clknet_1_0__leaf__03851_),
    .Y(net358));
 sky130_fd_sc_hd__inv_2 _20496__234 (.A(clknet_1_0__leaf__03851_),
    .Y(net359));
 sky130_fd_sc_hd__inv_2 _20497__235 (.A(clknet_1_0__leaf__03851_),
    .Y(net360));
 sky130_fd_sc_hd__inv_2 _20498__236 (.A(clknet_1_0__leaf__03851_),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 _20499__237 (.A(clknet_1_1__leaf__03851_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _20501__238 (.A(clknet_1_1__leaf__03852_),
    .Y(net363));
 sky130_fd_sc_hd__buf_1 _20500_ (.A(clknet_1_0__leaf__03846_),
    .X(_03852_));
 sky130_fd_sc_hd__inv_2 _20502__239 (.A(clknet_1_1__leaf__03852_),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _20503__240 (.A(clknet_1_1__leaf__03852_),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _20504__241 (.A(clknet_1_1__leaf__03852_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _20505__242 (.A(clknet_1_0__leaf__03852_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _20506__243 (.A(clknet_1_0__leaf__03852_),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _20507__244 (.A(clknet_1_0__leaf__03852_),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _20508__245 (.A(clknet_1_0__leaf__03852_),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _20509__246 (.A(clknet_1_0__leaf__03852_),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _20510__247 (.A(clknet_1_0__leaf__03852_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _20512__248 (.A(clknet_1_0__leaf__03853_),
    .Y(net373));
 sky130_fd_sc_hd__buf_1 _20511_ (.A(clknet_1_0__leaf__03846_),
    .X(_03853_));
 sky130_fd_sc_hd__inv_2 _20513__249 (.A(clknet_1_1__leaf__03853_),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _20514__250 (.A(clknet_1_1__leaf__03853_),
    .Y(net375));
 sky130_fd_sc_hd__inv_2 _20515__251 (.A(clknet_1_1__leaf__03853_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _20516__252 (.A(clknet_1_1__leaf__03853_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _20517__253 (.A(clknet_1_1__leaf__03853_),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _20518__254 (.A(clknet_1_1__leaf__03853_),
    .Y(net379));
 sky130_fd_sc_hd__inv_2 _20519__255 (.A(clknet_1_0__leaf__03853_),
    .Y(net380));
 sky130_fd_sc_hd__inv_2 _20520__256 (.A(clknet_1_0__leaf__03853_),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _20521__257 (.A(clknet_1_0__leaf__03853_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _20523__258 (.A(clknet_1_0__leaf__03854_),
    .Y(net383));
 sky130_fd_sc_hd__buf_1 _20522_ (.A(clknet_1_0__leaf__03846_),
    .X(_03854_));
 sky130_fd_sc_hd__inv_2 _20524__259 (.A(clknet_1_0__leaf__03854_),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _20525__260 (.A(clknet_1_0__leaf__03854_),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _20526__261 (.A(clknet_1_0__leaf__03854_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _20527__262 (.A(clknet_1_0__leaf__03854_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _20528__263 (.A(clknet_1_1__leaf__03854_),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _20529__264 (.A(clknet_1_1__leaf__03854_),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _20530__265 (.A(clknet_1_1__leaf__03854_),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _20531__266 (.A(clknet_1_1__leaf__03854_),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _20532__267 (.A(clknet_1_1__leaf__03854_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _20534__268 (.A(clknet_1_0__leaf__03855_),
    .Y(net393));
 sky130_fd_sc_hd__buf_1 _20533_ (.A(clknet_1_0__leaf__03846_),
    .X(_03855_));
 sky130_fd_sc_hd__inv_2 _20535__269 (.A(clknet_1_0__leaf__03855_),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _20536__270 (.A(clknet_1_1__leaf__03855_),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _20537__271 (.A(clknet_1_1__leaf__03855_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _20538__272 (.A(clknet_1_1__leaf__03855_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _20539__273 (.A(clknet_1_1__leaf__03855_),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _20540__274 (.A(clknet_1_0__leaf__03855_),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _20541__275 (.A(clknet_1_0__leaf__03855_),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _20542__276 (.A(clknet_1_1__leaf__03855_),
    .Y(net401));
 sky130_fd_sc_hd__inv_2 _20543__277 (.A(clknet_1_1__leaf__03855_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _20545__278 (.A(clknet_1_0__leaf__03856_),
    .Y(net403));
 sky130_fd_sc_hd__buf_1 _20544_ (.A(clknet_1_1__leaf__03846_),
    .X(_03856_));
 sky130_fd_sc_hd__inv_2 _20546__279 (.A(clknet_1_0__leaf__03856_),
    .Y(net404));
 sky130_fd_sc_hd__inv_2 _20547__280 (.A(clknet_1_0__leaf__03856_),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _20548__281 (.A(clknet_1_0__leaf__03856_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _20549__282 (.A(clknet_1_1__leaf__03856_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _20550__283 (.A(clknet_1_1__leaf__03856_),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _20551__284 (.A(clknet_1_1__leaf__03856_),
    .Y(net409));
 sky130_fd_sc_hd__inv_2 _20552__285 (.A(clknet_1_1__leaf__03856_),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _20553__286 (.A(clknet_1_1__leaf__03856_),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _20554__287 (.A(clknet_1_1__leaf__03856_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _20557__288 (.A(clknet_1_1__leaf__03858_),
    .Y(net413));
 sky130_fd_sc_hd__buf_1 _20555_ (.A(clknet_1_1__leaf__05825_),
    .X(_03857_));
 sky130_fd_sc_hd__buf_1 _20556_ (.A(clknet_1_1__leaf__03857_),
    .X(_03858_));
 sky130_fd_sc_hd__inv_2 _20558__289 (.A(clknet_1_1__leaf__03858_),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _20559__290 (.A(clknet_1_1__leaf__03858_),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _20560__291 (.A(clknet_1_1__leaf__03858_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _20561__292 (.A(clknet_1_1__leaf__03858_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _20562__293 (.A(clknet_1_1__leaf__03858_),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _20563__294 (.A(clknet_1_0__leaf__03858_),
    .Y(net419));
 sky130_fd_sc_hd__inv_2 _20564__295 (.A(clknet_1_0__leaf__03858_),
    .Y(net420));
 sky130_fd_sc_hd__inv_2 _20565__296 (.A(clknet_1_0__leaf__03858_),
    .Y(net421));
 sky130_fd_sc_hd__inv_2 _20566__297 (.A(clknet_1_0__leaf__03858_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _20568__298 (.A(clknet_1_1__leaf__03859_),
    .Y(net423));
 sky130_fd_sc_hd__buf_1 _20567_ (.A(clknet_1_1__leaf__03857_),
    .X(_03859_));
 sky130_fd_sc_hd__inv_2 _20569__299 (.A(clknet_1_1__leaf__03859_),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _20570__300 (.A(clknet_1_1__leaf__03859_),
    .Y(net425));
 sky130_fd_sc_hd__inv_2 _20571__301 (.A(clknet_1_1__leaf__03859_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _20572__302 (.A(clknet_1_1__leaf__03859_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _20573__303 (.A(clknet_1_1__leaf__03859_),
    .Y(net428));
 sky130_fd_sc_hd__inv_2 _20574__304 (.A(clknet_1_0__leaf__03859_),
    .Y(net429));
 sky130_fd_sc_hd__inv_2 _20575__305 (.A(clknet_1_0__leaf__03859_),
    .Y(net430));
 sky130_fd_sc_hd__inv_2 _20576__306 (.A(clknet_1_0__leaf__03859_),
    .Y(net431));
 sky130_fd_sc_hd__inv_2 _20577__307 (.A(clknet_1_0__leaf__03859_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _20579__308 (.A(clknet_1_1__leaf__03860_),
    .Y(net433));
 sky130_fd_sc_hd__buf_1 _20578_ (.A(clknet_1_1__leaf__03857_),
    .X(_03860_));
 sky130_fd_sc_hd__inv_2 _20580__309 (.A(clknet_1_1__leaf__03860_),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _20581__310 (.A(clknet_1_1__leaf__03860_),
    .Y(net435));
 sky130_fd_sc_hd__inv_2 _20582__311 (.A(clknet_1_1__leaf__03860_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _20583__312 (.A(clknet_1_1__leaf__03860_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _20584__313 (.A(clknet_1_0__leaf__03860_),
    .Y(net438));
 sky130_fd_sc_hd__inv_2 _20585__314 (.A(clknet_1_0__leaf__03860_),
    .Y(net439));
 sky130_fd_sc_hd__inv_2 _20586__315 (.A(clknet_1_0__leaf__03860_),
    .Y(net440));
 sky130_fd_sc_hd__inv_2 _20587__316 (.A(clknet_1_0__leaf__03860_),
    .Y(net441));
 sky130_fd_sc_hd__inv_2 _20588__317 (.A(clknet_1_0__leaf__03860_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _20590__318 (.A(clknet_1_1__leaf__03861_),
    .Y(net443));
 sky130_fd_sc_hd__buf_1 _20589_ (.A(clknet_1_1__leaf__03857_),
    .X(_03861_));
 sky130_fd_sc_hd__inv_2 _20591__319 (.A(clknet_1_1__leaf__03861_),
    .Y(net444));
 sky130_fd_sc_hd__inv_2 _20592__320 (.A(clknet_1_1__leaf__03861_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _20593__321 (.A(clknet_1_1__leaf__03861_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _20594__322 (.A(clknet_1_0__leaf__03861_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _20595__323 (.A(clknet_1_0__leaf__03861_),
    .Y(net448));
 sky130_fd_sc_hd__inv_2 _20596__324 (.A(clknet_1_0__leaf__03861_),
    .Y(net449));
 sky130_fd_sc_hd__inv_2 _20597__325 (.A(clknet_1_0__leaf__03861_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _20598__326 (.A(clknet_1_0__leaf__03861_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _20599__327 (.A(clknet_1_0__leaf__03861_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _20601__328 (.A(clknet_1_0__leaf__03862_),
    .Y(net453));
 sky130_fd_sc_hd__buf_1 _20600_ (.A(clknet_1_1__leaf__03857_),
    .X(_03862_));
 sky130_fd_sc_hd__inv_2 _20602__329 (.A(clknet_1_0__leaf__03862_),
    .Y(net454));
 sky130_fd_sc_hd__inv_2 _20603__330 (.A(clknet_1_0__leaf__03862_),
    .Y(net455));
 sky130_fd_sc_hd__inv_2 _20604__331 (.A(clknet_1_0__leaf__03862_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _20605__332 (.A(clknet_1_0__leaf__03862_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _20606__333 (.A(clknet_1_1__leaf__03862_),
    .Y(net458));
 sky130_fd_sc_hd__inv_2 _20607__334 (.A(clknet_1_1__leaf__03862_),
    .Y(net459));
 sky130_fd_sc_hd__inv_2 _20608__335 (.A(clknet_1_1__leaf__03862_),
    .Y(net460));
 sky130_fd_sc_hd__inv_2 _20609__336 (.A(clknet_1_1__leaf__03862_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _20610__337 (.A(clknet_1_1__leaf__03862_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _20612__338 (.A(clknet_1_0__leaf__03863_),
    .Y(net463));
 sky130_fd_sc_hd__buf_1 _20611_ (.A(clknet_1_1__leaf__03857_),
    .X(_03863_));
 sky130_fd_sc_hd__inv_2 _20613__339 (.A(clknet_1_1__leaf__03863_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _20614__340 (.A(clknet_1_1__leaf__03863_),
    .Y(net465));
 sky130_fd_sc_hd__inv_2 _20615__341 (.A(clknet_1_1__leaf__03863_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _20616__342 (.A(clknet_1_1__leaf__03863_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _20617__343 (.A(clknet_1_1__leaf__03863_),
    .Y(net468));
 sky130_fd_sc_hd__inv_2 _20618__344 (.A(clknet_1_0__leaf__03863_),
    .Y(net469));
 sky130_fd_sc_hd__inv_2 _20619__345 (.A(clknet_1_0__leaf__03863_),
    .Y(net470));
 sky130_fd_sc_hd__inv_2 _20620__346 (.A(clknet_1_0__leaf__03863_),
    .Y(net471));
 sky130_fd_sc_hd__inv_2 _20621__347 (.A(clknet_1_0__leaf__03863_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _20623__348 (.A(clknet_1_1__leaf__03864_),
    .Y(net473));
 sky130_fd_sc_hd__buf_1 _20622_ (.A(clknet_1_0__leaf__03857_),
    .X(_03864_));
 sky130_fd_sc_hd__inv_2 _20624__349 (.A(clknet_1_1__leaf__03864_),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _20625__350 (.A(clknet_1_1__leaf__03864_),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _20626__351 (.A(clknet_1_1__leaf__03864_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _20627__352 (.A(clknet_1_1__leaf__03864_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _20628__353 (.A(clknet_1_0__leaf__03864_),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _20629__354 (.A(clknet_1_0__leaf__03864_),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _20630__355 (.A(clknet_1_0__leaf__03864_),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _20631__356 (.A(clknet_1_0__leaf__03864_),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _20632__357 (.A(clknet_1_0__leaf__03864_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _20634__358 (.A(clknet_1_1__leaf__03865_),
    .Y(net483));
 sky130_fd_sc_hd__buf_1 _20633_ (.A(clknet_1_0__leaf__03857_),
    .X(_03865_));
 sky130_fd_sc_hd__inv_2 _20635__359 (.A(clknet_1_1__leaf__03865_),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _20636__360 (.A(clknet_1_1__leaf__03865_),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _20637__361 (.A(clknet_1_1__leaf__03865_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _20638__362 (.A(clknet_1_1__leaf__03865_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _20639__363 (.A(clknet_1_0__leaf__03865_),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _20640__364 (.A(clknet_1_0__leaf__03865_),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _20641__365 (.A(clknet_1_0__leaf__03865_),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _20642__366 (.A(clknet_1_0__leaf__03865_),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _20643__367 (.A(clknet_1_0__leaf__03865_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _20645__368 (.A(clknet_1_1__leaf__03866_),
    .Y(net493));
 sky130_fd_sc_hd__buf_1 _20644_ (.A(clknet_1_0__leaf__03857_),
    .X(_03866_));
 sky130_fd_sc_hd__inv_2 _20646__369 (.A(clknet_1_1__leaf__03866_),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _20647__370 (.A(clknet_1_1__leaf__03866_),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _20648__371 (.A(clknet_1_1__leaf__03866_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _20649__372 (.A(clknet_1_1__leaf__03866_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _20650__373 (.A(clknet_1_0__leaf__03866_),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _20651__374 (.A(clknet_1_0__leaf__03866_),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _20652__375 (.A(clknet_1_0__leaf__03866_),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _20653__376 (.A(clknet_1_0__leaf__03866_),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _20654__377 (.A(clknet_1_0__leaf__03866_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _20656__378 (.A(clknet_1_0__leaf__03867_),
    .Y(net503));
 sky130_fd_sc_hd__buf_1 _20655_ (.A(clknet_1_0__leaf__03857_),
    .X(_03867_));
 sky130_fd_sc_hd__inv_2 _20657__379 (.A(clknet_1_0__leaf__03867_),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _20658__380 (.A(clknet_1_0__leaf__03867_),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _20659__381 (.A(clknet_1_0__leaf__03867_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _20660__382 (.A(clknet_1_0__leaf__03867_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _20661__383 (.A(clknet_1_0__leaf__03867_),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _20662__384 (.A(clknet_1_1__leaf__03867_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _20663__385 (.A(clknet_1_1__leaf__03867_),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _20664__386 (.A(clknet_1_1__leaf__03867_),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _20665__387 (.A(clknet_1_1__leaf__03867_),
    .Y(net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__buf_1 _20666_ (.A(clknet_1_1__leaf__05825_),
    .X(_03868_));
 sky130_fd_sc_hd__inv_2 _20668__9 (.A(clknet_1_0__leaf__03868_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _20669__10 (.A(clknet_1_0__leaf__03868_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _20670__11 (.A(clknet_1_0__leaf__03868_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _20671__12 (.A(clknet_1_1__leaf__03868_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _20672__13 (.A(clknet_1_1__leaf__03868_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _20673__14 (.A(clknet_1_0__leaf__03868_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _20674__15 (.A(clknet_1_1__leaf__03868_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _20675__16 (.A(clknet_1_1__leaf__03868_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _20676__17 (.A(clknet_1_1__leaf__03868_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _20678__18 (.A(clknet_1_0__leaf__03869_),
    .Y(net143));
 sky130_fd_sc_hd__buf_1 _20677_ (.A(clknet_1_1__leaf__05825_),
    .X(_03869_));
 sky130_fd_sc_hd__inv_2 _20679__19 (.A(clknet_1_0__leaf__03869_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _20680__20 (.A(clknet_1_0__leaf__03869_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _20681__21 (.A(clknet_1_0__leaf__03869_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _20682__22 (.A(clknet_1_0__leaf__03869_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _20683__23 (.A(clknet_1_1__leaf__03869_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _20684__24 (.A(clknet_1_1__leaf__03869_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _20685__25 (.A(clknet_1_1__leaf__03869_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _20686__26 (.A(clknet_1_1__leaf__03869_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _20687__27 (.A(clknet_1_1__leaf__03869_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _19751__28 (.A(clknet_1_0__leaf__03504_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _20689__5 (.A(clknet_1_0__leaf__03503_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _20690__6 (.A(clknet_1_0__leaf__03503_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _20691__7 (.A(clknet_1_0__leaf__03503_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _20667__8 (.A(clknet_1_0__leaf__03868_),
    .Y(net133));
 sky130_fd_sc_hd__nor2_1 _20692_ (.A(\gpout5.clk_div[0] ),
    .B(net64),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_1 _20693_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .Y(_03870_));
 sky130_fd_sc_hd__or2_1 _20694_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .X(_03871_));
 sky130_fd_sc_hd__and3_1 _20695_ (.A(_09810_),
    .B(_03870_),
    .C(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__clkbuf_1 _20696_ (.A(_03872_),
    .X(_01599_));
 sky130_fd_sc_hd__nand2_1 _20697_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .Y(_03873_));
 sky130_fd_sc_hd__or2_1 _20698_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .X(_03874_));
 sky130_fd_sc_hd__clkbuf_4 _20699_ (.A(_03122_),
    .X(_03875_));
 sky130_fd_sc_hd__a32o_1 _20700_ (.A1(_03798_),
    .A2(_03873_),
    .A3(_03874_),
    .B1(_03875_),
    .B2(\rbzero.texV[-11] ),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _20701_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .X(_03876_));
 sky130_fd_sc_hd__nand2_1 _20702_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03877_));
 sky130_fd_sc_hd__nand3b_1 _20703_ (.A_N(_03873_),
    .B(_03876_),
    .C(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__a21bo_1 _20704_ (.A1(_03876_),
    .A2(_03877_),
    .B1_N(_03873_),
    .X(_03879_));
 sky130_fd_sc_hd__a32o_1 _20705_ (.A1(_03798_),
    .A2(_03878_),
    .A3(_03879_),
    .B1(_03875_),
    .B2(\rbzero.texV[-10] ),
    .X(_01601_));
 sky130_fd_sc_hd__clkbuf_4 _20706_ (.A(_09816_),
    .X(_03880_));
 sky130_fd_sc_hd__and2_1 _20707_ (.A(_03877_),
    .B(_03878_),
    .X(_03881_));
 sky130_fd_sc_hd__nor2_1 _20708_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _20709_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03883_));
 sky130_fd_sc_hd__and2b_1 _20710_ (.A_N(_03882_),
    .B(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__xnor2_1 _20711_ (.A(_03881_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__a22o_1 _20712_ (.A1(\rbzero.texV[-9] ),
    .A2(_09813_),
    .B1(_03880_),
    .B2(_03885_),
    .X(_01602_));
 sky130_fd_sc_hd__or2_1 _20713_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .X(_03886_));
 sky130_fd_sc_hd__nand2_1 _20714_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_03887_));
 sky130_fd_sc_hd__nand2_1 _20715_ (.A(_03886_),
    .B(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__o21ai_1 _20716_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03883_),
    .Y(_03889_));
 sky130_fd_sc_hd__xnor2_1 _20717_ (.A(_03888_),
    .B(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__a22o_1 _20718_ (.A1(\rbzero.texV[-8] ),
    .A2(_09813_),
    .B1(_03880_),
    .B2(_03890_),
    .X(_01603_));
 sky130_fd_sc_hd__nor2_1 _20719_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .Y(_03891_));
 sky130_fd_sc_hd__and2_1 _20720_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .X(_03892_));
 sky130_fd_sc_hd__a21boi_1 _20721_ (.A1(_03886_),
    .A2(_03889_),
    .B1_N(_03887_),
    .Y(_03893_));
 sky130_fd_sc_hd__o21ai_1 _20722_ (.A1(_03891_),
    .A2(_03892_),
    .B1(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__or3_1 _20723_ (.A(_03891_),
    .B(_03892_),
    .C(_03893_),
    .X(_03895_));
 sky130_fd_sc_hd__a32o_1 _20724_ (.A1(_03798_),
    .A2(_03894_),
    .A3(_03895_),
    .B1(_03875_),
    .B2(\rbzero.texV[-7] ),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_1 _20725_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_03896_));
 sky130_fd_sc_hd__o21bai_1 _20726_ (.A1(_03891_),
    .A2(_03893_),
    .B1_N(_03892_),
    .Y(_03897_));
 sky130_fd_sc_hd__xnor2_1 _20727_ (.A(_03896_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__a22o_1 _20728_ (.A1(\rbzero.texV[-6] ),
    .A2(_09813_),
    .B1(_03880_),
    .B2(_03898_),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _20729_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_03899_));
 sky130_fd_sc_hd__and2_1 _20730_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .X(_03900_));
 sky130_fd_sc_hd__a21o_1 _20731_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_03897_),
    .X(_03901_));
 sky130_fd_sc_hd__o21ai_1 _20732_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__or3_1 _20733_ (.A(_03899_),
    .B(_03900_),
    .C(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__o21ai_1 _20734_ (.A1(_03899_),
    .A2(_03900_),
    .B1(_03902_),
    .Y(_03904_));
 sky130_fd_sc_hd__a32o_1 _20735_ (.A1(_03798_),
    .A2(_03903_),
    .A3(_03904_),
    .B1(_03875_),
    .B2(\rbzero.texV[-5] ),
    .X(_01606_));
 sky130_fd_sc_hd__xnor2_1 _20736_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_03905_));
 sky130_fd_sc_hd__o21bai_1 _20737_ (.A1(_03899_),
    .A2(_03902_),
    .B1_N(_03900_),
    .Y(_03906_));
 sky130_fd_sc_hd__xnor2_1 _20738_ (.A(_03905_),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__a22o_1 _20739_ (.A1(\rbzero.texV[-4] ),
    .A2(_09813_),
    .B1(_03880_),
    .B2(_03907_),
    .X(_01607_));
 sky130_fd_sc_hd__nor2_1 _20740_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03908_));
 sky130_fd_sc_hd__nand2_1 _20741_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03909_));
 sky130_fd_sc_hd__and2b_1 _20742_ (.A_N(_03908_),
    .B(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__a21o_1 _20743_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_03906_),
    .X(_03911_));
 sky130_fd_sc_hd__o21ai_1 _20744_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__xnor2_1 _20745_ (.A(_03910_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__a22o_1 _20746_ (.A1(\rbzero.texV[-3] ),
    .A2(_03875_),
    .B1(_03880_),
    .B2(_03913_),
    .X(_01608_));
 sky130_fd_sc_hd__or2_1 _20747_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .X(_03914_));
 sky130_fd_sc_hd__nand2_1 _20748_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .Y(_03915_));
 sky130_fd_sc_hd__o21ai_1 _20749_ (.A1(_03908_),
    .A2(_03912_),
    .B1(_03909_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand3_1 _20750_ (.A(_03914_),
    .B(_03915_),
    .C(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__a21o_1 _20751_ (.A1(_03914_),
    .A2(_03915_),
    .B1(_03916_),
    .X(_03918_));
 sky130_fd_sc_hd__a32o_1 _20752_ (.A1(_03798_),
    .A2(_03917_),
    .A3(_03918_),
    .B1(_03613_),
    .B2(\rbzero.texV[-2] ),
    .X(_01609_));
 sky130_fd_sc_hd__nor2_1 _20753_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .Y(_03919_));
 sky130_fd_sc_hd__and2_1 _20754_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .X(_03920_));
 sky130_fd_sc_hd__or2_1 _20755_ (.A(_03919_),
    .B(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__a21boi_1 _20756_ (.A1(_03914_),
    .A2(_03916_),
    .B1_N(_03915_),
    .Y(_03922_));
 sky130_fd_sc_hd__xor2_1 _20757_ (.A(_03921_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__a22o_1 _20758_ (.A1(\rbzero.texV[-1] ),
    .A2(_03875_),
    .B1(_03880_),
    .B2(_03923_),
    .X(_01610_));
 sky130_fd_sc_hd__or2_1 _20759_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .X(_03924_));
 sky130_fd_sc_hd__nand2_1 _20760_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .Y(_03925_));
 sky130_fd_sc_hd__nor2_1 _20761_ (.A(_03921_),
    .B(_03922_),
    .Y(_03926_));
 sky130_fd_sc_hd__a211o_1 _20762_ (.A1(_03924_),
    .A2(_03925_),
    .B1(_03920_),
    .C1(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__o211a_1 _20763_ (.A1(_03920_),
    .A2(_03926_),
    .B1(_03924_),
    .C1(_03925_),
    .X(_03928_));
 sky130_fd_sc_hd__inv_2 _20764_ (.A(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__a32o_1 _20765_ (.A1(_03798_),
    .A2(_03927_),
    .A3(_03929_),
    .B1(_03613_),
    .B2(\rbzero.texV[0] ),
    .X(_01611_));
 sky130_fd_sc_hd__or2_1 _20766_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_1 _20767_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _20768_ (.A(_03925_),
    .B(_03929_),
    .Y(_03932_));
 sky130_fd_sc_hd__and3_1 _20769_ (.A(_03930_),
    .B(_03931_),
    .C(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__inv_2 _20770_ (.A(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__a21o_1 _20771_ (.A1(_03930_),
    .A2(_03931_),
    .B1(_03932_),
    .X(_03935_));
 sky130_fd_sc_hd__a32o_1 _20772_ (.A1(_03798_),
    .A2(_03934_),
    .A3(_03935_),
    .B1(_03613_),
    .B2(\rbzero.texV[1] ),
    .X(_01612_));
 sky130_fd_sc_hd__or2_1 _20773_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .X(_03936_));
 sky130_fd_sc_hd__nand2_1 _20774_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _20775_ (.A(_03931_),
    .B(_03934_),
    .Y(_03938_));
 sky130_fd_sc_hd__a21o_1 _20776_ (.A1(_03936_),
    .A2(_03937_),
    .B1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__and3_1 _20777_ (.A(_03936_),
    .B(_03937_),
    .C(_03938_),
    .X(_03940_));
 sky130_fd_sc_hd__inv_2 _20778_ (.A(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__a32o_1 _20779_ (.A1(_03798_),
    .A2(_03939_),
    .A3(_03941_),
    .B1(_03613_),
    .B2(\rbzero.texV[2] ),
    .X(_01613_));
 sky130_fd_sc_hd__or2_1 _20780_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .X(_03942_));
 sky130_fd_sc_hd__nand2_1 _20781_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _20782_ (.A(_03937_),
    .B(_03941_),
    .Y(_03944_));
 sky130_fd_sc_hd__and3_1 _20783_ (.A(_03942_),
    .B(_03943_),
    .C(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__inv_2 _20784_ (.A(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__a21o_1 _20785_ (.A1(_03942_),
    .A2(_03943_),
    .B1(_03944_),
    .X(_03947_));
 sky130_fd_sc_hd__a32o_1 _20786_ (.A1(_03798_),
    .A2(_03946_),
    .A3(_03947_),
    .B1(_03613_),
    .B2(\rbzero.texV[3] ),
    .X(_01614_));
 sky130_fd_sc_hd__or2_1 _20787_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .X(_03948_));
 sky130_fd_sc_hd__nand2_1 _20788_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_1 _20789_ (.A(_03943_),
    .B(_03946_),
    .Y(_03950_));
 sky130_fd_sc_hd__a21o_1 _20790_ (.A1(_03948_),
    .A2(_03949_),
    .B1(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__nand3_1 _20791_ (.A(_03948_),
    .B(_03949_),
    .C(_03950_),
    .Y(_03952_));
 sky130_fd_sc_hd__a32o_1 _20792_ (.A1(_09816_),
    .A2(_03951_),
    .A3(_03952_),
    .B1(_03613_),
    .B2(\rbzero.texV[4] ),
    .X(_01615_));
 sky130_fd_sc_hd__a21boi_1 _20793_ (.A1(_03948_),
    .A2(_03950_),
    .B1_N(_03949_),
    .Y(_03953_));
 sky130_fd_sc_hd__nor2_1 _20794_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03954_));
 sky130_fd_sc_hd__nand2_1 _20795_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03955_));
 sky130_fd_sc_hd__and2b_1 _20796_ (.A_N(_03954_),
    .B(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__xnor2_1 _20797_ (.A(_03953_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__a22o_1 _20798_ (.A1(\rbzero.texV[5] ),
    .A2(_03875_),
    .B1(_03880_),
    .B2(_03957_),
    .X(_01616_));
 sky130_fd_sc_hd__or2_1 _20799_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .X(_03958_));
 sky130_fd_sc_hd__nand2_1 _20800_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_03959_));
 sky130_fd_sc_hd__nand2_1 _20801_ (.A(_03958_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__o21ai_1 _20802_ (.A1(_03953_),
    .A2(_03954_),
    .B1(_03955_),
    .Y(_03961_));
 sky130_fd_sc_hd__xnor2_1 _20803_ (.A(_03960_),
    .B(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__a22o_1 _20804_ (.A1(\rbzero.texV[6] ),
    .A2(_03875_),
    .B1(_03880_),
    .B2(_03962_),
    .X(_01617_));
 sky130_fd_sc_hd__nor2_1 _20805_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03963_));
 sky130_fd_sc_hd__nand2_1 _20806_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03964_));
 sky130_fd_sc_hd__and2b_1 _20807_ (.A_N(_03963_),
    .B(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__a21boi_1 _20808_ (.A1(_03958_),
    .A2(_03961_),
    .B1_N(_03959_),
    .Y(_03966_));
 sky130_fd_sc_hd__xnor2_1 _20809_ (.A(_03965_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__a22o_1 _20810_ (.A1(\rbzero.texV[7] ),
    .A2(_03875_),
    .B1(_03880_),
    .B2(_03967_),
    .X(_01618_));
 sky130_fd_sc_hd__or2_1 _20811_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .X(_03968_));
 sky130_fd_sc_hd__nand2_1 _20812_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_03969_));
 sky130_fd_sc_hd__o21ai_1 _20813_ (.A1(_03963_),
    .A2(_03966_),
    .B1(_03964_),
    .Y(_03970_));
 sky130_fd_sc_hd__a21o_1 _20814_ (.A1(_03968_),
    .A2(_03969_),
    .B1(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__nand3_1 _20815_ (.A(_03968_),
    .B(_03969_),
    .C(_03970_),
    .Y(_03972_));
 sky130_fd_sc_hd__a32o_1 _20816_ (.A1(_09816_),
    .A2(_03971_),
    .A3(_03972_),
    .B1(_03613_),
    .B2(\rbzero.texV[8] ),
    .X(_01619_));
 sky130_fd_sc_hd__or2_1 _20817_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .X(_03973_));
 sky130_fd_sc_hd__nand2_1 _20818_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_03974_));
 sky130_fd_sc_hd__a21o_1 _20819_ (.A1(\rbzero.traced_texa[8] ),
    .A2(\rbzero.texV[8] ),
    .B1(_03970_),
    .X(_03975_));
 sky130_fd_sc_hd__nand4_1 _20820_ (.A(_03968_),
    .B(_03973_),
    .C(_03974_),
    .D(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__a22o_1 _20821_ (.A1(_03973_),
    .A2(_03974_),
    .B1(_03975_),
    .B2(_03968_),
    .X(_03977_));
 sky130_fd_sc_hd__a32o_1 _20822_ (.A1(_09816_),
    .A2(_03976_),
    .A3(_03977_),
    .B1(_03613_),
    .B2(\rbzero.texV[9] ),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_1 _20823_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_03978_));
 sky130_fd_sc_hd__and3_1 _20824_ (.A(_03974_),
    .B(_03976_),
    .C(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__a21oi_1 _20825_ (.A1(_03974_),
    .A2(_03976_),
    .B1(_03978_),
    .Y(_03980_));
 sky130_fd_sc_hd__nor2_1 _20826_ (.A(_03979_),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__a22o_1 _20827_ (.A1(\rbzero.texV[10] ),
    .A2(_03875_),
    .B1(_03880_),
    .B2(_03981_),
    .X(_01621_));
 sky130_fd_sc_hd__o21ai_1 _20828_ (.A1(_04493_),
    .A2(_08207_),
    .B1(_04495_),
    .Y(_03982_));
 sky130_fd_sc_hd__nand2_1 _20829_ (.A(_04495_),
    .B(_09805_),
    .Y(_03983_));
 sky130_fd_sc_hd__a21o_1 _20830_ (.A1(_05095_),
    .A2(_03983_),
    .B1(_06331_),
    .X(_03984_));
 sky130_fd_sc_hd__mux2_1 _20831_ (.A0(_03982_),
    .A1(_04495_),
    .S(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__and2_1 _20832_ (.A(_08128_),
    .B(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__clkbuf_1 _20833_ (.A(_03986_),
    .X(_01622_));
 sky130_fd_sc_hd__nand2_1 _20834_ (.A(_04493_),
    .B(_04495_),
    .Y(_03987_));
 sky130_fd_sc_hd__o211a_1 _20835_ (.A1(_03987_),
    .A2(_03984_),
    .B1(_04500_),
    .C1(_04487_),
    .X(_01623_));
 sky130_fd_sc_hd__nor2_1 _20836_ (.A(_03987_),
    .B(_03984_),
    .Y(_03988_));
 sky130_fd_sc_hd__a21oi_1 _20837_ (.A1(_04486_),
    .A2(_03988_),
    .B1(_08201_),
    .Y(_03989_));
 sky130_fd_sc_hd__o21a_1 _20838_ (.A1(_04486_),
    .A2(_03988_),
    .B1(_03989_),
    .X(_01624_));
 sky130_fd_sc_hd__a21boi_1 _20839_ (.A1(_04486_),
    .A2(_04493_),
    .B1_N(\rbzero.trace_state[3] ),
    .Y(_03990_));
 sky130_fd_sc_hd__o31a_1 _20840_ (.A1(_08304_),
    .A2(_03984_),
    .A3(_03990_),
    .B1(_01633_),
    .X(_01625_));
 sky130_fd_sc_hd__and2_2 _20841_ (.A(_08190_),
    .B(clknet_1_0__leaf__05775_),
    .X(_03991_));
 sky130_fd_sc_hd__buf_1 _20842_ (.A(_03991_),
    .X(_01626_));
 sky130_fd_sc_hd__and2_2 _20843_ (.A(_08190_),
    .B(clknet_1_0__leaf__05832_),
    .X(_03992_));
 sky130_fd_sc_hd__buf_1 _20844_ (.A(_03992_),
    .X(_01627_));
 sky130_fd_sc_hd__and2_2 _20845_ (.A(_08190_),
    .B(clknet_1_0__leaf__05887_),
    .X(_03993_));
 sky130_fd_sc_hd__buf_1 _20846_ (.A(_03993_),
    .X(_01628_));
 sky130_fd_sc_hd__and2_2 _20847_ (.A(_09810_),
    .B(clknet_1_1__leaf__05942_),
    .X(_03994_));
 sky130_fd_sc_hd__buf_1 _20848_ (.A(_03994_),
    .X(_01629_));
 sky130_fd_sc_hd__and2_2 _20849_ (.A(_09810_),
    .B(clknet_1_0__leaf__06001_),
    .X(_03995_));
 sky130_fd_sc_hd__buf_1 _20850_ (.A(_03995_),
    .X(_01630_));
 sky130_fd_sc_hd__and2_2 _20851_ (.A(_09810_),
    .B(clknet_1_0__leaf__06050_),
    .X(_03996_));
 sky130_fd_sc_hd__buf_1 _20852_ (.A(_03996_),
    .X(_01631_));
 sky130_fd_sc_hd__nor2_1 _20853_ (.A(\rbzero.hsync ),
    .B(net64),
    .Y(_01632_));
 sky130_fd_sc_hd__a22o_1 _20854_ (.A1(\rbzero.traced_texVinit[0] ),
    .A2(_09836_),
    .B1(_09835_),
    .B2(_09193_),
    .X(_01634_));
 sky130_fd_sc_hd__a22o_1 _20855_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(_09836_),
    .B1(_09835_),
    .B2(_09914_),
    .X(_01635_));
 sky130_fd_sc_hd__inv_2 _20856_ (.A(_09183_),
    .Y(_03997_));
 sky130_fd_sc_hd__a22o_1 _20857_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(_09836_),
    .B1(_09835_),
    .B2(_03997_),
    .X(_01636_));
 sky130_fd_sc_hd__buf_4 _20858_ (.A(_09825_),
    .X(_03998_));
 sky130_fd_sc_hd__a22o_1 _20859_ (.A1(\rbzero.traced_texVinit[3] ),
    .A2(_09836_),
    .B1(_03998_),
    .B2(_09926_),
    .X(_01637_));
 sky130_fd_sc_hd__inv_2 _20860_ (.A(_09422_),
    .Y(_03999_));
 sky130_fd_sc_hd__a22o_1 _20861_ (.A1(\rbzero.traced_texVinit[4] ),
    .A2(_09836_),
    .B1(_03998_),
    .B2(_03999_),
    .X(_01638_));
 sky130_fd_sc_hd__a22o_1 _20862_ (.A1(\rbzero.traced_texVinit[5] ),
    .A2(_09836_),
    .B1(_03998_),
    .B2(_09947_),
    .X(_01639_));
 sky130_fd_sc_hd__a22o_1 _20863_ (.A1(\rbzero.traced_texVinit[6] ),
    .A2(_09836_),
    .B1(_03998_),
    .B2(_09673_),
    .X(_01640_));
 sky130_fd_sc_hd__a22o_1 _20864_ (.A1(\rbzero.traced_texVinit[7] ),
    .A2(_09836_),
    .B1(_03998_),
    .B2(_09797_),
    .X(_01641_));
 sky130_fd_sc_hd__buf_4 _20865_ (.A(_09821_),
    .X(_04000_));
 sky130_fd_sc_hd__a22o_1 _20866_ (.A1(\rbzero.traced_texVinit[8] ),
    .A2(_04000_),
    .B1(_03998_),
    .B2(_10092_),
    .X(_01642_));
 sky130_fd_sc_hd__a22o_1 _20867_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(_04000_),
    .B1(_03998_),
    .B2(_10211_),
    .X(_01643_));
 sky130_fd_sc_hd__a22o_1 _20868_ (.A1(\rbzero.traced_texVinit[10] ),
    .A2(_04000_),
    .B1(_03998_),
    .B2(_10333_),
    .X(_01644_));
 sky130_fd_sc_hd__nor2_1 _20869_ (.A(\gpout0.clk_div[0] ),
    .B(net64),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _20870_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .Y(_04001_));
 sky130_fd_sc_hd__or2_1 _20871_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .X(_04002_));
 sky130_fd_sc_hd__and3_1 _20872_ (.A(_09810_),
    .B(_04001_),
    .C(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__clkbuf_1 _20873_ (.A(_04003_),
    .X(_01646_));
 sky130_fd_sc_hd__or2_1 _20874_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_04004_));
 sky130_fd_sc_hd__and3_1 _20875_ (.A(_09825_),
    .B(_02543_),
    .C(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__a21o_1 _20876_ (.A1(\rbzero.wall_tracer.rayAddendX[-9] ),
    .A2(_09823_),
    .B1(_04005_),
    .X(_01647_));
 sky130_fd_sc_hd__xor2_1 _20877_ (.A(_02543_),
    .B(_02546_),
    .X(_04006_));
 sky130_fd_sc_hd__a22o_1 _20878_ (.A1(\rbzero.wall_tracer.rayAddendX[-8] ),
    .A2(_04000_),
    .B1(_03998_),
    .B2(_04006_),
    .X(_01648_));
 sky130_fd_sc_hd__and2b_1 _20879_ (.A_N(_02542_),
    .B(_02548_),
    .X(_04007_));
 sky130_fd_sc_hd__xnor2_1 _20880_ (.A(_02547_),
    .B(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__a22o_1 _20881_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_04000_),
    .B1(_03998_),
    .B2(_04008_),
    .X(_01649_));
 sky130_fd_sc_hd__nand2_1 _20882_ (.A(_02541_),
    .B(_02550_),
    .Y(_04009_));
 sky130_fd_sc_hd__xnor2_1 _20883_ (.A(_02549_),
    .B(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__a22o_1 _20884_ (.A1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .A2(_04000_),
    .B1(_02611_),
    .B2(_04010_),
    .X(_01650_));
 sky130_fd_sc_hd__xor2_1 _20885_ (.A(_05172_),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_04011_));
 sky130_fd_sc_hd__a22o_1 _20886_ (.A1(\rbzero.wall_tracer.rayAddendY[-9] ),
    .A2(_04000_),
    .B1(_02611_),
    .B2(_04011_),
    .X(_01651_));
 sky130_fd_sc_hd__a22o_1 _20887_ (.A1(_05172_),
    .A2(\rbzero.wall_tracer.rayAddendY[-9] ),
    .B1(_02778_),
    .B2(_02779_),
    .X(_04012_));
 sky130_fd_sc_hd__a32o_1 _20888_ (.A1(_09826_),
    .A2(_02780_),
    .A3(_04012_),
    .B1(_04000_),
    .B2(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_01652_));
 sky130_fd_sc_hd__and2b_1 _20889_ (.A_N(_02777_),
    .B(_02782_),
    .X(_04013_));
 sky130_fd_sc_hd__xnor2_1 _20890_ (.A(_02781_),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__a22o_1 _20891_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_04000_),
    .B1(_02611_),
    .B2(_04014_),
    .X(_01653_));
 sky130_fd_sc_hd__nand2_1 _20892_ (.A(_02776_),
    .B(_02784_),
    .Y(_04015_));
 sky130_fd_sc_hd__xnor2_1 _20893_ (.A(_02783_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__a22o_1 _20894_ (.A1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .A2(_04000_),
    .B1(_02611_),
    .B2(_04016_),
    .X(_01654_));
 sky130_fd_sc_hd__nor2_1 _20895_ (.A(\gpout1.clk_div[0] ),
    .B(net64),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_1 _20896_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .Y(_04017_));
 sky130_fd_sc_hd__or2_1 _20897_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .X(_04018_));
 sky130_fd_sc_hd__and3_1 _20898_ (.A(_09810_),
    .B(_04017_),
    .C(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__clkbuf_1 _20899_ (.A(_04019_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_1 _20900_ (.A(\gpout2.clk_div[0] ),
    .B(net64),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _20901_ (.A(\gpout2.clk_div[1] ),
    .B(\gpout2.clk_div[0] ),
    .Y(_04020_));
 sky130_fd_sc_hd__or2_1 _20902_ (.A(\gpout2.clk_div[1] ),
    .B(\gpout2.clk_div[0] ),
    .X(_04021_));
 sky130_fd_sc_hd__and3_1 _20903_ (.A(_09810_),
    .B(_04020_),
    .C(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_1 _20904_ (.A(_04022_),
    .X(_01658_));
 sky130_fd_sc_hd__nor2_1 _20905_ (.A(\gpout3.clk_div[0] ),
    .B(net64),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _20906_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .Y(_04023_));
 sky130_fd_sc_hd__or2_1 _20907_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .X(_04024_));
 sky130_fd_sc_hd__and3_1 _20908_ (.A(_09810_),
    .B(_04023_),
    .C(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__clkbuf_1 _20909_ (.A(_04025_),
    .X(_01660_));
 sky130_fd_sc_hd__nor2_1 _20910_ (.A(\gpout4.clk_div[0] ),
    .B(net64),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _20911_ (.A(\gpout4.clk_div[0] ),
    .B(\gpout4.clk_div[1] ),
    .Y(_04026_));
 sky130_fd_sc_hd__or2_1 _20912_ (.A(\gpout4.clk_div[0] ),
    .B(\gpout4.clk_div[1] ),
    .X(_04027_));
 sky130_fd_sc_hd__and3_1 _20913_ (.A(_03150_),
    .B(_04026_),
    .C(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_1 _20914_ (.A(_04028_),
    .X(_01662_));
 sky130_fd_sc_hd__dfxtp_1 _20915_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00000_),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20916_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00001_),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20917_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00386_),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20918_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00387_),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20919_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00388_),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20920_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00389_),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20921_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00390_),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20922_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00391_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_2 _20923_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00392_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20924_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00393_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20925_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00394_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20926_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00395_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20927_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00396_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20928_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00397_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20929_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00398_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00399_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20931_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00400_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20932_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00401_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20933_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00402_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00403_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20935_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00404_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20936_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00405_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20937_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20938_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20939_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20940_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20941_ (.CLK(clknet_4_15_0_i_clk),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20942_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20943_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_4 _20944_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00413_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20945_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00414_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _20946_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00415_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20947_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00416_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20948_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00417_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20949_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00418_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _20950_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00419_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20951_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00420_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_4 _20952_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00421_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _20953_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00422_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20954_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00423_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_4 _20955_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00424_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20956_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00425_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20957_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00426_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20958_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00427_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_4 _20959_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00428_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20960_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00429_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20961_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00430_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_4 _20962_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00431_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20963_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00432_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_4 _20964_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00433_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_4 _20965_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00434_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20966_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_2 _20967_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20970_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20973_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20976_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20977_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20979_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20984_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20985_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00457_),
    .Q(\reg_rgb[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00458_),
    .Q(\reg_rgb[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00459_),
    .Q(\reg_rgb[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00460_),
    .Q(\reg_rgb[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20992_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00461_),
    .Q(\reg_rgb[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20993_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00462_),
    .Q(\reg_rgb[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20994_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00463_),
    .Q(\rbzero.wall_hot[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20995_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00464_),
    .Q(\rbzero.wall_hot[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20996_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00465_),
    .Q(\rbzero.side_hot ));
 sky130_fd_sc_hd__dfxtp_2 _20997_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00466_),
    .Q(\rbzero.texu_hot[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20998_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00467_),
    .Q(\rbzero.texu_hot[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20999_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00468_),
    .Q(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21000_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00469_),
    .Q(\rbzero.texu_hot[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21001_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00470_),
    .Q(\rbzero.texu_hot[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21002_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00471_),
    .Q(\rbzero.texu_hot[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21003_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00472_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21004_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00473_),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_4 _21005_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00474_),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21006_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00475_),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21007_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00476_),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21008_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00477_),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21009_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00478_),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21010_ (.CLK(clknet_leaf_107_i_clk),
    .D(_00479_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_4 _21011_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00480_),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21012_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00481_),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_4 _21013_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00482_),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _21014_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00483_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21015_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00484_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21016_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00485_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21017_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00486_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21018_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00487_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00488_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21020_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00489_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21021_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00490_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21022_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00491_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21023_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00492_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21024_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00493_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21025_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00494_),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21026_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00495_),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21027_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00496_),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21028_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00497_),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21029_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00498_),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00499_),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21031_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00500_),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21032_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00501_),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21033_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00502_),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21034_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00503_),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00504_),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00505_),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21037_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00506_),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21038_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00507_),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21039_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00508_),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21040_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00509_),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21041_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00510_),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21042_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00511_),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21043_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00512_),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21044_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00513_),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21045_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00514_),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21046_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00515_),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21047_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00516_),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21048_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00517_),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21049_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00518_),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21050_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00519_),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21051_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00520_),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21052_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00521_),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21053_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00522_),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21054_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00523_),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21055_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00524_),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21056_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00525_),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21057_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00526_),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21058_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00527_),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21059_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00528_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_2 _21060_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00529_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21061_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00530_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21062_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00531_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00532_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00533_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00534_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00535_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00536_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21068_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00537_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00538_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00539_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21071_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00540_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21073_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21074_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21080_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21081_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21088_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21091_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21092_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21093_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21097_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21098_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21099_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21100_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21101_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21102_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21103_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00572_),
    .Q(\rbzero.spi_registers.new_texadd[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21104_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00573_),
    .Q(\rbzero.spi_registers.new_texadd[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21105_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00574_),
    .Q(\rbzero.spi_registers.new_texadd[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21106_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00575_),
    .Q(\rbzero.spi_registers.new_texadd[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21107_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00576_),
    .Q(\rbzero.spi_registers.new_texadd[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21108_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00577_),
    .Q(\rbzero.spi_registers.new_texadd[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21109_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00578_),
    .Q(\rbzero.spi_registers.new_texadd[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21110_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00579_),
    .Q(\rbzero.spi_registers.new_texadd[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21111_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00580_),
    .Q(\rbzero.spi_registers.new_texadd[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21112_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00581_),
    .Q(\rbzero.spi_registers.new_texadd[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21113_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00582_),
    .Q(\rbzero.spi_registers.new_texadd[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21114_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00583_),
    .Q(\rbzero.spi_registers.new_texadd[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21115_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00584_),
    .Q(\rbzero.spi_registers.new_texadd[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21116_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00585_),
    .Q(\rbzero.spi_registers.new_texadd[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21117_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00586_),
    .Q(\rbzero.spi_registers.new_texadd[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21118_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00587_),
    .Q(\rbzero.spi_registers.new_texadd[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21119_ (.CLK(clknet_leaf_134_i_clk),
    .D(_00588_),
    .Q(\rbzero.spi_registers.new_texadd[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21120_ (.CLK(clknet_leaf_134_i_clk),
    .D(_00589_),
    .Q(\rbzero.spi_registers.new_texadd[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00590_),
    .Q(\rbzero.spi_registers.new_texadd[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21122_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00591_),
    .Q(\rbzero.spi_registers.new_texadd[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00592_),
    .Q(\rbzero.spi_registers.new_texadd[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00593_),
    .Q(\rbzero.spi_registers.new_texadd[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21125_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00594_),
    .Q(\rbzero.spi_registers.new_texadd[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00595_),
    .Q(\rbzero.spi_registers.new_texadd[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21127_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00596_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21128_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00597_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21129_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00598_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21130_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00599_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21131_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00600_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00601_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21133_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00602_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21134_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00603_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21135_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00604_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21136_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00605_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00606_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21138_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00607_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21139_ (.CLK(clknet_4_11_0_i_clk),
    .D(_00608_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21140_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00609_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21141_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00610_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21142_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00611_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21143_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00612_),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_2 _21144_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00613_),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_1 _21145_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00614_),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_4 _21146_ (.CLK(clknet_4_6_0_i_clk),
    .D(_00615_),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_4 _21147_ (.CLK(clknet_leaf_110_i_clk),
    .D(_00616_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21148_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00617_),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21149_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00618_),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_1 _21150_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00619_),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_1 _21151_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00620_),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_1 _21152_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00621_),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_4 _21153_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00622_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21154_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00623_),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21155_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00624_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21156_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00625_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21157_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00626_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21158_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00627_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21159_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00628_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00629_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00630_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21162_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00631_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21163_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00632_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21164_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00633_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00634_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21166_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00635_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00636_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00637_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00638_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00639_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21171_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00640_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00641_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21173_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00642_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00643_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21175_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00644_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21176_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00645_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21177_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00646_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00647_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00648_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00649_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(clknet_leaf_128_i_clk),
    .D(_00650_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21182_ (.CLK(clknet_leaf_128_i_clk),
    .D(_00651_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(clknet_leaf_128_i_clk),
    .D(_00652_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21184_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00653_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(clknet_leaf_128_i_clk),
    .D(_00654_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(clknet_leaf_123_i_clk),
    .D(_00655_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00656_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00657_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21189_ (.CLK(clknet_leaf_125_i_clk),
    .D(_00658_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(clknet_leaf_126_i_clk),
    .D(_00659_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(clknet_leaf_127_i_clk),
    .D(_00660_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(clknet_leaf_127_i_clk),
    .D(_00661_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(clknet_leaf_127_i_clk),
    .D(_00662_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(clknet_leaf_126_i_clk),
    .D(_00663_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21195_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00664_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21196_ (.CLK(clknet_leaf_127_i_clk),
    .D(_00665_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00666_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21198_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00667_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00668_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00669_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00670_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00671_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00672_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00673_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21205_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00674_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21206_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00675_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00676_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(clknet_leaf_124_i_clk),
    .D(_00677_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21209_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00678_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21210_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00679_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00680_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21212_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00681_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00682_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21214_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00683_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21215_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00684_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21216_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00685_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00686_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00687_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00688_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21220_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00689_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00690_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00691_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00692_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00693_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21225_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00694_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21226_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00695_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21227_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00696_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00697_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00698_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00699_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00700_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00701_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00702_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00703_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00704_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00705_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00706_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00707_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00708_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00709_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00710_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00711_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00712_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00713_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21245_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00714_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00715_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21247_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00716_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21248_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00717_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00718_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00719_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00720_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00721_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00722_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00723_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00724_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00725_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00726_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21258_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00727_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21259_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00728_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21260_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00729_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21261_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00730_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21262_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00731_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21263_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00732_),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _21264_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00733_),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21265_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00734_),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _21266_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00735_),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _21267_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00736_),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(clknet_leaf_133_i_clk),
    .D(_00737_),
    .Q(\rbzero.spi_registers.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _21269_ (.CLK(clknet_leaf_134_i_clk),
    .D(_00738_),
    .Q(\rbzero.spi_registers.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(clknet_leaf_134_i_clk),
    .D(_00739_),
    .Q(\rbzero.spi_registers.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(clknet_leaf_135_i_clk),
    .D(_00740_),
    .Q(\rbzero.spi_registers.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(clknet_leaf_135_i_clk),
    .D(_00741_),
    .Q(\rbzero.spi_registers.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00742_),
    .Q(\rbzero.spi_registers.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00743_),
    .Q(\rbzero.spi_registers.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21275_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00744_),
    .Q(\rbzero.spi_registers.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_2 _21276_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00745_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21277_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00746_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21278_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00747_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00748_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21280_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00749_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00750_),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00751_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00752_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(clknet_leaf_130_i_clk),
    .D(_00753_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00754_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00755_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00756_),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00757_),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00758_),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00759_),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00760_),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00761_),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21293_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00762_),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21294_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00763_),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00764_),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00765_),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21297_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00766_),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00767_),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00768_),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00769_),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21301_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00770_),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00771_),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00772_),
    .Q(\rbzero.map_overlay.i_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00773_),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00774_),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00775_),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00776_),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00777_),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21309_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00778_),
    .Q(\rbzero.map_overlay.i_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21310_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00779_),
    .Q(\rbzero.mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00780_),
    .Q(\rbzero.mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00781_),
    .Q(\rbzero.mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00782_),
    .Q(\rbzero.mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00783_),
    .Q(\rbzero.spi_registers.texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00784_),
    .Q(\rbzero.spi_registers.texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00785_),
    .Q(\rbzero.spi_registers.texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00786_),
    .Q(\rbzero.spi_registers.texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00787_),
    .Q(\rbzero.spi_registers.texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00788_),
    .Q(\rbzero.spi_registers.texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00789_),
    .Q(\rbzero.spi_registers.texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00790_),
    .Q(\rbzero.spi_registers.texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00791_),
    .Q(\rbzero.spi_registers.texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00792_),
    .Q(\rbzero.spi_registers.texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00793_),
    .Q(\rbzero.spi_registers.texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00794_),
    .Q(\rbzero.spi_registers.texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00795_),
    .Q(\rbzero.spi_registers.texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00796_),
    .Q(\rbzero.spi_registers.texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00797_),
    .Q(\rbzero.spi_registers.texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00798_),
    .Q(\rbzero.spi_registers.texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00799_),
    .Q(\rbzero.spi_registers.texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00800_),
    .Q(\rbzero.spi_registers.texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00801_),
    .Q(\rbzero.spi_registers.texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00802_),
    .Q(\rbzero.spi_registers.texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00803_),
    .Q(\rbzero.spi_registers.texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00804_),
    .Q(\rbzero.spi_registers.texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00805_),
    .Q(\rbzero.spi_registers.texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00806_),
    .Q(\rbzero.spi_registers.texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00807_),
    .Q(\rbzero.spi_registers.texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00808_),
    .Q(\rbzero.spi_registers.texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00809_),
    .Q(\rbzero.spi_registers.texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00810_),
    .Q(\rbzero.spi_registers.texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00811_),
    .Q(\rbzero.spi_registers.texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00812_),
    .Q(\rbzero.spi_registers.texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00813_),
    .Q(\rbzero.spi_registers.texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00814_),
    .Q(\rbzero.spi_registers.texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00815_),
    .Q(\rbzero.spi_registers.texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00816_),
    .Q(\rbzero.spi_registers.texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00817_),
    .Q(\rbzero.spi_registers.texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00818_),
    .Q(\rbzero.spi_registers.texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00819_),
    .Q(\rbzero.spi_registers.texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00820_),
    .Q(\rbzero.spi_registers.texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00821_),
    .Q(\rbzero.spi_registers.texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00822_),
    .Q(\rbzero.spi_registers.texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00823_),
    .Q(\rbzero.spi_registers.texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(clknet_leaf_135_i_clk),
    .D(_00824_),
    .Q(\rbzero.spi_registers.texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(clknet_leaf_135_i_clk),
    .D(_00825_),
    .Q(\rbzero.spi_registers.texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(clknet_leaf_135_i_clk),
    .D(_00826_),
    .Q(\rbzero.spi_registers.texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00827_),
    .Q(\rbzero.spi_registers.texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00828_),
    .Q(\rbzero.spi_registers.texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00829_),
    .Q(\rbzero.spi_registers.texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00830_),
    .Q(\rbzero.spi_registers.texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00831_),
    .Q(\rbzero.spi_registers.texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00832_),
    .Q(\rbzero.spi_registers.texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00833_),
    .Q(\rbzero.spi_registers.texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00834_),
    .Q(\rbzero.spi_registers.texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00835_),
    .Q(\rbzero.spi_registers.texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00836_),
    .Q(\rbzero.spi_registers.texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00837_),
    .Q(\rbzero.spi_registers.texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00838_),
    .Q(\rbzero.spi_registers.texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00839_),
    .Q(\rbzero.spi_registers.texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00840_),
    .Q(\rbzero.spi_registers.texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00841_),
    .Q(\rbzero.spi_registers.texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00842_),
    .Q(\rbzero.spi_registers.texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00843_),
    .Q(\rbzero.spi_registers.texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00844_),
    .Q(\rbzero.spi_registers.texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00845_),
    .Q(\rbzero.spi_registers.texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00846_),
    .Q(\rbzero.spi_registers.texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00847_),
    .Q(\rbzero.spi_registers.texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00848_),
    .Q(\rbzero.spi_registers.texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00849_),
    .Q(\rbzero.spi_registers.texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00850_),
    .Q(\rbzero.spi_registers.texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00851_),
    .Q(\rbzero.spi_registers.texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00852_),
    .Q(\rbzero.spi_registers.texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00853_),
    .Q(\rbzero.spi_registers.texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00854_),
    .Q(\rbzero.spi_registers.texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00855_),
    .Q(\rbzero.spi_registers.texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00856_),
    .Q(\rbzero.spi_registers.texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00857_),
    .Q(\rbzero.spi_registers.texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00858_),
    .Q(\rbzero.spi_registers.texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00859_),
    .Q(\rbzero.spi_registers.texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00860_),
    .Q(\rbzero.spi_registers.texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00861_),
    .Q(\rbzero.spi_registers.texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00862_),
    .Q(\rbzero.spi_registers.texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00863_),
    .Q(\rbzero.spi_registers.texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00864_),
    .Q(\rbzero.spi_registers.texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00865_),
    .Q(\rbzero.spi_registers.texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00866_),
    .Q(\rbzero.spi_registers.texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00867_),
    .Q(\rbzero.spi_registers.texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00868_),
    .Q(\rbzero.spi_registers.texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00869_),
    .Q(\rbzero.spi_registers.texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00870_),
    .Q(\rbzero.spi_registers.texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(clknet_leaf_134_i_clk),
    .D(_00871_),
    .Q(\rbzero.spi_registers.texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(clknet_leaf_134_i_clk),
    .D(_00872_),
    .Q(\rbzero.spi_registers.texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00873_),
    .Q(\rbzero.spi_registers.texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00874_),
    .Q(\rbzero.spi_registers.texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00875_),
    .Q(\rbzero.spi_registers.texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00876_),
    .Q(\rbzero.spi_registers.texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00877_),
    .Q(\rbzero.spi_registers.texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21409_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00878_),
    .Q(\rbzero.spi_registers.texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21410_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00879_),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21411_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00880_),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21412_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00881_),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21413_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00882_),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00883_),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00884_),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21416_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00885_),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00886_),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00887_),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21419_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00888_),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00889_),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00890_),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00891_),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00892_),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21424_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00893_),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21425_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00894_),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00895_),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00896_),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00897_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00898_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00899_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21431_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00900_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21432_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00901_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21433_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00902_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21434_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00903_),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00904_),
    .Q(\rbzero.spi_registers.new_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21436_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00905_),
    .Q(\rbzero.spi_registers.new_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21437_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00906_),
    .Q(\rbzero.spi_registers.new_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21438_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00907_),
    .Q(\rbzero.spi_registers.new_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00908_),
    .Q(\rbzero.spi_registers.new_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21440_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00909_),
    .Q(\rbzero.spi_registers.new_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21441_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00910_),
    .Q(\rbzero.spi_registers.got_new_sky ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00911_),
    .Q(\rbzero.spi_registers.new_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00912_),
    .Q(\rbzero.spi_registers.new_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00913_),
    .Q(\rbzero.spi_registers.new_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00914_),
    .Q(\rbzero.spi_registers.new_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00915_),
    .Q(\rbzero.spi_registers.new_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21447_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00916_),
    .Q(\rbzero.spi_registers.new_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00917_),
    .Q(\rbzero.spi_registers.got_new_floor ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00918_),
    .Q(\rbzero.spi_registers.new_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21450_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00919_),
    .Q(\rbzero.spi_registers.new_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00920_),
    .Q(\rbzero.spi_registers.new_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00921_),
    .Q(\rbzero.spi_registers.new_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00922_),
    .Q(\rbzero.spi_registers.new_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00923_),
    .Q(\rbzero.spi_registers.new_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00924_),
    .Q(\rbzero.spi_registers.got_new_leak ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00925_),
    .Q(\rbzero.spi_registers.new_other[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00926_),
    .Q(\rbzero.spi_registers.new_other[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00927_),
    .Q(\rbzero.spi_registers.new_other[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00928_),
    .Q(\rbzero.spi_registers.new_other[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21460_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00929_),
    .Q(\rbzero.spi_registers.new_other[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21461_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00930_),
    .Q(\rbzero.spi_registers.new_other[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21462_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00931_),
    .Q(\rbzero.spi_registers.new_other[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21463_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00932_),
    .Q(\rbzero.spi_registers.new_other[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00933_),
    .Q(\rbzero.spi_registers.new_other[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21465_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00934_),
    .Q(\rbzero.spi_registers.new_other[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00935_),
    .Q(\rbzero.spi_registers.got_new_other ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00936_),
    .Q(\rbzero.spi_registers.new_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21468_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00937_),
    .Q(\rbzero.spi_registers.new_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21469_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00938_),
    .Q(\rbzero.spi_registers.new_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21470_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00939_),
    .Q(\rbzero.spi_registers.new_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(clknet_leaf_38_i_clk),
    .D(_00940_),
    .Q(\rbzero.spi_registers.new_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21472_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00941_),
    .Q(\rbzero.spi_registers.new_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21473_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00942_),
    .Q(\rbzero.spi_registers.got_new_vshift ));
 sky130_fd_sc_hd__dfxtp_1 _21474_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00943_),
    .Q(\rbzero.spi_registers.new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00944_),
    .Q(\rbzero.spi_registers.got_new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21476_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00945_),
    .Q(\rbzero.spi_registers.new_mapd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00946_),
    .Q(\rbzero.spi_registers.new_mapd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00947_),
    .Q(\rbzero.spi_registers.new_mapd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00948_),
    .Q(\rbzero.spi_registers.new_mapd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00949_),
    .Q(\rbzero.spi_registers.new_mapd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00950_),
    .Q(\rbzero.spi_registers.new_mapd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00951_),
    .Q(\rbzero.spi_registers.new_mapd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21483_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00952_),
    .Q(\rbzero.spi_registers.new_mapd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00953_),
    .Q(\rbzero.spi_registers.new_mapd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00954_),
    .Q(\rbzero.spi_registers.new_mapd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21486_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00955_),
    .Q(\rbzero.spi_registers.new_mapd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00956_),
    .Q(\rbzero.spi_registers.new_mapd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21488_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00957_),
    .Q(\rbzero.spi_registers.new_mapd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21489_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00958_),
    .Q(\rbzero.spi_registers.new_mapd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21490_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00959_),
    .Q(\rbzero.spi_registers.new_mapd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21491_ (.CLK(clknet_leaf_131_i_clk),
    .D(_00960_),
    .Q(\rbzero.spi_registers.new_mapd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21492_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00961_),
    .Q(\rbzero.spi_registers.got_new_mapd ));
 sky130_fd_sc_hd__dfxtp_1 _21493_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00962_),
    .Q(\rbzero.spi_registers.got_new_texadd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00963_),
    .Q(\rbzero.spi_registers.got_new_texadd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21495_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00964_),
    .Q(\rbzero.spi_registers.got_new_texadd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21496_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00965_),
    .Q(\rbzero.spi_registers.got_new_texadd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21497_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00966_),
    .Q(\rbzero.spi_registers.new_texadd[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21498_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00967_),
    .Q(\rbzero.spi_registers.new_texadd[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21499_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00968_),
    .Q(\rbzero.spi_registers.new_texadd[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21500_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00969_),
    .Q(\rbzero.spi_registers.new_texadd[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21501_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00970_),
    .Q(\rbzero.spi_registers.new_texadd[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21502_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00971_),
    .Q(\rbzero.spi_registers.new_texadd[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21503_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00972_),
    .Q(\rbzero.spi_registers.new_texadd[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21504_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00973_),
    .Q(\rbzero.spi_registers.new_texadd[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00974_),
    .Q(\rbzero.spi_registers.new_texadd[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21506_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00975_),
    .Q(\rbzero.spi_registers.new_texadd[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00976_),
    .Q(\rbzero.spi_registers.new_texadd[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00977_),
    .Q(\rbzero.spi_registers.new_texadd[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00978_),
    .Q(\rbzero.spi_registers.new_texadd[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21510_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00979_),
    .Q(\rbzero.spi_registers.new_texadd[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21511_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00980_),
    .Q(\rbzero.spi_registers.new_texadd[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21512_ (.CLK(clknet_leaf_132_i_clk),
    .D(_00981_),
    .Q(\rbzero.spi_registers.new_texadd[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21513_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00982_),
    .Q(\rbzero.spi_registers.new_texadd[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21514_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00983_),
    .Q(\rbzero.spi_registers.new_texadd[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21515_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00984_),
    .Q(\rbzero.spi_registers.new_texadd[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21516_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00985_),
    .Q(\rbzero.spi_registers.new_texadd[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21517_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00986_),
    .Q(\rbzero.spi_registers.new_texadd[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21518_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00987_),
    .Q(\rbzero.spi_registers.new_texadd[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00988_),
    .Q(\rbzero.spi_registers.new_texadd[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00989_),
    .Q(\rbzero.spi_registers.new_texadd[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21521_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00990_),
    .Q(\rbzero.spi_registers.new_texadd[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21522_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00991_),
    .Q(\rbzero.spi_registers.new_texadd[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21523_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00992_),
    .Q(\rbzero.spi_registers.new_texadd[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21524_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00993_),
    .Q(\rbzero.spi_registers.new_texadd[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00994_),
    .Q(\rbzero.spi_registers.new_texadd[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00995_),
    .Q(\rbzero.spi_registers.new_texadd[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00996_),
    .Q(\rbzero.spi_registers.new_texadd[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21528_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00997_),
    .Q(\rbzero.spi_registers.new_texadd[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21529_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00998_),
    .Q(\rbzero.spi_registers.new_texadd[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00999_),
    .Q(\rbzero.spi_registers.new_texadd[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21531_ (.CLK(clknet_leaf_9_i_clk),
    .D(_01000_),
    .Q(\rbzero.spi_registers.new_texadd[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21532_ (.CLK(clknet_leaf_0_i_clk),
    .D(_01001_),
    .Q(\rbzero.spi_registers.new_texadd[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(clknet_leaf_0_i_clk),
    .D(_01002_),
    .Q(\rbzero.spi_registers.new_texadd[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21534_ (.CLK(clknet_leaf_9_i_clk),
    .D(_01003_),
    .Q(\rbzero.spi_registers.new_texadd[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21535_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01004_),
    .Q(\rbzero.spi_registers.new_texadd[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(clknet_leaf_3_i_clk),
    .D(_01005_),
    .Q(\rbzero.spi_registers.new_texadd[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21537_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01006_),
    .Q(\rbzero.spi_registers.new_texadd[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01007_),
    .Q(\rbzero.spi_registers.new_texadd[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21539_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01008_),
    .Q(\rbzero.spi_registers.new_texadd[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01009_),
    .Q(\rbzero.spi_registers.new_texadd[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21541_ (.CLK(clknet_leaf_10_i_clk),
    .D(_01010_),
    .Q(\rbzero.spi_registers.new_texadd[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21542_ (.CLK(clknet_leaf_11_i_clk),
    .D(_01011_),
    .Q(\rbzero.spi_registers.new_texadd[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21543_ (.CLK(clknet_leaf_11_i_clk),
    .D(_01012_),
    .Q(\rbzero.spi_registers.new_texadd[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(clknet_leaf_16_i_clk),
    .D(_01013_),
    .Q(\rbzero.spi_registers.new_texadd[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21545_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01014_),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _21546_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01015_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01016_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21548_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01017_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01018_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21550_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01019_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01020_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21552_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01021_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21553_ (.CLK(net153),
    .D(_01022_),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21554_ (.CLK(net154),
    .D(_01023_),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(net155),
    .D(_01024_),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21556_ (.CLK(net156),
    .D(_01025_),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21557_ (.CLK(net157),
    .D(_01026_),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21558_ (.CLK(net158),
    .D(_01027_),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21559_ (.CLK(net159),
    .D(_01028_),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(net160),
    .D(_01029_),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(net161),
    .D(_01030_),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(net162),
    .D(_01031_),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(net163),
    .D(_01032_),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(net164),
    .D(_01033_),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(net165),
    .D(_01034_),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21566_ (.CLK(net166),
    .D(_01035_),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(net167),
    .D(_01036_),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21568_ (.CLK(net168),
    .D(_01037_),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(net169),
    .D(_01038_),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(net170),
    .D(_01039_),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(net171),
    .D(_01040_),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21572_ (.CLK(net172),
    .D(_01041_),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(net173),
    .D(_01042_),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(net174),
    .D(_01043_),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(net175),
    .D(_01044_),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(net176),
    .D(_01045_),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21577_ (.CLK(net177),
    .D(_01046_),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21578_ (.CLK(net178),
    .D(_01047_),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21579_ (.CLK(net179),
    .D(_01048_),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(net180),
    .D(_01049_),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21581_ (.CLK(net181),
    .D(_01050_),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21582_ (.CLK(net182),
    .D(_01051_),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(net183),
    .D(_01052_),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21584_ (.CLK(net184),
    .D(_01053_),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21585_ (.CLK(net185),
    .D(_01054_),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21586_ (.CLK(net186),
    .D(_01055_),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21587_ (.CLK(net187),
    .D(_01056_),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21588_ (.CLK(net188),
    .D(_01057_),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21589_ (.CLK(net189),
    .D(_01058_),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21590_ (.CLK(net190),
    .D(_01059_),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21591_ (.CLK(net191),
    .D(_01060_),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(net192),
    .D(_01061_),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21593_ (.CLK(net193),
    .D(_01062_),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21594_ (.CLK(net194),
    .D(_01063_),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(net195),
    .D(_01064_),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21596_ (.CLK(net196),
    .D(_01065_),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21597_ (.CLK(net197),
    .D(_01066_),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(net198),
    .D(_01067_),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21599_ (.CLK(net199),
    .D(_01068_),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21600_ (.CLK(net200),
    .D(_01069_),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21601_ (.CLK(net201),
    .D(_01070_),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21602_ (.CLK(net202),
    .D(_01071_),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21603_ (.CLK(net203),
    .D(_01072_),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21604_ (.CLK(net204),
    .D(_01073_),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21605_ (.CLK(net205),
    .D(_01074_),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21606_ (.CLK(net206),
    .D(_01075_),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(net207),
    .D(_01076_),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(net208),
    .D(_01077_),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21609_ (.CLK(net209),
    .D(_01078_),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(net210),
    .D(_01079_),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(net211),
    .D(_01080_),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(net212),
    .D(_01081_),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(net213),
    .D(_01082_),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21614_ (.CLK(net214),
    .D(_01083_),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(net215),
    .D(_01084_),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(net216),
    .D(_01085_),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01086_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21618_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01087_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21619_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01088_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01089_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01090_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01091_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01092_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01093_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01094_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21626_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01095_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01096_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01097_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21629_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01098_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21630_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01099_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21631_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01100_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21632_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01101_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01102_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21634_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01103_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21635_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01104_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21636_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01105_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21637_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01106_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21638_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01107_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01108_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21640_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01109_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21641_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01110_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21642_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01111_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21643_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01112_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01113_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21645_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01114_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21646_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01115_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21647_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01116_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21648_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01117_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21649_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01118_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21650_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01119_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21651_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01120_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01121_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01122_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01123_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21655_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01124_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01125_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01126_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01127_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21659_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01128_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01129_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01130_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(clknet_leaf_104_i_clk),
    .D(_01131_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01132_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01133_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01134_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01135_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21667_ (.CLK(clknet_leaf_119_i_clk),
    .D(_01136_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(clknet_leaf_119_i_clk),
    .D(_01137_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21669_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01138_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21670_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01139_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21671_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01140_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21672_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01141_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21673_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01142_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21674_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01143_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21675_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01144_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01145_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21677_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01146_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01147_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01148_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01149_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01150_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21682_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01151_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01152_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01153_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21685_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01154_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21686_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01155_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21687_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01156_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01157_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21689_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01158_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21690_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01159_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21691_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01160_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01161_),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21693_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01162_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21694_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01163_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21695_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01164_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21696_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01165_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01166_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21698_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01167_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21699_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01168_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01169_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(clknet_leaf_103_i_clk),
    .D(_01170_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21702_ (.CLK(clknet_leaf_104_i_clk),
    .D(_01171_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21703_ (.CLK(clknet_leaf_103_i_clk),
    .D(_01172_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21704_ (.CLK(clknet_leaf_104_i_clk),
    .D(_01173_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _21705_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01174_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21706_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01175_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21707_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01176_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21708_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01177_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21709_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01178_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21710_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01179_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21711_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01180_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21712_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01181_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21713_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01182_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21714_ (.CLK(clknet_leaf_103_i_clk),
    .D(_01183_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21715_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01184_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21716_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01185_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21717_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01186_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21718_ (.CLK(clknet_leaf_102_i_clk),
    .D(_01187_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21719_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01188_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21720_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01189_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21721_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01190_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21722_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01191_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21723_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01192_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21724_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01193_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21725_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01194_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21726_ (.CLK(clknet_leaf_119_i_clk),
    .D(_01195_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21727_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01196_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01197_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01198_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01199_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21731_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01200_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21732_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01201_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21733_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01202_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21734_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01203_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21735_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01204_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21736_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01205_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21737_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01206_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21738_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01207_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21739_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01208_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21740_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01209_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21741_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01210_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21742_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01211_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21743_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01212_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21744_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01213_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21745_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01214_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21746_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01215_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21747_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01216_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21748_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01217_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21749_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01218_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_4 _21750_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01219_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21751_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01220_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21752_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01221_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21753_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01222_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21754_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01223_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_4 _21755_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01224_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21756_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01225_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21757_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01226_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21758_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01227_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21759_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01228_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01229_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01230_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21762_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01231_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_4 _21763_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01232_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_4 _21764_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01233_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21765_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01234_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_4 _21766_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01235_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_4 _21767_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01236_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21768_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01237_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _21769_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01238_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21770_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01239_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21771_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01240_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21772_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01241_),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21773_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01242_),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01243_),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_1 _21775_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01244_),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21776_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01245_),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21777_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01246_),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21778_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01247_),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21779_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01248_),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01249_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21781_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01250_),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21782_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01251_),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21783_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01252_),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21784_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01253_),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(clknet_leaf_19_i_clk),
    .D(_01254_),
    .Q(\rbzero.spi_registers.new_texadd[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21786_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01255_),
    .Q(\rbzero.spi_registers.new_texadd[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21787_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01256_),
    .Q(\rbzero.spi_registers.new_texadd[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21788_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01257_),
    .Q(\rbzero.spi_registers.new_texadd[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21789_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01258_),
    .Q(\rbzero.spi_registers.new_texadd[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21790_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01259_),
    .Q(\rbzero.spi_registers.new_texadd[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21791_ (.CLK(clknet_leaf_19_i_clk),
    .D(_01260_),
    .Q(\rbzero.spi_registers.new_texadd[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21792_ (.CLK(clknet_leaf_20_i_clk),
    .D(_01261_),
    .Q(\rbzero.spi_registers.new_texadd[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21793_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01262_),
    .Q(\rbzero.spi_registers.new_texadd[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21794_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01263_),
    .Q(\rbzero.spi_registers.new_texadd[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21795_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01264_),
    .Q(\rbzero.spi_registers.new_texadd[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21796_ (.CLK(clknet_leaf_2_i_clk),
    .D(_01265_),
    .Q(\rbzero.spi_registers.new_texadd[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01266_),
    .Q(\rbzero.spi_registers.new_texadd[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21798_ (.CLK(clknet_leaf_5_i_clk),
    .D(_01267_),
    .Q(\rbzero.spi_registers.new_texadd[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21799_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01268_),
    .Q(\rbzero.spi_registers.new_texadd[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21800_ (.CLK(clknet_leaf_2_i_clk),
    .D(_01269_),
    .Q(\rbzero.spi_registers.new_texadd[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01270_),
    .Q(\rbzero.spi_registers.new_texadd[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21802_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01271_),
    .Q(\rbzero.spi_registers.new_texadd[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21803_ (.CLK(clknet_leaf_0_i_clk),
    .D(_01272_),
    .Q(\rbzero.spi_registers.new_texadd[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21804_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01273_),
    .Q(\rbzero.spi_registers.new_texadd[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(clknet_leaf_11_i_clk),
    .D(_01274_),
    .Q(\rbzero.spi_registers.new_texadd[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(clknet_leaf_11_i_clk),
    .D(_01275_),
    .Q(\rbzero.spi_registers.new_texadd[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21807_ (.CLK(clknet_leaf_11_i_clk),
    .D(_01276_),
    .Q(\rbzero.spi_registers.new_texadd[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(clknet_leaf_12_i_clk),
    .D(_01277_),
    .Q(\rbzero.spi_registers.new_texadd[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(net217),
    .D(_01278_),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(net218),
    .D(_01279_),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(net219),
    .D(_01280_),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(net220),
    .D(_01281_),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(net221),
    .D(_01282_),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(net222),
    .D(_01283_),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21815_ (.CLK(net223),
    .D(_01284_),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21816_ (.CLK(net224),
    .D(_01285_),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21817_ (.CLK(net225),
    .D(_01286_),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(net226),
    .D(_01287_),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21819_ (.CLK(net227),
    .D(_01288_),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21820_ (.CLK(net228),
    .D(_01289_),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(net229),
    .D(_01290_),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21822_ (.CLK(net230),
    .D(_01291_),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21823_ (.CLK(net231),
    .D(_01292_),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21824_ (.CLK(net232),
    .D(_01293_),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21825_ (.CLK(net233),
    .D(_01294_),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21826_ (.CLK(net234),
    .D(_01295_),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21827_ (.CLK(net235),
    .D(_01296_),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21828_ (.CLK(net236),
    .D(_01297_),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21829_ (.CLK(net237),
    .D(_01298_),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21830_ (.CLK(net238),
    .D(_01299_),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21831_ (.CLK(net239),
    .D(_01300_),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21832_ (.CLK(net240),
    .D(_01301_),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21833_ (.CLK(net241),
    .D(_01302_),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(net242),
    .D(_01303_),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(net243),
    .D(_01304_),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(net244),
    .D(_01305_),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(net245),
    .D(_01306_),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(net246),
    .D(_01307_),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21839_ (.CLK(net247),
    .D(_01308_),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(net248),
    .D(_01309_),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21841_ (.CLK(net249),
    .D(_01310_),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21842_ (.CLK(net250),
    .D(_01311_),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21843_ (.CLK(net251),
    .D(_01312_),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21844_ (.CLK(net252),
    .D(_01313_),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(net253),
    .D(_01314_),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21846_ (.CLK(net254),
    .D(_01315_),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21847_ (.CLK(net255),
    .D(_01316_),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21848_ (.CLK(net256),
    .D(_01317_),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(net257),
    .D(_01318_),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(net258),
    .D(_01319_),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(net259),
    .D(_01320_),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(net260),
    .D(_01321_),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21853_ (.CLK(net261),
    .D(_01322_),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(net262),
    .D(_01323_),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(net263),
    .D(_01324_),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(net264),
    .D(_01325_),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(net265),
    .D(_01326_),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(net266),
    .D(_01327_),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(net267),
    .D(_01328_),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(net268),
    .D(_01329_),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(net269),
    .D(_01330_),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(net270),
    .D(_01331_),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21863_ (.CLK(net271),
    .D(_01332_),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(net272),
    .D(_01333_),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(net273),
    .D(_01334_),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(net274),
    .D(_01335_),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(net275),
    .D(_01336_),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(net276),
    .D(_01337_),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(net277),
    .D(_01338_),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(net278),
    .D(_01339_),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(net279),
    .D(_01340_),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(net280),
    .D(_01341_),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21873_ (.CLK(net281),
    .D(_01342_),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21874_ (.CLK(net282),
    .D(_01343_),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(net283),
    .D(_01344_),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(net284),
    .D(_01345_),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(net285),
    .D(_01346_),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21878_ (.CLK(net286),
    .D(_01347_),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21879_ (.CLK(net287),
    .D(_01348_),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21880_ (.CLK(net288),
    .D(_01349_),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(net289),
    .D(_01350_),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21882_ (.CLK(net290),
    .D(_01351_),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(net291),
    .D(_01352_),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(net292),
    .D(_01353_),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(net293),
    .D(_01354_),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(net294),
    .D(_01355_),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(net295),
    .D(_01356_),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(net296),
    .D(_01357_),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(net297),
    .D(_01358_),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(net298),
    .D(_01359_),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(net299),
    .D(_01360_),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(net300),
    .D(_01361_),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(net301),
    .D(_01362_),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(net302),
    .D(_01363_),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21895_ (.CLK(net303),
    .D(_01364_),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(net304),
    .D(_01365_),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(net305),
    .D(_01366_),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21898_ (.CLK(net306),
    .D(_01367_),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(net307),
    .D(_01368_),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(net308),
    .D(_01369_),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(net309),
    .D(_01370_),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(net310),
    .D(_01371_),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(net311),
    .D(_01372_),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(net312),
    .D(_01373_),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(net313),
    .D(_01374_),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(net314),
    .D(_01375_),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(net315),
    .D(_01376_),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(net316),
    .D(_01377_),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21909_ (.CLK(net317),
    .D(_01378_),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(net318),
    .D(_01379_),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21911_ (.CLK(net319),
    .D(_01380_),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(net320),
    .D(_01381_),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(net321),
    .D(_01382_),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(net322),
    .D(_01383_),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21915_ (.CLK(net323),
    .D(_01384_),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(net324),
    .D(_01385_),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(net325),
    .D(_01386_),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(net326),
    .D(_01387_),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(net327),
    .D(_01388_),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(net328),
    .D(_01389_),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(net329),
    .D(_01390_),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(net330),
    .D(_01391_),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(net331),
    .D(_01392_),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(net332),
    .D(_01393_),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(net333),
    .D(_01394_),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21926_ (.CLK(net334),
    .D(_01395_),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(net335),
    .D(_01396_),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(net336),
    .D(_01397_),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(net337),
    .D(_01398_),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21930_ (.CLK(net338),
    .D(_01399_),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21931_ (.CLK(net339),
    .D(_01400_),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(net340),
    .D(_01401_),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(net341),
    .D(_01402_),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(net342),
    .D(_01403_),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(net343),
    .D(_01404_),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(net344),
    .D(_01405_),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(net345),
    .D(_01406_),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(net346),
    .D(_01407_),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(net347),
    .D(_01408_),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(net348),
    .D(_01409_),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(net349),
    .D(_01410_),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(net350),
    .D(_01411_),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(net351),
    .D(_01412_),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21944_ (.CLK(net352),
    .D(_01413_),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(net353),
    .D(_01414_),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21946_ (.CLK(net354),
    .D(_01415_),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21947_ (.CLK(net355),
    .D(_01416_),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21948_ (.CLK(net356),
    .D(_01417_),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21949_ (.CLK(net357),
    .D(_01418_),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21950_ (.CLK(net358),
    .D(_01419_),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(net359),
    .D(_01420_),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(net360),
    .D(_01421_),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(net361),
    .D(_01422_),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(net362),
    .D(_01423_),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(net363),
    .D(_01424_),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(net364),
    .D(_01425_),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(net365),
    .D(_01426_),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21958_ (.CLK(net366),
    .D(_01427_),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(net367),
    .D(_01428_),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21960_ (.CLK(net368),
    .D(_01429_),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(net369),
    .D(_01430_),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(net370),
    .D(_01431_),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21963_ (.CLK(net371),
    .D(_01432_),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(net372),
    .D(_01433_),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(net373),
    .D(_01434_),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(net374),
    .D(_01435_),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21967_ (.CLK(net375),
    .D(_01436_),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(net376),
    .D(_01437_),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(net377),
    .D(_01438_),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(net378),
    .D(_01439_),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21971_ (.CLK(net379),
    .D(_01440_),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(net380),
    .D(_01441_),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(net381),
    .D(_01442_),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(net382),
    .D(_01443_),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(net383),
    .D(_01444_),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(net384),
    .D(_01445_),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(net385),
    .D(_01446_),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(net386),
    .D(_01447_),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(net387),
    .D(_01448_),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(net388),
    .D(_01449_),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(net389),
    .D(_01450_),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(net390),
    .D(_01451_),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(net391),
    .D(_01452_),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(net392),
    .D(_01453_),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(net393),
    .D(_01454_),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(net394),
    .D(_01455_),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(net395),
    .D(_01456_),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(net396),
    .D(_01457_),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(net397),
    .D(_01458_),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(net398),
    .D(_01459_),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21991_ (.CLK(net399),
    .D(_01460_),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21992_ (.CLK(net400),
    .D(_01461_),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(net401),
    .D(_01462_),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(net402),
    .D(_01463_),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(net403),
    .D(_01464_),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(net404),
    .D(_01465_),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(net405),
    .D(_01466_),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21998_ (.CLK(net406),
    .D(_01467_),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(net407),
    .D(_01468_),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(net408),
    .D(_01469_),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(net409),
    .D(_01470_),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(net410),
    .D(_01471_),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(net411),
    .D(_01472_),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(net412),
    .D(_01473_),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(net413),
    .D(_01474_),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(net414),
    .D(_01475_),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(net415),
    .D(_01476_),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(net416),
    .D(_01477_),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(net417),
    .D(_01478_),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(net418),
    .D(_01479_),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(net419),
    .D(_01480_),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22012_ (.CLK(net420),
    .D(_01481_),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22013_ (.CLK(net421),
    .D(_01482_),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(net422),
    .D(_01483_),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(net423),
    .D(_01484_),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(net424),
    .D(_01485_),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(net425),
    .D(_01486_),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(net426),
    .D(_01487_),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(net427),
    .D(_01488_),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(net428),
    .D(_01489_),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(net429),
    .D(_01490_),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22022_ (.CLK(net430),
    .D(_01491_),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(net431),
    .D(_01492_),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(net432),
    .D(_01493_),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(net433),
    .D(_01494_),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(net434),
    .D(_01495_),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(net435),
    .D(_01496_),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(net436),
    .D(_01497_),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(net437),
    .D(_01498_),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(net438),
    .D(_01499_),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(net439),
    .D(_01500_),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(net440),
    .D(_01501_),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22033_ (.CLK(net441),
    .D(_01502_),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(net442),
    .D(_01503_),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(net443),
    .D(_01504_),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22036_ (.CLK(net444),
    .D(_01505_),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(net445),
    .D(_01506_),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(net446),
    .D(_01507_),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(net447),
    .D(_01508_),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(net448),
    .D(_01509_),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(net449),
    .D(_01510_),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(net450),
    .D(_01511_),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(net451),
    .D(_01512_),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(net452),
    .D(_01513_),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(net453),
    .D(_01514_),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22046_ (.CLK(net454),
    .D(_01515_),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22047_ (.CLK(net455),
    .D(_01516_),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22048_ (.CLK(net456),
    .D(_01517_),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22049_ (.CLK(net457),
    .D(_01518_),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22050_ (.CLK(net458),
    .D(_01519_),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22051_ (.CLK(net459),
    .D(_01520_),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22052_ (.CLK(net460),
    .D(_01521_),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22053_ (.CLK(net461),
    .D(_01522_),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22054_ (.CLK(net462),
    .D(_01523_),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22055_ (.CLK(net463),
    .D(_01524_),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22056_ (.CLK(net464),
    .D(_01525_),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22057_ (.CLK(net465),
    .D(_01526_),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22058_ (.CLK(net466),
    .D(_01527_),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22059_ (.CLK(net467),
    .D(_01528_),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22060_ (.CLK(net468),
    .D(_01529_),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22061_ (.CLK(net469),
    .D(_01530_),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22062_ (.CLK(net470),
    .D(_01531_),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22063_ (.CLK(net471),
    .D(_01532_),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22064_ (.CLK(net472),
    .D(_01533_),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22065_ (.CLK(net473),
    .D(_01534_),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22066_ (.CLK(net474),
    .D(_01535_),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22067_ (.CLK(net475),
    .D(_01536_),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22068_ (.CLK(net476),
    .D(_01537_),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22069_ (.CLK(net477),
    .D(_01538_),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22070_ (.CLK(net478),
    .D(_01539_),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22071_ (.CLK(net479),
    .D(_01540_),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22072_ (.CLK(net480),
    .D(_01541_),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22073_ (.CLK(net481),
    .D(_01542_),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22074_ (.CLK(net482),
    .D(_01543_),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22075_ (.CLK(net483),
    .D(_01544_),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22076_ (.CLK(net484),
    .D(_01545_),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22077_ (.CLK(net485),
    .D(_01546_),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22078_ (.CLK(net486),
    .D(_01547_),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22079_ (.CLK(net487),
    .D(_01548_),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22080_ (.CLK(net488),
    .D(_01549_),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22081_ (.CLK(net489),
    .D(_01550_),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22082_ (.CLK(net490),
    .D(_01551_),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22083_ (.CLK(net491),
    .D(_01552_),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22084_ (.CLK(net492),
    .D(_01553_),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22085_ (.CLK(net493),
    .D(_01554_),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22086_ (.CLK(net494),
    .D(_01555_),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22087_ (.CLK(net495),
    .D(_01556_),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22088_ (.CLK(net496),
    .D(_01557_),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22089_ (.CLK(net497),
    .D(_01558_),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22090_ (.CLK(net498),
    .D(_01559_),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22091_ (.CLK(net499),
    .D(_01560_),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22092_ (.CLK(net500),
    .D(_01561_),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22093_ (.CLK(net501),
    .D(_01562_),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22094_ (.CLK(net502),
    .D(_01563_),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22095_ (.CLK(net503),
    .D(_01564_),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22096_ (.CLK(net504),
    .D(_01565_),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22097_ (.CLK(net505),
    .D(_01566_),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22098_ (.CLK(net506),
    .D(_01567_),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22099_ (.CLK(net507),
    .D(_01568_),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22100_ (.CLK(net508),
    .D(_01569_),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22101_ (.CLK(net509),
    .D(_01570_),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22102_ (.CLK(net510),
    .D(_01571_),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22103_ (.CLK(net511),
    .D(_01572_),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22104_ (.CLK(net512),
    .D(_01573_),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22105_ (.CLK(net133),
    .D(_01574_),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22106_ (.CLK(net134),
    .D(_01575_),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22107_ (.CLK(net135),
    .D(_01576_),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22108_ (.CLK(net136),
    .D(_01577_),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22109_ (.CLK(net137),
    .D(_01578_),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22110_ (.CLK(net138),
    .D(_01579_),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22111_ (.CLK(net139),
    .D(_01580_),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22112_ (.CLK(net140),
    .D(_01581_),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22113_ (.CLK(net141),
    .D(_01582_),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22114_ (.CLK(net142),
    .D(_01583_),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22115_ (.CLK(net143),
    .D(_01584_),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22116_ (.CLK(net144),
    .D(_01585_),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22117_ (.CLK(net145),
    .D(_01586_),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22118_ (.CLK(net146),
    .D(_01587_),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22119_ (.CLK(net147),
    .D(_01588_),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22120_ (.CLK(net148),
    .D(_01589_),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22121_ (.CLK(net149),
    .D(_01590_),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22122_ (.CLK(net150),
    .D(_01591_),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22123_ (.CLK(net151),
    .D(_01592_),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22124_ (.CLK(net152),
    .D(_01593_),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22125_ (.CLK(net129),
    .D(_01594_),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22126_ (.CLK(net130),
    .D(_01595_),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22127_ (.CLK(net131),
    .D(_01596_),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22128_ (.CLK(net132),
    .D(_01597_),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22129_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01598_),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22130_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01599_),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22131_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01600_),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _22132_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01601_),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _22133_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01602_),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22134_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01603_),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22135_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01604_),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22136_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01605_),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22137_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01606_),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _22138_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01607_),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _22139_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01608_),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _22140_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01609_),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _22141_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01610_),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _22142_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01611_),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22143_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01612_),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22144_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01613_),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22145_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01614_),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22146_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01615_),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22147_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01616_),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22148_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01617_),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22149_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01618_),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22150_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01619_),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22151_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01620_),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22152_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01621_),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22153_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01622_),
    .Q(\rbzero.trace_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22154_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01623_),
    .Q(\rbzero.trace_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22155_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01624_),
    .Q(\rbzero.trace_state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _22156_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01625_),
    .Q(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22157_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01626_),
    .Q(\reg_gpout[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22158_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01627_),
    .Q(\reg_gpout[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22159_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01628_),
    .Q(\reg_gpout[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22160_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01629_),
    .Q(\reg_gpout[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22161_ (.CLK(clknet_leaf_49_i_clk),
    .D(_01630_),
    .Q(\reg_gpout[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22162_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01631_),
    .Q(\reg_gpout[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22163_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01632_),
    .Q(reg_hsync));
 sky130_fd_sc_hd__dfxtp_1 _22164_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01633_),
    .Q(reg_vsync));
 sky130_fd_sc_hd__dfxtp_1 _22165_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01634_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22166_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01635_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22167_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01636_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22168_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01637_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22169_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01638_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22170_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01639_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22171_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01640_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22172_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01641_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22173_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01642_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22174_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01643_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22175_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01644_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22176_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01645_),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22177_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01646_),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22178_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01647_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22179_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01648_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22180_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01649_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22181_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01650_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22182_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01651_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22183_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01652_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22184_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01653_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22185_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01654_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22186_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01655_),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22187_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01656_),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22188_ (.CLK(clknet_leaf_49_i_clk),
    .D(_01657_),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22189_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01658_),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22190_ (.CLK(clknet_leaf_49_i_clk),
    .D(_01659_),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22191_ (.CLK(clknet_leaf_49_i_clk),
    .D(_01660_),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22192_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01661_),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22193_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01662_),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.HI(net111));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_122 (.HI(net122));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_124 (.HI(net124));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_125 (.HI(net125));
 sky130_fd_sc_hd__inv_2 _11504__1 (.A(clknet_opt_3_1_i_clk),
    .Y(net126));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.HI(net110));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(i_debug_map_overlay),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(i_debug_trace_overlay),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(i_debug_vec_overlay),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(i_gpout0_sel[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(i_gpout0_sel[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(i_gpout0_sel[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(i_gpout0_sel[3]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(i_gpout0_sel[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(i_gpout0_sel[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(i_gpout1_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__buf_6 input11 (.A(i_gpout1_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(i_gpout1_sel[2]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(i_gpout1_sel[3]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(i_gpout1_sel[4]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(i_gpout1_sel[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_8 input16 (.A(i_gpout2_sel[0]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(i_gpout2_sel[1]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(i_gpout2_sel[2]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(i_gpout2_sel[3]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(i_gpout2_sel[4]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(i_gpout2_sel[5]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(i_gpout3_sel[0]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(i_gpout3_sel[1]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(i_gpout3_sel[2]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(i_gpout3_sel[3]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(i_gpout3_sel[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(i_gpout3_sel[5]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(i_gpout4_sel[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(i_gpout4_sel[1]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input30 (.A(i_gpout4_sel[2]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 input31 (.A(i_gpout4_sel[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(i_gpout4_sel[4]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(i_gpout4_sel[5]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(i_gpout5_sel[0]),
    .X(net34));
 sky130_fd_sc_hd__buf_6 input35 (.A(i_gpout5_sel[1]),
    .X(net35));
 sky130_fd_sc_hd__buf_6 input36 (.A(i_gpout5_sel[2]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(i_gpout5_sel[3]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(i_gpout5_sel[4]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(i_gpout5_sel[5]),
    .X(net39));
 sky130_fd_sc_hd__buf_8 input40 (.A(i_mode[0]),
    .X(net40));
 sky130_fd_sc_hd__buf_8 input41 (.A(i_mode[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 input42 (.A(i_mode[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(i_reg_csb),
    .X(net43));
 sky130_fd_sc_hd__buf_6 input44 (.A(i_reg_mosi),
    .X(net44));
 sky130_fd_sc_hd__buf_6 input45 (.A(i_reg_outs_enb),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input46 (.A(i_reg_sclk),
    .X(net46));
 sky130_fd_sc_hd__buf_6 input47 (.A(i_reset_lock_a),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_reset_lock_b),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(i_test_wb_clk_i),
    .X(net49));
 sky130_fd_sc_hd__buf_6 input50 (.A(i_tex_in[0]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 input51 (.A(i_tex_in[1]),
    .X(net51));
 sky130_fd_sc_hd__buf_6 input52 (.A(i_tex_in[2]),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input53 (.A(i_tex_in[3]),
    .X(net53));
 sky130_fd_sc_hd__buf_6 input54 (.A(i_vec_csb),
    .X(net54));
 sky130_fd_sc_hd__buf_4 input55 (.A(i_vec_mosi),
    .X(net55));
 sky130_fd_sc_hd__buf_6 input56 (.A(i_vec_sclk),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(o_hsync));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(o_reset));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(o_tex_csb));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(o_tex_out0));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net126),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(o_vsync));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_76 (.LO(net76));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_leaf_39_i_clk),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 net99_3 (.A(clknet_leaf_38_i_clk),
    .Y(net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_opt_2_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_opt_4_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_101_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_102_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_103_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_104_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_105_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_i_clk (.A(clknet_opt_6_0_i_clk),
    .X(clknet_leaf_106_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_107_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_108_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_110_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_111_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_i_clk (.A(clknet_opt_5_0_i_clk),
    .X(clknet_leaf_112_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_113_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_114_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_115_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_116_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_117_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_118_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_119_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_120_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_121_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_122_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_123_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_124_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_125_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_126_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_127_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_128_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_129_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_130_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_131_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_132_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_133_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_134_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_135_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_1_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_2_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_1_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_2_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_1_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_2_2_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_1_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_2_3_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_2_0_1_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_2_0_1_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_2_1_1_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_2_1_1_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_2_2_1_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_2_2_1_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_2_3_1_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_2_3_1_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_opt_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_opt_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_1_i_clk (.A(clknet_opt_3_0_i_clk),
    .X(clknet_opt_3_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_0_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_opt_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_0_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_opt_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_0_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_opt_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05775_ (.A(_05775_),
    .X(clknet_0__05775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05775_ (.A(clknet_0__05775_),
    .X(clknet_1_0__leaf__05775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05775_ (.A(clknet_0__05775_),
    .X(clknet_1_1__leaf__05775_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__06050_ (.A(_06050_),
    .X(clknet_0__06050_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__06050_ (.A(clknet_0__06050_),
    .X(clknet_1_0__leaf__06050_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__06050_ (.A(clknet_0__06050_),
    .X(clknet_1_1__leaf__06050_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05825_ (.A(_05825_),
    .X(clknet_0__05825_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05825_ (.A(clknet_0__05825_),
    .X(clknet_1_0__leaf__05825_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05825_ (.A(clknet_0__05825_),
    .X(clknet_1_1__leaf__05825_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03869_ (.A(_03869_),
    .X(clknet_0__03869_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03869_ (.A(clknet_0__03869_),
    .X(clknet_1_0__leaf__03869_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03869_ (.A(clknet_0__03869_),
    .X(clknet_1_1__leaf__03869_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03868_ (.A(_03868_),
    .X(clknet_0__03868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03868_ (.A(clknet_0__03868_),
    .X(clknet_1_0__leaf__03868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03868_ (.A(clknet_0__03868_),
    .X(clknet_1_1__leaf__03868_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03857_ (.A(_03857_),
    .X(clknet_0__03857_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03857_ (.A(clknet_0__03857_),
    .X(clknet_1_0__leaf__03857_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03857_ (.A(clknet_0__03857_),
    .X(clknet_1_1__leaf__03857_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03867_ (.A(_03867_),
    .X(clknet_0__03867_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03867_ (.A(clknet_0__03867_),
    .X(clknet_1_0__leaf__03867_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03867_ (.A(clknet_0__03867_),
    .X(clknet_1_1__leaf__03867_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03866_ (.A(_03866_),
    .X(clknet_0__03866_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03866_ (.A(clknet_0__03866_),
    .X(clknet_1_0__leaf__03866_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03866_ (.A(clknet_0__03866_),
    .X(clknet_1_1__leaf__03866_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03865_ (.A(_03865_),
    .X(clknet_0__03865_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03865_ (.A(clknet_0__03865_),
    .X(clknet_1_0__leaf__03865_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03865_ (.A(clknet_0__03865_),
    .X(clknet_1_1__leaf__03865_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03864_ (.A(_03864_),
    .X(clknet_0__03864_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03864_ (.A(clknet_0__03864_),
    .X(clknet_1_0__leaf__03864_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03864_ (.A(clknet_0__03864_),
    .X(clknet_1_1__leaf__03864_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03863_ (.A(_03863_),
    .X(clknet_0__03863_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03863_ (.A(clknet_0__03863_),
    .X(clknet_1_0__leaf__03863_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03863_ (.A(clknet_0__03863_),
    .X(clknet_1_1__leaf__03863_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03862_ (.A(_03862_),
    .X(clknet_0__03862_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03862_ (.A(clknet_0__03862_),
    .X(clknet_1_0__leaf__03862_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03862_ (.A(clknet_0__03862_),
    .X(clknet_1_1__leaf__03862_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03861_ (.A(_03861_),
    .X(clknet_0__03861_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03861_ (.A(clknet_0__03861_),
    .X(clknet_1_0__leaf__03861_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03861_ (.A(clknet_0__03861_),
    .X(clknet_1_1__leaf__03861_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03860_ (.A(_03860_),
    .X(clknet_0__03860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03860_ (.A(clknet_0__03860_),
    .X(clknet_1_0__leaf__03860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03860_ (.A(clknet_0__03860_),
    .X(clknet_1_1__leaf__03860_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03859_ (.A(_03859_),
    .X(clknet_0__03859_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03859_ (.A(clknet_0__03859_),
    .X(clknet_1_0__leaf__03859_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03859_ (.A(clknet_0__03859_),
    .X(clknet_1_1__leaf__03859_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03858_ (.A(_03858_),
    .X(clknet_0__03858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03858_ (.A(clknet_0__03858_),
    .X(clknet_1_0__leaf__03858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03858_ (.A(clknet_0__03858_),
    .X(clknet_1_1__leaf__03858_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03846_ (.A(_03846_),
    .X(clknet_0__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03846_ (.A(clknet_0__03846_),
    .X(clknet_1_0__leaf__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03846_ (.A(clknet_0__03846_),
    .X(clknet_1_1__leaf__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03856_ (.A(_03856_),
    .X(clknet_0__03856_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03856_ (.A(clknet_0__03856_),
    .X(clknet_1_0__leaf__03856_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03856_ (.A(clknet_0__03856_),
    .X(clknet_1_1__leaf__03856_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03855_ (.A(_03855_),
    .X(clknet_0__03855_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03855_ (.A(clknet_0__03855_),
    .X(clknet_1_0__leaf__03855_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03855_ (.A(clknet_0__03855_),
    .X(clknet_1_1__leaf__03855_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03854_ (.A(_03854_),
    .X(clknet_0__03854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03854_ (.A(clknet_0__03854_),
    .X(clknet_1_0__leaf__03854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03854_ (.A(clknet_0__03854_),
    .X(clknet_1_1__leaf__03854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03853_ (.A(_03853_),
    .X(clknet_0__03853_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03853_ (.A(clknet_0__03853_),
    .X(clknet_1_0__leaf__03853_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03853_ (.A(clknet_0__03853_),
    .X(clknet_1_1__leaf__03853_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03852_ (.A(_03852_),
    .X(clknet_0__03852_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03852_ (.A(clknet_0__03852_),
    .X(clknet_1_0__leaf__03852_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03852_ (.A(clknet_0__03852_),
    .X(clknet_1_1__leaf__03852_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03851_ (.A(_03851_),
    .X(clknet_0__03851_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03851_ (.A(clknet_0__03851_),
    .X(clknet_1_0__leaf__03851_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03851_ (.A(clknet_0__03851_),
    .X(clknet_1_1__leaf__03851_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03850_ (.A(_03850_),
    .X(clknet_0__03850_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03850_ (.A(clknet_0__03850_),
    .X(clknet_1_0__leaf__03850_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03850_ (.A(clknet_0__03850_),
    .X(clknet_1_1__leaf__03850_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03849_ (.A(_03849_),
    .X(clknet_0__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03849_ (.A(clknet_0__03849_),
    .X(clknet_1_0__leaf__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03849_ (.A(clknet_0__03849_),
    .X(clknet_1_1__leaf__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03848_ (.A(_03848_),
    .X(clknet_0__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03848_ (.A(clknet_0__03848_),
    .X(clknet_1_0__leaf__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03848_ (.A(clknet_0__03848_),
    .X(clknet_1_1__leaf__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03847_ (.A(_03847_),
    .X(clknet_0__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03847_ (.A(clknet_0__03847_),
    .X(clknet_1_0__leaf__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03847_ (.A(clknet_0__03847_),
    .X(clknet_1_1__leaf__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03510_ (.A(_03510_),
    .X(clknet_0__03510_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03510_ (.A(clknet_0__03510_),
    .X(clknet_1_0__leaf__03510_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03510_ (.A(clknet_0__03510_),
    .X(clknet_1_1__leaf__03510_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03845_ (.A(_03845_),
    .X(clknet_0__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03845_ (.A(clknet_0__03845_),
    .X(clknet_1_0__leaf__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03845_ (.A(clknet_0__03845_),
    .X(clknet_1_1__leaf__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03844_ (.A(_03844_),
    .X(clknet_0__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03844_ (.A(clknet_0__03844_),
    .X(clknet_1_0__leaf__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03844_ (.A(clknet_0__03844_),
    .X(clknet_1_1__leaf__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03843_ (.A(_03843_),
    .X(clknet_0__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03843_ (.A(clknet_0__03843_),
    .X(clknet_1_0__leaf__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03843_ (.A(clknet_0__03843_),
    .X(clknet_1_1__leaf__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03842_ (.A(_03842_),
    .X(clknet_0__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03842_ (.A(clknet_0__03842_),
    .X(clknet_1_0__leaf__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03842_ (.A(clknet_0__03842_),
    .X(clknet_1_1__leaf__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03841_ (.A(_03841_),
    .X(clknet_0__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03841_ (.A(clknet_0__03841_),
    .X(clknet_1_0__leaf__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03841_ (.A(clknet_0__03841_),
    .X(clknet_1_1__leaf__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03840_ (.A(_03840_),
    .X(clknet_0__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03840_ (.A(clknet_0__03840_),
    .X(clknet_1_0__leaf__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03840_ (.A(clknet_0__03840_),
    .X(clknet_1_1__leaf__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03839_ (.A(_03839_),
    .X(clknet_0__03839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03839_ (.A(clknet_0__03839_),
    .X(clknet_1_0__leaf__03839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03839_ (.A(clknet_0__03839_),
    .X(clknet_1_1__leaf__03839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03838_ (.A(_03838_),
    .X(clknet_0__03838_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03838_ (.A(clknet_0__03838_),
    .X(clknet_1_0__leaf__03838_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03838_ (.A(clknet_0__03838_),
    .X(clknet_1_1__leaf__03838_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03837_ (.A(_03837_),
    .X(clknet_0__03837_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03837_ (.A(clknet_0__03837_),
    .X(clknet_1_0__leaf__03837_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03837_ (.A(clknet_0__03837_),
    .X(clknet_1_1__leaf__03837_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03511_ (.A(_03511_),
    .X(clknet_0__03511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03511_ (.A(clknet_0__03511_),
    .X(clknet_1_0__leaf__03511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03511_ (.A(clknet_0__03511_),
    .X(clknet_1_1__leaf__03511_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03503_ (.A(_03503_),
    .X(clknet_0__03503_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03503_ (.A(clknet_0__03503_),
    .X(clknet_1_0__leaf__03503_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03503_ (.A(clknet_0__03503_),
    .X(clknet_1_1__leaf__03503_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03509_ (.A(_03509_),
    .X(clknet_0__03509_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03509_ (.A(clknet_0__03509_),
    .X(clknet_1_0__leaf__03509_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03509_ (.A(clknet_0__03509_),
    .X(clknet_1_1__leaf__03509_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03508_ (.A(_03508_),
    .X(clknet_0__03508_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03508_ (.A(clknet_0__03508_),
    .X(clknet_1_0__leaf__03508_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03508_ (.A(clknet_0__03508_),
    .X(clknet_1_1__leaf__03508_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03507_ (.A(_03507_),
    .X(clknet_0__03507_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03507_ (.A(clknet_0__03507_),
    .X(clknet_1_0__leaf__03507_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03507_ (.A(clknet_0__03507_),
    .X(clknet_1_1__leaf__03507_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03506_ (.A(_03506_),
    .X(clknet_0__03506_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03506_ (.A(clknet_0__03506_),
    .X(clknet_1_0__leaf__03506_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03506_ (.A(clknet_0__03506_),
    .X(clknet_1_1__leaf__03506_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03505_ (.A(_03505_),
    .X(clknet_0__03505_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03505_ (.A(clknet_0__03505_),
    .X(clknet_1_0__leaf__03505_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03505_ (.A(clknet_0__03505_),
    .X(clknet_1_1__leaf__03505_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03504_ (.A(_03504_),
    .X(clknet_0__03504_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03504_ (.A(clknet_0__03504_),
    .X(clknet_1_0__leaf__03504_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03504_ (.A(clknet_0__03504_),
    .X(clknet_1_1__leaf__03504_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__06001_ (.A(_06001_),
    .X(clknet_0__06001_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__06001_ (.A(clknet_0__06001_),
    .X(clknet_1_0__leaf__06001_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__06001_ (.A(clknet_0__06001_),
    .X(clknet_1_1__leaf__06001_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05942_ (.A(_05942_),
    .X(clknet_0__05942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05942_ (.A(clknet_0__05942_),
    .X(clknet_1_0__leaf__05942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05942_ (.A(clknet_0__05942_),
    .X(clknet_1_1__leaf__05942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05887_ (.A(_05887_),
    .X(clknet_0__05887_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05887_ (.A(clknet_0__05887_),
    .X(clknet_1_0__leaf__05887_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05887_ (.A(clknet_0__05887_),
    .X(clknet_1_1__leaf__05887_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05832_ (.A(_05832_),
    .X(clknet_0__05832_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05832_ (.A(clknet_0__05832_),
    .X(clknet_1_0__leaf__05832_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05832_ (.A(clknet_0__05832_),
    .X(clknet_1_1__leaf__05832_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rbzero.tex_r1[40] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\rbzero.spi_registers.new_mapd[4] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\rbzero.texu_hot[2] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\rbzero.texu_hot[3] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\rbzero.texu_hot[4] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\rbzero.spi_registers.new_mapd[10] ),
    .X(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01902_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02768_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_03139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_05711_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_05712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_08078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_08090_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_08201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_08201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_08201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_08201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_09691_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_09828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_06163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_06420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_08194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_09831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_09878_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net49));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_980 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1171 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1247 ();
 assign o_rgb[0] = net76;
 assign o_rgb[10] = net84;
 assign o_rgb[11] = net85;
 assign o_rgb[12] = net86;
 assign o_rgb[13] = net87;
 assign o_rgb[16] = net88;
 assign o_rgb[17] = net89;
 assign o_rgb[18] = net90;
 assign o_rgb[19] = net91;
 assign o_rgb[1] = net77;
 assign o_rgb[20] = net92;
 assign o_rgb[21] = net93;
 assign o_rgb[2] = net78;
 assign o_rgb[3] = net79;
 assign o_rgb[4] = net80;
 assign o_rgb[5] = net81;
 assign o_rgb[8] = net82;
 assign o_rgb[9] = net83;
 assign ones[0] = net110;
 assign ones[10] = net120;
 assign ones[11] = net121;
 assign ones[12] = net122;
 assign ones[13] = net123;
 assign ones[14] = net124;
 assign ones[15] = net125;
 assign ones[1] = net111;
 assign ones[2] = net112;
 assign ones[3] = net113;
 assign ones[4] = net114;
 assign ones[5] = net115;
 assign ones[6] = net116;
 assign ones[7] = net117;
 assign ones[8] = net118;
 assign ones[9] = net119;
 assign zeros[0] = net94;
 assign zeros[10] = net104;
 assign zeros[11] = net105;
 assign zeros[12] = net106;
 assign zeros[13] = net107;
 assign zeros[14] = net108;
 assign zeros[15] = net109;
 assign zeros[1] = net95;
 assign zeros[2] = net96;
 assign zeros[3] = net97;
 assign zeros[4] = net98;
 assign zeros[5] = net99;
 assign zeros[6] = net100;
 assign zeros[7] = net101;
 assign zeros[8] = net102;
 assign zeros[9] = net103;
endmodule

