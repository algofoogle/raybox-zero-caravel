magic
tech sky130A
magscale 1 2
timestamp 1698855527
<< nwell >>
rect 1066 116677 116418 116998
rect 1066 115589 116418 116155
rect 1066 114501 116418 115067
rect 1066 113413 116418 113979
rect 1066 112325 116418 112891
rect 1066 111237 116418 111803
rect 1066 110149 116418 110715
rect 1066 109061 116418 109627
rect 1066 107973 116418 108539
rect 1066 106885 116418 107451
rect 1066 105797 116418 106363
rect 1066 104709 116418 105275
rect 1066 103621 116418 104187
rect 1066 102533 116418 103099
rect 1066 101445 116418 102011
rect 1066 100357 116418 100923
rect 1066 99269 116418 99835
rect 1066 98181 116418 98747
rect 1066 97093 116418 97659
rect 1066 96005 116418 96571
rect 1066 94917 116418 95483
rect 1066 93829 116418 94395
rect 1066 92741 116418 93307
rect 1066 91653 116418 92219
rect 1066 90565 116418 91131
rect 1066 89477 116418 90043
rect 1066 88389 116418 88955
rect 1066 87301 116418 87867
rect 1066 86213 116418 86779
rect 1066 85125 116418 85691
rect 1066 84037 116418 84603
rect 1066 82949 116418 83515
rect 1066 81861 116418 82427
rect 1066 80773 116418 81339
rect 1066 79685 116418 80251
rect 1066 78597 116418 79163
rect 1066 77509 116418 78075
rect 1066 76421 116418 76987
rect 1066 75333 116418 75899
rect 1066 74245 116418 74811
rect 1066 73157 116418 73723
rect 1066 72069 116418 72635
rect 1066 70981 116418 71547
rect 1066 69893 116418 70459
rect 1066 68805 116418 69371
rect 1066 67717 116418 68283
rect 1066 66629 116418 67195
rect 1066 65541 116418 66107
rect 1066 64453 116418 65019
rect 1066 63365 116418 63931
rect 1066 62277 116418 62843
rect 1066 61189 116418 61755
rect 1066 60101 116418 60667
rect 1066 59013 116418 59579
rect 1066 57925 116418 58491
rect 1066 56837 116418 57403
rect 1066 55749 116418 56315
rect 1066 54661 116418 55227
rect 1066 53573 116418 54139
rect 1066 52485 116418 53051
rect 1066 51397 116418 51963
rect 1066 50309 116418 50875
rect 1066 49221 116418 49787
rect 1066 48133 116418 48699
rect 1066 47045 116418 47611
rect 1066 45957 116418 46523
rect 1066 44869 116418 45435
rect 1066 43781 116418 44347
rect 1066 42693 116418 43259
rect 1066 41605 116418 42171
rect 1066 40517 116418 41083
rect 1066 39429 116418 39995
rect 1066 38341 116418 38907
rect 1066 37253 116418 37819
rect 1066 36165 116418 36731
rect 1066 35077 116418 35643
rect 1066 33989 116418 34555
rect 1066 32901 116418 33467
rect 1066 31813 116418 32379
rect 1066 30725 116418 31291
rect 1066 29637 116418 30203
rect 1066 28549 116418 29115
rect 1066 27461 116418 28027
rect 1066 26373 116418 26939
rect 1066 25285 116418 25851
rect 1066 24197 116418 24763
rect 1066 23109 116418 23675
rect 1066 22021 116418 22587
rect 1066 20933 116418 21499
rect 1066 19845 116418 20411
rect 1066 18757 116418 19323
rect 1066 17669 116418 18235
rect 1066 16581 116418 17147
rect 1066 15493 116418 16059
rect 1066 14405 116418 14971
rect 1066 13317 116418 13883
rect 1066 12229 116418 12795
rect 1066 11141 116418 11707
rect 1066 10053 116418 10619
rect 1066 8965 116418 9531
rect 1066 7877 116418 8443
rect 1066 6789 116418 7355
rect 1066 5701 116418 6267
rect 1066 4613 116418 5179
rect 1066 3525 116418 4091
rect 1066 2437 116418 3003
<< obsli1 >>
rect 1104 2159 116380 116977
<< obsm1 >>
rect 1104 1844 116380 117008
<< metal2 >>
rect 1306 118858 1362 119658
rect 3698 118858 3754 119658
rect 6090 118858 6146 119658
rect 8482 118858 8538 119658
rect 10874 118858 10930 119658
rect 13266 118858 13322 119658
rect 15658 118858 15714 119658
rect 18050 118858 18106 119658
rect 20442 118858 20498 119658
rect 22834 118858 22890 119658
rect 25226 118858 25282 119658
rect 27618 118858 27674 119658
rect 30010 118858 30066 119658
rect 32402 118858 32458 119658
rect 34794 118858 34850 119658
rect 37186 118858 37242 119658
rect 39578 118858 39634 119658
rect 41970 118858 42026 119658
rect 44362 118858 44418 119658
rect 46754 118858 46810 119658
rect 49146 118858 49202 119658
rect 51538 118858 51594 119658
rect 53930 118858 53986 119658
rect 56322 118858 56378 119658
rect 58714 118858 58770 119658
rect 61106 118858 61162 119658
rect 63498 118858 63554 119658
rect 65890 118858 65946 119658
rect 68282 118858 68338 119658
rect 70674 118858 70730 119658
rect 73066 118858 73122 119658
rect 75458 118858 75514 119658
rect 77850 118858 77906 119658
rect 80242 118858 80298 119658
rect 82634 118858 82690 119658
rect 85026 118858 85082 119658
rect 87418 118858 87474 119658
rect 89810 118858 89866 119658
rect 92202 118858 92258 119658
rect 94594 118858 94650 119658
rect 96986 118858 97042 119658
rect 99378 118858 99434 119658
rect 101770 118858 101826 119658
rect 104162 118858 104218 119658
rect 106554 118858 106610 119658
rect 108946 118858 109002 119658
rect 111338 118858 111394 119658
rect 113730 118858 113786 119658
rect 116122 118858 116178 119658
rect 2502 0 2558 800
rect 5538 0 5594 800
rect 8574 0 8630 800
rect 11610 0 11666 800
rect 14646 0 14702 800
rect 17682 0 17738 800
rect 20718 0 20774 800
rect 23754 0 23810 800
rect 26790 0 26846 800
rect 29826 0 29882 800
rect 32862 0 32918 800
rect 35898 0 35954 800
rect 38934 0 38990 800
rect 41970 0 42026 800
rect 45006 0 45062 800
rect 48042 0 48098 800
rect 51078 0 51134 800
rect 54114 0 54170 800
rect 57150 0 57206 800
rect 60186 0 60242 800
rect 63222 0 63278 800
rect 66258 0 66314 800
rect 69294 0 69350 800
rect 72330 0 72386 800
rect 75366 0 75422 800
rect 78402 0 78458 800
rect 81438 0 81494 800
rect 84474 0 84530 800
rect 87510 0 87566 800
rect 90546 0 90602 800
rect 93582 0 93638 800
rect 96618 0 96674 800
rect 99654 0 99710 800
rect 102690 0 102746 800
rect 105726 0 105782 800
rect 108762 0 108818 800
rect 111798 0 111854 800
rect 114834 0 114890 800
<< obsm2 >>
rect 1584 118802 3642 118858
rect 3810 118802 6034 118858
rect 6202 118802 8426 118858
rect 8594 118802 10818 118858
rect 10986 118802 13210 118858
rect 13378 118802 15602 118858
rect 15770 118802 17994 118858
rect 18162 118802 20386 118858
rect 20554 118802 22778 118858
rect 22946 118802 25170 118858
rect 25338 118802 27562 118858
rect 27730 118802 29954 118858
rect 30122 118802 32346 118858
rect 32514 118802 34738 118858
rect 34906 118802 37130 118858
rect 37298 118802 39522 118858
rect 39690 118802 41914 118858
rect 42082 118802 44306 118858
rect 44474 118802 46698 118858
rect 46866 118802 49090 118858
rect 49258 118802 51482 118858
rect 51650 118802 53874 118858
rect 54042 118802 56266 118858
rect 56434 118802 58658 118858
rect 58826 118802 61050 118858
rect 61218 118802 63442 118858
rect 63610 118802 65834 118858
rect 66002 118802 68226 118858
rect 68394 118802 70618 118858
rect 70786 118802 73010 118858
rect 73178 118802 75402 118858
rect 75570 118802 77794 118858
rect 77962 118802 80186 118858
rect 80354 118802 82578 118858
rect 82746 118802 84970 118858
rect 85138 118802 87362 118858
rect 87530 118802 89754 118858
rect 89922 118802 92146 118858
rect 92314 118802 94538 118858
rect 94706 118802 96930 118858
rect 97098 118802 99322 118858
rect 99490 118802 101714 118858
rect 101882 118802 104106 118858
rect 104274 118802 106498 118858
rect 106666 118802 108890 118858
rect 109058 118802 111282 118858
rect 111450 118802 113674 118858
rect 113842 118802 116066 118858
rect 1584 856 116176 118802
rect 1584 734 2446 856
rect 2614 734 5482 856
rect 5650 734 8518 856
rect 8686 734 11554 856
rect 11722 734 14590 856
rect 14758 734 17626 856
rect 17794 734 20662 856
rect 20830 734 23698 856
rect 23866 734 26734 856
rect 26902 734 29770 856
rect 29938 734 32806 856
rect 32974 734 35842 856
rect 36010 734 38878 856
rect 39046 734 41914 856
rect 42082 734 44950 856
rect 45118 734 47986 856
rect 48154 734 51022 856
rect 51190 734 54058 856
rect 54226 734 57094 856
rect 57262 734 60130 856
rect 60298 734 63166 856
rect 63334 734 66202 856
rect 66370 734 69238 856
rect 69406 734 72274 856
rect 72442 734 75310 856
rect 75478 734 78346 856
rect 78514 734 81382 856
rect 81550 734 84418 856
rect 84586 734 87454 856
rect 87622 734 90490 856
rect 90658 734 93526 856
rect 93694 734 96562 856
rect 96730 734 99598 856
rect 99766 734 102634 856
rect 102802 734 105670 856
rect 105838 734 108706 856
rect 108874 734 111742 856
rect 111910 734 114778 856
rect 114946 734 116176 856
<< metal3 >>
rect 116714 116832 117514 116952
rect 116714 113976 117514 114096
rect 116714 111120 117514 111240
rect 116714 108264 117514 108384
rect 116714 105408 117514 105528
rect 116714 102552 117514 102672
rect 116714 99696 117514 99816
rect 116714 96840 117514 96960
rect 116714 93984 117514 94104
rect 116714 91128 117514 91248
rect 116714 88272 117514 88392
rect 116714 85416 117514 85536
rect 116714 82560 117514 82680
rect 116714 79704 117514 79824
rect 116714 76848 117514 76968
rect 116714 73992 117514 74112
rect 116714 71136 117514 71256
rect 116714 68280 117514 68400
rect 116714 65424 117514 65544
rect 116714 62568 117514 62688
rect 116714 59712 117514 59832
rect 116714 56856 117514 56976
rect 116714 54000 117514 54120
rect 116714 51144 117514 51264
rect 116714 48288 117514 48408
rect 116714 45432 117514 45552
rect 116714 42576 117514 42696
rect 116714 39720 117514 39840
rect 116714 36864 117514 36984
rect 116714 34008 117514 34128
rect 116714 31152 117514 31272
rect 116714 28296 117514 28416
rect 116714 25440 117514 25560
rect 116714 22584 117514 22704
rect 116714 19728 117514 19848
rect 116714 16872 117514 16992
rect 116714 14016 117514 14136
rect 116714 11160 117514 11280
rect 116714 8304 117514 8424
rect 116714 5448 117514 5568
rect 116714 2592 117514 2712
<< obsm3 >>
rect 4210 116752 116634 116993
rect 4210 114176 116714 116752
rect 4210 113896 116634 114176
rect 4210 111320 116714 113896
rect 4210 111040 116634 111320
rect 4210 108464 116714 111040
rect 4210 108184 116634 108464
rect 4210 105608 116714 108184
rect 4210 105328 116634 105608
rect 4210 102752 116714 105328
rect 4210 102472 116634 102752
rect 4210 99896 116714 102472
rect 4210 99616 116634 99896
rect 4210 97040 116714 99616
rect 4210 96760 116634 97040
rect 4210 94184 116714 96760
rect 4210 93904 116634 94184
rect 4210 91328 116714 93904
rect 4210 91048 116634 91328
rect 4210 88472 116714 91048
rect 4210 88192 116634 88472
rect 4210 85616 116714 88192
rect 4210 85336 116634 85616
rect 4210 82760 116714 85336
rect 4210 82480 116634 82760
rect 4210 79904 116714 82480
rect 4210 79624 116634 79904
rect 4210 77048 116714 79624
rect 4210 76768 116634 77048
rect 4210 74192 116714 76768
rect 4210 73912 116634 74192
rect 4210 71336 116714 73912
rect 4210 71056 116634 71336
rect 4210 68480 116714 71056
rect 4210 68200 116634 68480
rect 4210 65624 116714 68200
rect 4210 65344 116634 65624
rect 4210 62768 116714 65344
rect 4210 62488 116634 62768
rect 4210 59912 116714 62488
rect 4210 59632 116634 59912
rect 4210 57056 116714 59632
rect 4210 56776 116634 57056
rect 4210 54200 116714 56776
rect 4210 53920 116634 54200
rect 4210 51344 116714 53920
rect 4210 51064 116634 51344
rect 4210 48488 116714 51064
rect 4210 48208 116634 48488
rect 4210 45632 116714 48208
rect 4210 45352 116634 45632
rect 4210 42776 116714 45352
rect 4210 42496 116634 42776
rect 4210 39920 116714 42496
rect 4210 39640 116634 39920
rect 4210 37064 116714 39640
rect 4210 36784 116634 37064
rect 4210 34208 116714 36784
rect 4210 33928 116634 34208
rect 4210 31352 116714 33928
rect 4210 31072 116634 31352
rect 4210 28496 116714 31072
rect 4210 28216 116634 28496
rect 4210 25640 116714 28216
rect 4210 25360 116634 25640
rect 4210 22784 116714 25360
rect 4210 22504 116634 22784
rect 4210 19928 116714 22504
rect 4210 19648 116634 19928
rect 4210 17072 116714 19648
rect 4210 16792 116634 17072
rect 4210 14216 116714 16792
rect 4210 13936 116634 14216
rect 4210 11360 116714 13936
rect 4210 11080 116634 11360
rect 4210 8504 116714 11080
rect 4210 8224 116634 8504
rect 4210 5648 116714 8224
rect 4210 5368 116634 5648
rect 4210 2792 116714 5368
rect 4210 2512 116634 2792
rect 4210 2143 116714 2512
<< metal4 >>
rect 4208 2128 4528 117008
rect 19568 2128 19888 117008
rect 34928 2128 35248 117008
rect 50288 2128 50608 117008
rect 65648 2128 65968 117008
rect 81008 2128 81328 117008
rect 96368 2128 96688 117008
rect 111728 2128 112048 117008
<< obsm4 >>
rect 26371 2483 34848 116653
rect 35328 2483 50208 116653
rect 50688 2483 65568 116653
rect 66048 2483 80928 116653
rect 81408 2483 96288 116653
rect 96768 2483 111648 116653
rect 112128 2483 115309 116653
<< labels >>
rlabel metal3 s 116714 2592 117514 2712 6 i_clk
port 1 nsew signal input
rlabel metal3 s 116714 71136 117514 71256 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 116714 51144 117514 51264 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 116714 16872 117514 16992 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 116714 19728 117514 19848 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 116714 22584 117514 22704 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 116714 25440 117514 25560 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 116714 28296 117514 28416 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 116714 31152 117514 31272 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 116714 34008 117514 34128 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 116714 36864 117514 36984 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 116714 39720 117514 39840 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 116714 42576 117514 42696 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 116714 45432 117514 45552 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 116714 48288 117514 48408 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 116714 54000 117514 54120 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 116714 56856 117514 56976 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 116714 59712 117514 59832 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 116714 62568 117514 62688 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 116714 65424 117514 65544 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 116714 68280 117514 68400 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 116714 73992 117514 74112 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 116714 76848 117514 76968 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 116714 79704 117514 79824 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 116714 82560 117514 82680 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 116714 85416 117514 85536 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 116714 88272 117514 88392 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 116714 91128 117514 91248 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 116714 93984 117514 94104 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 116714 96840 117514 96960 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 116714 99696 117514 99816 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 116714 102552 117514 102672 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 116714 105408 117514 105528 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 116714 108264 117514 108384 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 116714 111120 117514 111240 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 116714 113976 117514 114096 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 116714 5448 117514 5568 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 116714 8304 117514 8424 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 116714 11160 117514 11280 6 i_reg_outs_enb
port 47 nsew signal input
rlabel metal3 s 116714 14016 117514 14136 6 i_reg_sclk
port 48 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 i_reset_lock_a
port 49 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 i_reset_lock_b
port 50 nsew signal input
rlabel metal3 s 116714 116832 117514 116952 6 i_spare_0
port 51 nsew signal input
rlabel metal2 s 1306 118858 1362 119658 6 i_spare_1
port 52 nsew signal input
rlabel metal2 s 10874 118858 10930 119658 6 i_tex_in[0]
port 53 nsew signal input
rlabel metal2 s 8482 118858 8538 119658 6 i_tex_in[1]
port 54 nsew signal input
rlabel metal2 s 6090 118858 6146 119658 6 i_tex_in[2]
port 55 nsew signal input
rlabel metal2 s 3698 118858 3754 119658 6 i_tex_in[3]
port 56 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 i_vec_csb
port 57 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 i_vec_mosi
port 58 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 i_vec_sclk
port 59 nsew signal input
rlabel metal2 s 25226 118858 25282 119658 6 o_gpout[0]
port 60 nsew signal output
rlabel metal2 s 22834 118858 22890 119658 6 o_gpout[1]
port 61 nsew signal output
rlabel metal2 s 20442 118858 20498 119658 6 o_gpout[2]
port 62 nsew signal output
rlabel metal2 s 18050 118858 18106 119658 6 o_gpout[3]
port 63 nsew signal output
rlabel metal2 s 15658 118858 15714 119658 6 o_gpout[4]
port 64 nsew signal output
rlabel metal2 s 13266 118858 13322 119658 6 o_gpout[5]
port 65 nsew signal output
rlabel metal2 s 39578 118858 39634 119658 6 o_hsync
port 66 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 o_reset
port 67 nsew signal output
rlabel metal2 s 2502 0 2558 800 6 o_rgb[0]
port 68 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 o_rgb[10]
port 69 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 o_rgb[11]
port 70 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 o_rgb[12]
port 71 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 o_rgb[13]
port 72 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 o_rgb[14]
port 73 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 o_rgb[15]
port 74 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 o_rgb[16]
port 75 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 o_rgb[17]
port 76 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 o_rgb[18]
port 77 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 o_rgb[19]
port 78 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 o_rgb[1]
port 79 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 o_rgb[20]
port 80 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 o_rgb[21]
port 81 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 o_rgb[22]
port 82 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 o_rgb[23]
port 83 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 o_rgb[2]
port 84 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 o_rgb[3]
port 85 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 o_rgb[4]
port 86 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 o_rgb[5]
port 87 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 o_rgb[6]
port 88 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 o_rgb[7]
port 89 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 o_rgb[8]
port 90 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 o_rgb[9]
port 91 nsew signal output
rlabel metal2 s 34794 118858 34850 119658 6 o_tex_csb
port 92 nsew signal output
rlabel metal2 s 32402 118858 32458 119658 6 o_tex_oeb0
port 93 nsew signal output
rlabel metal2 s 30010 118858 30066 119658 6 o_tex_out0
port 94 nsew signal output
rlabel metal2 s 27618 118858 27674 119658 6 o_tex_sclk
port 95 nsew signal output
rlabel metal2 s 37186 118858 37242 119658 6 o_vsync
port 96 nsew signal output
rlabel metal2 s 116122 118858 116178 119658 6 ones[0]
port 97 nsew signal output
rlabel metal2 s 92202 118858 92258 119658 6 ones[10]
port 98 nsew signal output
rlabel metal2 s 89810 118858 89866 119658 6 ones[11]
port 99 nsew signal output
rlabel metal2 s 87418 118858 87474 119658 6 ones[12]
port 100 nsew signal output
rlabel metal2 s 85026 118858 85082 119658 6 ones[13]
port 101 nsew signal output
rlabel metal2 s 82634 118858 82690 119658 6 ones[14]
port 102 nsew signal output
rlabel metal2 s 80242 118858 80298 119658 6 ones[15]
port 103 nsew signal output
rlabel metal2 s 113730 118858 113786 119658 6 ones[1]
port 104 nsew signal output
rlabel metal2 s 111338 118858 111394 119658 6 ones[2]
port 105 nsew signal output
rlabel metal2 s 108946 118858 109002 119658 6 ones[3]
port 106 nsew signal output
rlabel metal2 s 106554 118858 106610 119658 6 ones[4]
port 107 nsew signal output
rlabel metal2 s 104162 118858 104218 119658 6 ones[5]
port 108 nsew signal output
rlabel metal2 s 101770 118858 101826 119658 6 ones[6]
port 109 nsew signal output
rlabel metal2 s 99378 118858 99434 119658 6 ones[7]
port 110 nsew signal output
rlabel metal2 s 96986 118858 97042 119658 6 ones[8]
port 111 nsew signal output
rlabel metal2 s 94594 118858 94650 119658 6 ones[9]
port 112 nsew signal output
rlabel metal4 s 4208 2128 4528 117008 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117008 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117008 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117008 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117008 6 vssd1
port 114 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117008 6 vssd1
port 114 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117008 6 vssd1
port 114 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117008 6 vssd1
port 114 nsew ground bidirectional
rlabel metal2 s 77850 118858 77906 119658 6 zeros[0]
port 115 nsew signal output
rlabel metal2 s 53930 118858 53986 119658 6 zeros[10]
port 116 nsew signal output
rlabel metal2 s 51538 118858 51594 119658 6 zeros[11]
port 117 nsew signal output
rlabel metal2 s 49146 118858 49202 119658 6 zeros[12]
port 118 nsew signal output
rlabel metal2 s 46754 118858 46810 119658 6 zeros[13]
port 119 nsew signal output
rlabel metal2 s 44362 118858 44418 119658 6 zeros[14]
port 120 nsew signal output
rlabel metal2 s 41970 118858 42026 119658 6 zeros[15]
port 121 nsew signal output
rlabel metal2 s 75458 118858 75514 119658 6 zeros[1]
port 122 nsew signal output
rlabel metal2 s 73066 118858 73122 119658 6 zeros[2]
port 123 nsew signal output
rlabel metal2 s 70674 118858 70730 119658 6 zeros[3]
port 124 nsew signal output
rlabel metal2 s 68282 118858 68338 119658 6 zeros[4]
port 125 nsew signal output
rlabel metal2 s 65890 118858 65946 119658 6 zeros[5]
port 126 nsew signal output
rlabel metal2 s 63498 118858 63554 119658 6 zeros[6]
port 127 nsew signal output
rlabel metal2 s 61106 118858 61162 119658 6 zeros[7]
port 128 nsew signal output
rlabel metal2 s 58714 118858 58770 119658 6 zeros[8]
port 129 nsew signal output
rlabel metal2 s 56322 118858 56378 119658 6 zeros[9]
port 130 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 117514 119658
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32733700
string GDS_FILE /home/zerotoasic/asic_tools/caravel_user_project/openlane/top_ew_algofoogle/runs/23_11_02_02_43/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1473130
<< end >>

