magic
tech sky130A
magscale 1 2
timestamp 1699028990
<< nwell >>
rect 1066 116677 116602 117243
rect 1066 115589 116602 116155
rect 1066 114501 116602 115067
rect 1066 113413 116602 113979
rect 1066 112325 116602 112891
rect 1066 111237 116602 111803
rect 1066 110149 116602 110715
rect 1066 109061 116602 109627
rect 1066 107973 116602 108539
rect 1066 106885 116602 107451
rect 1066 105797 116602 106363
rect 1066 104709 116602 105275
rect 1066 103621 116602 104187
rect 1066 102533 116602 103099
rect 1066 101445 116602 102011
rect 1066 100357 116602 100923
rect 1066 99269 116602 99835
rect 1066 98181 116602 98747
rect 1066 97093 116602 97659
rect 1066 96005 116602 96571
rect 1066 94917 116602 95483
rect 1066 93829 116602 94395
rect 1066 92741 116602 93307
rect 1066 91653 116602 92219
rect 1066 90565 116602 91131
rect 1066 89477 116602 90043
rect 1066 88389 116602 88955
rect 1066 87301 116602 87867
rect 1066 86213 116602 86779
rect 1066 85125 116602 85691
rect 1066 84037 116602 84603
rect 1066 82949 116602 83515
rect 1066 81861 116602 82427
rect 1066 80773 116602 81339
rect 1066 79685 116602 80251
rect 1066 78597 116602 79163
rect 1066 77509 116602 78075
rect 1066 76421 116602 76987
rect 1066 75333 116602 75899
rect 1066 74245 116602 74811
rect 1066 73157 116602 73723
rect 1066 72069 116602 72635
rect 1066 70981 116602 71547
rect 1066 69893 116602 70459
rect 1066 68805 116602 69371
rect 1066 67717 116602 68283
rect 1066 66629 116602 67195
rect 1066 65541 116602 66107
rect 1066 64453 116602 65019
rect 1066 63365 116602 63931
rect 1066 62277 116602 62843
rect 1066 61189 116602 61755
rect 1066 60101 116602 60667
rect 1066 59013 116602 59579
rect 1066 57925 116602 58491
rect 1066 56837 116602 57403
rect 1066 55749 116602 56315
rect 1066 54661 116602 55227
rect 1066 53573 116602 54139
rect 1066 52485 116602 53051
rect 1066 51397 116602 51963
rect 1066 50309 116602 50875
rect 1066 49221 116602 49787
rect 1066 48133 116602 48699
rect 1066 47045 116602 47611
rect 1066 45957 116602 46523
rect 1066 44869 116602 45435
rect 1066 43781 116602 44347
rect 1066 42693 116602 43259
rect 1066 41605 116602 42171
rect 1066 40517 116602 41083
rect 1066 39429 116602 39995
rect 1066 38341 116602 38907
rect 1066 37253 116602 37819
rect 1066 36165 116602 36731
rect 1066 35077 116602 35643
rect 1066 33989 116602 34555
rect 1066 32901 116602 33467
rect 1066 31813 116602 32379
rect 1066 30725 116602 31291
rect 1066 29637 116602 30203
rect 1066 28549 116602 29115
rect 1066 27461 116602 28027
rect 1066 26373 116602 26939
rect 1066 25285 116602 25851
rect 1066 24197 116602 24763
rect 1066 23109 116602 23675
rect 1066 22021 116602 22587
rect 1066 20933 116602 21499
rect 1066 19845 116602 20411
rect 1066 18757 116602 19323
rect 1066 17669 116602 18235
rect 1066 16581 116602 17147
rect 1066 15493 116602 16059
rect 1066 14405 116602 14971
rect 1066 13317 116602 13883
rect 1066 12229 116602 12795
rect 1066 11141 116602 11707
rect 1066 10053 116602 10619
rect 1066 8965 116602 9531
rect 1066 7877 116602 8443
rect 1066 6789 116602 7355
rect 1066 5701 116602 6267
rect 1066 4613 116602 5179
rect 1066 3525 116602 4091
rect 1066 2437 116602 3003
<< obsli1 >>
rect 1104 2159 116564 117521
<< obsm1 >>
rect 1104 2128 117010 119264
<< metal2 >>
rect 1398 119102 1454 119902
rect 3790 119102 3846 119902
rect 6182 119102 6238 119902
rect 8574 119102 8630 119902
rect 10966 119102 11022 119902
rect 13358 119102 13414 119902
rect 15750 119102 15806 119902
rect 18142 119102 18198 119902
rect 20534 119102 20590 119902
rect 22926 119102 22982 119902
rect 25318 119102 25374 119902
rect 27710 119102 27766 119902
rect 30102 119102 30158 119902
rect 32494 119102 32550 119902
rect 34886 119102 34942 119902
rect 37278 119102 37334 119902
rect 39670 119102 39726 119902
rect 42062 119102 42118 119902
rect 44454 119102 44510 119902
rect 46846 119102 46902 119902
rect 49238 119102 49294 119902
rect 51630 119102 51686 119902
rect 54022 119102 54078 119902
rect 56414 119102 56470 119902
rect 58806 119102 58862 119902
rect 61198 119102 61254 119902
rect 63590 119102 63646 119902
rect 65982 119102 66038 119902
rect 68374 119102 68430 119902
rect 70766 119102 70822 119902
rect 73158 119102 73214 119902
rect 75550 119102 75606 119902
rect 77942 119102 77998 119902
rect 80334 119102 80390 119902
rect 82726 119102 82782 119902
rect 85118 119102 85174 119902
rect 87510 119102 87566 119902
rect 89902 119102 89958 119902
rect 92294 119102 92350 119902
rect 94686 119102 94742 119902
rect 97078 119102 97134 119902
rect 99470 119102 99526 119902
rect 101862 119102 101918 119902
rect 104254 119102 104310 119902
rect 106646 119102 106702 119902
rect 109038 119102 109094 119902
rect 111430 119102 111486 119902
rect 113822 119102 113878 119902
rect 116214 119102 116270 119902
rect 2686 0 2742 800
rect 5722 0 5778 800
rect 8758 0 8814 800
rect 11794 0 11850 800
rect 14830 0 14886 800
rect 17866 0 17922 800
rect 20902 0 20958 800
rect 23938 0 23994 800
rect 26974 0 27030 800
rect 30010 0 30066 800
rect 33046 0 33102 800
rect 36082 0 36138 800
rect 39118 0 39174 800
rect 42154 0 42210 800
rect 45190 0 45246 800
rect 48226 0 48282 800
rect 51262 0 51318 800
rect 54298 0 54354 800
rect 57334 0 57390 800
rect 60370 0 60426 800
rect 63406 0 63462 800
rect 66442 0 66498 800
rect 69478 0 69534 800
rect 72514 0 72570 800
rect 75550 0 75606 800
rect 78586 0 78642 800
rect 81622 0 81678 800
rect 84658 0 84714 800
rect 87694 0 87750 800
rect 90730 0 90786 800
rect 93766 0 93822 800
rect 96802 0 96858 800
rect 99838 0 99894 800
rect 102874 0 102930 800
rect 105910 0 105966 800
rect 108946 0 109002 800
rect 111982 0 112038 800
rect 115018 0 115074 800
<< obsm2 >>
rect 2700 119046 3734 119270
rect 3902 119046 6126 119270
rect 6294 119046 8518 119270
rect 8686 119046 10910 119270
rect 11078 119046 13302 119270
rect 13470 119046 15694 119270
rect 15862 119046 18086 119270
rect 18254 119046 20478 119270
rect 20646 119046 22870 119270
rect 23038 119046 25262 119270
rect 25430 119046 27654 119270
rect 27822 119046 30046 119270
rect 30214 119046 32438 119270
rect 32606 119046 34830 119270
rect 34998 119046 37222 119270
rect 37390 119046 39614 119270
rect 39782 119046 42006 119270
rect 42174 119046 44398 119270
rect 44566 119046 46790 119270
rect 46958 119046 49182 119270
rect 49350 119046 51574 119270
rect 51742 119046 53966 119270
rect 54134 119046 56358 119270
rect 56526 119046 58750 119270
rect 58918 119046 61142 119270
rect 61310 119046 63534 119270
rect 63702 119046 65926 119270
rect 66094 119046 68318 119270
rect 68486 119046 70710 119270
rect 70878 119046 73102 119270
rect 73270 119046 75494 119270
rect 75662 119046 77886 119270
rect 78054 119046 80278 119270
rect 80446 119046 82670 119270
rect 82838 119046 85062 119270
rect 85230 119046 87454 119270
rect 87622 119046 89846 119270
rect 90014 119046 92238 119270
rect 92406 119046 94630 119270
rect 94798 119046 97022 119270
rect 97190 119046 99414 119270
rect 99582 119046 101806 119270
rect 101974 119046 104198 119270
rect 104366 119046 106590 119270
rect 106758 119046 108982 119270
rect 109150 119046 111374 119270
rect 111542 119046 113766 119270
rect 113934 119046 116158 119270
rect 116326 119046 117004 119270
rect 2700 856 117004 119046
rect 2798 734 5666 856
rect 5834 734 8702 856
rect 8870 734 11738 856
rect 11906 734 14774 856
rect 14942 734 17810 856
rect 17978 734 20846 856
rect 21014 734 23882 856
rect 24050 734 26918 856
rect 27086 734 29954 856
rect 30122 734 32990 856
rect 33158 734 36026 856
rect 36194 734 39062 856
rect 39230 734 42098 856
rect 42266 734 45134 856
rect 45302 734 48170 856
rect 48338 734 51206 856
rect 51374 734 54242 856
rect 54410 734 57278 856
rect 57446 734 60314 856
rect 60482 734 63350 856
rect 63518 734 66386 856
rect 66554 734 69422 856
rect 69590 734 72458 856
rect 72626 734 75494 856
rect 75662 734 78530 856
rect 78698 734 81566 856
rect 81734 734 84602 856
rect 84770 734 87638 856
rect 87806 734 90674 856
rect 90842 734 93710 856
rect 93878 734 96746 856
rect 96914 734 99782 856
rect 99950 734 102818 856
rect 102986 734 105854 856
rect 106022 734 108890 856
rect 109058 734 111926 856
rect 112094 734 114962 856
rect 115130 734 117004 856
<< metal3 >>
rect 116958 114248 117758 114368
rect 116958 111528 117758 111648
rect 116958 108808 117758 108928
rect 116958 106088 117758 106208
rect 116958 103368 117758 103488
rect 116958 100648 117758 100768
rect 116958 97928 117758 98048
rect 116958 95208 117758 95328
rect 116958 92488 117758 92608
rect 116958 89768 117758 89888
rect 116958 87048 117758 87168
rect 116958 84328 117758 84448
rect 116958 81608 117758 81728
rect 116958 78888 117758 79008
rect 116958 76168 117758 76288
rect 116958 73448 117758 73568
rect 116958 70728 117758 70848
rect 116958 68008 117758 68128
rect 116958 65288 117758 65408
rect 116958 62568 117758 62688
rect 116958 59848 117758 59968
rect 116958 57128 117758 57248
rect 116958 54408 117758 54528
rect 116958 51688 117758 51808
rect 116958 48968 117758 49088
rect 116958 46248 117758 46368
rect 116958 43528 117758 43648
rect 116958 40808 117758 40928
rect 116958 38088 117758 38208
rect 116958 35368 117758 35488
rect 116958 32648 117758 32768
rect 116958 29928 117758 30048
rect 116958 27208 117758 27328
rect 116958 24488 117758 24608
rect 116958 21768 117758 21888
rect 116958 19048 117758 19168
rect 116958 16328 117758 16448
rect 116958 13608 117758 13728
rect 116958 10888 117758 11008
rect 116958 8168 117758 8288
rect 116958 5448 117758 5568
<< obsm3 >>
rect 3509 114448 116958 117741
rect 3509 114168 116878 114448
rect 3509 111728 116958 114168
rect 3509 111448 116878 111728
rect 3509 109008 116958 111448
rect 3509 108728 116878 109008
rect 3509 106288 116958 108728
rect 3509 106008 116878 106288
rect 3509 103568 116958 106008
rect 3509 103288 116878 103568
rect 3509 100848 116958 103288
rect 3509 100568 116878 100848
rect 3509 98128 116958 100568
rect 3509 97848 116878 98128
rect 3509 95408 116958 97848
rect 3509 95128 116878 95408
rect 3509 92688 116958 95128
rect 3509 92408 116878 92688
rect 3509 89968 116958 92408
rect 3509 89688 116878 89968
rect 3509 87248 116958 89688
rect 3509 86968 116878 87248
rect 3509 84528 116958 86968
rect 3509 84248 116878 84528
rect 3509 81808 116958 84248
rect 3509 81528 116878 81808
rect 3509 79088 116958 81528
rect 3509 78808 116878 79088
rect 3509 76368 116958 78808
rect 3509 76088 116878 76368
rect 3509 73648 116958 76088
rect 3509 73368 116878 73648
rect 3509 70928 116958 73368
rect 3509 70648 116878 70928
rect 3509 68208 116958 70648
rect 3509 67928 116878 68208
rect 3509 65488 116958 67928
rect 3509 65208 116878 65488
rect 3509 62768 116958 65208
rect 3509 62488 116878 62768
rect 3509 60048 116958 62488
rect 3509 59768 116878 60048
rect 3509 57328 116958 59768
rect 3509 57048 116878 57328
rect 3509 54608 116958 57048
rect 3509 54328 116878 54608
rect 3509 51888 116958 54328
rect 3509 51608 116878 51888
rect 3509 49168 116958 51608
rect 3509 48888 116878 49168
rect 3509 46448 116958 48888
rect 3509 46168 116878 46448
rect 3509 43728 116958 46168
rect 3509 43448 116878 43728
rect 3509 41008 116958 43448
rect 3509 40728 116878 41008
rect 3509 38288 116958 40728
rect 3509 38008 116878 38288
rect 3509 35568 116958 38008
rect 3509 35288 116878 35568
rect 3509 32848 116958 35288
rect 3509 32568 116878 32848
rect 3509 30128 116958 32568
rect 3509 29848 116878 30128
rect 3509 27408 116958 29848
rect 3509 27128 116878 27408
rect 3509 24688 116958 27128
rect 3509 24408 116878 24688
rect 3509 21968 116958 24408
rect 3509 21688 116878 21968
rect 3509 19248 116958 21688
rect 3509 18968 116878 19248
rect 3509 16528 116958 18968
rect 3509 16248 116878 16528
rect 3509 13808 116958 16248
rect 3509 13528 116878 13808
rect 3509 11088 116958 13528
rect 3509 10808 116878 11088
rect 3509 8368 116958 10808
rect 3509 8088 116878 8368
rect 3509 5648 116958 8088
rect 3509 5368 116878 5648
rect 3509 2143 116958 5368
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
<< obsm4 >>
rect 6499 2619 19488 116245
rect 19968 2619 34848 116245
rect 35328 2619 50208 116245
rect 50688 2619 65568 116245
rect 66048 2619 80928 116245
rect 81408 2619 96288 116245
rect 96768 2619 111648 116245
rect 112128 2619 114757 116245
<< labels >>
rlabel metal3 s 116958 5448 117758 5568 6 i_clk
port 1 nsew signal input
rlabel metal3 s 116958 70728 117758 70848 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 116958 51688 117758 51808 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 116958 19048 117758 19168 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 116958 21768 117758 21888 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 116958 24488 117758 24608 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 116958 27208 117758 27328 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 116958 29928 117758 30048 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 116958 32648 117758 32768 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 116958 35368 117758 35488 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 116958 38088 117758 38208 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 116958 40808 117758 40928 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 116958 43528 117758 43648 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 116958 46248 117758 46368 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 116958 48968 117758 49088 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 116958 54408 117758 54528 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 116958 57128 117758 57248 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 116958 59848 117758 59968 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 116958 62568 117758 62688 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 116958 65288 117758 65408 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 116958 68008 117758 68128 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 116958 73448 117758 73568 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 116958 76168 117758 76288 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 116958 78888 117758 79008 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 116958 81608 117758 81728 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 116958 84328 117758 84448 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 116958 87048 117758 87168 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 116958 89768 117758 89888 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 116958 92488 117758 92608 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 116958 95208 117758 95328 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 116958 97928 117758 98048 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 116958 100648 117758 100768 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 116958 103368 117758 103488 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 116958 106088 117758 106208 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 116958 108808 117758 108928 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 116958 111528 117758 111648 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 116958 8168 117758 8288 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 116958 10888 117758 11008 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 116958 13608 117758 13728 6 i_reg_outs_enb
port 47 nsew signal input
rlabel metal3 s 116958 16328 117758 16448 6 i_reg_sclk
port 48 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 i_reset_lock_a
port 49 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 i_reset_lock_b
port 50 nsew signal input
rlabel metal3 s 116958 114248 117758 114368 6 i_spare_0
port 51 nsew signal input
rlabel metal2 s 1398 119102 1454 119902 6 i_spare_1
port 52 nsew signal input
rlabel metal2 s 10966 119102 11022 119902 6 i_tex_in[0]
port 53 nsew signal input
rlabel metal2 s 8574 119102 8630 119902 6 i_tex_in[1]
port 54 nsew signal input
rlabel metal2 s 6182 119102 6238 119902 6 i_tex_in[2]
port 55 nsew signal input
rlabel metal2 s 3790 119102 3846 119902 6 i_tex_in[3]
port 56 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 i_vec_csb
port 57 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 i_vec_mosi
port 58 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 i_vec_sclk
port 59 nsew signal input
rlabel metal2 s 25318 119102 25374 119902 6 o_gpout[0]
port 60 nsew signal output
rlabel metal2 s 22926 119102 22982 119902 6 o_gpout[1]
port 61 nsew signal output
rlabel metal2 s 20534 119102 20590 119902 6 o_gpout[2]
port 62 nsew signal output
rlabel metal2 s 18142 119102 18198 119902 6 o_gpout[3]
port 63 nsew signal output
rlabel metal2 s 15750 119102 15806 119902 6 o_gpout[4]
port 64 nsew signal output
rlabel metal2 s 13358 119102 13414 119902 6 o_gpout[5]
port 65 nsew signal output
rlabel metal2 s 39670 119102 39726 119902 6 o_hsync
port 66 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 o_reset
port 67 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 o_rgb[0]
port 68 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 o_rgb[10]
port 69 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 o_rgb[11]
port 70 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 o_rgb[12]
port 71 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 o_rgb[13]
port 72 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 o_rgb[14]
port 73 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 o_rgb[15]
port 74 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 o_rgb[16]
port 75 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 o_rgb[17]
port 76 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 o_rgb[18]
port 77 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 o_rgb[19]
port 78 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 o_rgb[1]
port 79 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 o_rgb[20]
port 80 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 o_rgb[21]
port 81 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 o_rgb[22]
port 82 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 o_rgb[23]
port 83 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 o_rgb[2]
port 84 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 o_rgb[3]
port 85 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 o_rgb[4]
port 86 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 o_rgb[5]
port 87 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 o_rgb[6]
port 88 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 o_rgb[7]
port 89 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 o_rgb[8]
port 90 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 o_rgb[9]
port 91 nsew signal output
rlabel metal2 s 34886 119102 34942 119902 6 o_tex_csb
port 92 nsew signal output
rlabel metal2 s 32494 119102 32550 119902 6 o_tex_oeb0
port 93 nsew signal output
rlabel metal2 s 30102 119102 30158 119902 6 o_tex_out0
port 94 nsew signal output
rlabel metal2 s 27710 119102 27766 119902 6 o_tex_sclk
port 95 nsew signal output
rlabel metal2 s 37278 119102 37334 119902 6 o_vsync
port 96 nsew signal output
rlabel metal2 s 116214 119102 116270 119902 6 ones[0]
port 97 nsew signal output
rlabel metal2 s 92294 119102 92350 119902 6 ones[10]
port 98 nsew signal output
rlabel metal2 s 89902 119102 89958 119902 6 ones[11]
port 99 nsew signal output
rlabel metal2 s 87510 119102 87566 119902 6 ones[12]
port 100 nsew signal output
rlabel metal2 s 85118 119102 85174 119902 6 ones[13]
port 101 nsew signal output
rlabel metal2 s 82726 119102 82782 119902 6 ones[14]
port 102 nsew signal output
rlabel metal2 s 80334 119102 80390 119902 6 ones[15]
port 103 nsew signal output
rlabel metal2 s 113822 119102 113878 119902 6 ones[1]
port 104 nsew signal output
rlabel metal2 s 111430 119102 111486 119902 6 ones[2]
port 105 nsew signal output
rlabel metal2 s 109038 119102 109094 119902 6 ones[3]
port 106 nsew signal output
rlabel metal2 s 106646 119102 106702 119902 6 ones[4]
port 107 nsew signal output
rlabel metal2 s 104254 119102 104310 119902 6 ones[5]
port 108 nsew signal output
rlabel metal2 s 101862 119102 101918 119902 6 ones[6]
port 109 nsew signal output
rlabel metal2 s 99470 119102 99526 119902 6 ones[7]
port 110 nsew signal output
rlabel metal2 s 97078 119102 97134 119902 6 ones[8]
port 111 nsew signal output
rlabel metal2 s 94686 119102 94742 119902 6 ones[9]
port 112 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 113 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 114 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 114 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 114 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 114 nsew ground bidirectional
rlabel metal2 s 77942 119102 77998 119902 6 zeros[0]
port 115 nsew signal output
rlabel metal2 s 54022 119102 54078 119902 6 zeros[10]
port 116 nsew signal output
rlabel metal2 s 51630 119102 51686 119902 6 zeros[11]
port 117 nsew signal output
rlabel metal2 s 49238 119102 49294 119902 6 zeros[12]
port 118 nsew signal output
rlabel metal2 s 46846 119102 46902 119902 6 zeros[13]
port 119 nsew signal output
rlabel metal2 s 44454 119102 44510 119902 6 zeros[14]
port 120 nsew signal output
rlabel metal2 s 42062 119102 42118 119902 6 zeros[15]
port 121 nsew signal output
rlabel metal2 s 75550 119102 75606 119902 6 zeros[1]
port 122 nsew signal output
rlabel metal2 s 73158 119102 73214 119902 6 zeros[2]
port 123 nsew signal output
rlabel metal2 s 70766 119102 70822 119902 6 zeros[3]
port 124 nsew signal output
rlabel metal2 s 68374 119102 68430 119902 6 zeros[4]
port 125 nsew signal output
rlabel metal2 s 65982 119102 66038 119902 6 zeros[5]
port 126 nsew signal output
rlabel metal2 s 63590 119102 63646 119902 6 zeros[6]
port 127 nsew signal output
rlabel metal2 s 61198 119102 61254 119902 6 zeros[7]
port 128 nsew signal output
rlabel metal2 s 58806 119102 58862 119902 6 zeros[8]
port 129 nsew signal output
rlabel metal2 s 56414 119102 56470 119902 6 zeros[9]
port 130 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 117758 119902
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 42283366
string GDS_FILE /home/zerotoasic/asic_tools/raybox-zero-caravel/openlane/top_ew_algofoogle/runs/23_11_04_02_43/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1542014
<< end >>

