// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_outs_enb,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_spare_0,
    i_spare_1,
    i_test_wb_clk_i,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_outs_enb;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_spare_0;
 input i_spare_1;
 input i_test_wb_clk_i;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire _00000_;
 wire _00001_;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire clknet_leaf_0_i_clk;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net77;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net78;
 wire net93;
 wire net94;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net111;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdx[5] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_mapdy[5] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.side_hot ;
 wire \rbzero.spi_registers.got_new_floor ;
 wire \rbzero.spi_registers.got_new_leak ;
 wire \rbzero.spi_registers.got_new_mapd ;
 wire \rbzero.spi_registers.got_new_other ;
 wire \rbzero.spi_registers.got_new_sky ;
 wire \rbzero.spi_registers.got_new_texadd0 ;
 wire \rbzero.spi_registers.got_new_texadd1 ;
 wire \rbzero.spi_registers.got_new_texadd2 ;
 wire \rbzero.spi_registers.got_new_texadd3 ;
 wire \rbzero.spi_registers.got_new_vinf ;
 wire \rbzero.spi_registers.got_new_vshift ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.new_floor[0] ;
 wire \rbzero.spi_registers.new_floor[1] ;
 wire \rbzero.spi_registers.new_floor[2] ;
 wire \rbzero.spi_registers.new_floor[3] ;
 wire \rbzero.spi_registers.new_floor[4] ;
 wire \rbzero.spi_registers.new_floor[5] ;
 wire \rbzero.spi_registers.new_leak[0] ;
 wire \rbzero.spi_registers.new_leak[1] ;
 wire \rbzero.spi_registers.new_leak[2] ;
 wire \rbzero.spi_registers.new_leak[3] ;
 wire \rbzero.spi_registers.new_leak[4] ;
 wire \rbzero.spi_registers.new_leak[5] ;
 wire \rbzero.spi_registers.new_mapd[0] ;
 wire \rbzero.spi_registers.new_mapd[10] ;
 wire \rbzero.spi_registers.new_mapd[11] ;
 wire \rbzero.spi_registers.new_mapd[12] ;
 wire \rbzero.spi_registers.new_mapd[13] ;
 wire \rbzero.spi_registers.new_mapd[14] ;
 wire \rbzero.spi_registers.new_mapd[15] ;
 wire \rbzero.spi_registers.new_mapd[1] ;
 wire \rbzero.spi_registers.new_mapd[2] ;
 wire \rbzero.spi_registers.new_mapd[3] ;
 wire \rbzero.spi_registers.new_mapd[4] ;
 wire \rbzero.spi_registers.new_mapd[5] ;
 wire \rbzero.spi_registers.new_mapd[6] ;
 wire \rbzero.spi_registers.new_mapd[7] ;
 wire \rbzero.spi_registers.new_mapd[8] ;
 wire \rbzero.spi_registers.new_mapd[9] ;
 wire \rbzero.spi_registers.new_other[0] ;
 wire \rbzero.spi_registers.new_other[10] ;
 wire \rbzero.spi_registers.new_other[1] ;
 wire \rbzero.spi_registers.new_other[2] ;
 wire \rbzero.spi_registers.new_other[3] ;
 wire \rbzero.spi_registers.new_other[4] ;
 wire \rbzero.spi_registers.new_other[6] ;
 wire \rbzero.spi_registers.new_other[7] ;
 wire \rbzero.spi_registers.new_other[8] ;
 wire \rbzero.spi_registers.new_other[9] ;
 wire \rbzero.spi_registers.new_sky[0] ;
 wire \rbzero.spi_registers.new_sky[1] ;
 wire \rbzero.spi_registers.new_sky[2] ;
 wire \rbzero.spi_registers.new_sky[3] ;
 wire \rbzero.spi_registers.new_sky[4] ;
 wire \rbzero.spi_registers.new_sky[5] ;
 wire \rbzero.spi_registers.new_texadd0[0] ;
 wire \rbzero.spi_registers.new_texadd0[10] ;
 wire \rbzero.spi_registers.new_texadd0[11] ;
 wire \rbzero.spi_registers.new_texadd0[12] ;
 wire \rbzero.spi_registers.new_texadd0[13] ;
 wire \rbzero.spi_registers.new_texadd0[14] ;
 wire \rbzero.spi_registers.new_texadd0[15] ;
 wire \rbzero.spi_registers.new_texadd0[16] ;
 wire \rbzero.spi_registers.new_texadd0[17] ;
 wire \rbzero.spi_registers.new_texadd0[18] ;
 wire \rbzero.spi_registers.new_texadd0[19] ;
 wire \rbzero.spi_registers.new_texadd0[1] ;
 wire \rbzero.spi_registers.new_texadd0[20] ;
 wire \rbzero.spi_registers.new_texadd0[21] ;
 wire \rbzero.spi_registers.new_texadd0[22] ;
 wire \rbzero.spi_registers.new_texadd0[23] ;
 wire \rbzero.spi_registers.new_texadd0[2] ;
 wire \rbzero.spi_registers.new_texadd0[3] ;
 wire \rbzero.spi_registers.new_texadd0[4] ;
 wire \rbzero.spi_registers.new_texadd0[5] ;
 wire \rbzero.spi_registers.new_texadd0[6] ;
 wire \rbzero.spi_registers.new_texadd0[7] ;
 wire \rbzero.spi_registers.new_texadd0[8] ;
 wire \rbzero.spi_registers.new_texadd0[9] ;
 wire \rbzero.spi_registers.new_texadd1[0] ;
 wire \rbzero.spi_registers.new_texadd1[10] ;
 wire \rbzero.spi_registers.new_texadd1[11] ;
 wire \rbzero.spi_registers.new_texadd1[12] ;
 wire \rbzero.spi_registers.new_texadd1[13] ;
 wire \rbzero.spi_registers.new_texadd1[14] ;
 wire \rbzero.spi_registers.new_texadd1[15] ;
 wire \rbzero.spi_registers.new_texadd1[16] ;
 wire \rbzero.spi_registers.new_texadd1[17] ;
 wire \rbzero.spi_registers.new_texadd1[18] ;
 wire \rbzero.spi_registers.new_texadd1[19] ;
 wire \rbzero.spi_registers.new_texadd1[1] ;
 wire \rbzero.spi_registers.new_texadd1[20] ;
 wire \rbzero.spi_registers.new_texadd1[21] ;
 wire \rbzero.spi_registers.new_texadd1[22] ;
 wire \rbzero.spi_registers.new_texadd1[23] ;
 wire \rbzero.spi_registers.new_texadd1[2] ;
 wire \rbzero.spi_registers.new_texadd1[3] ;
 wire \rbzero.spi_registers.new_texadd1[4] ;
 wire \rbzero.spi_registers.new_texadd1[5] ;
 wire \rbzero.spi_registers.new_texadd1[6] ;
 wire \rbzero.spi_registers.new_texadd1[7] ;
 wire \rbzero.spi_registers.new_texadd1[8] ;
 wire \rbzero.spi_registers.new_texadd1[9] ;
 wire \rbzero.spi_registers.new_texadd2[0] ;
 wire \rbzero.spi_registers.new_texadd2[10] ;
 wire \rbzero.spi_registers.new_texadd2[11] ;
 wire \rbzero.spi_registers.new_texadd2[12] ;
 wire \rbzero.spi_registers.new_texadd2[13] ;
 wire \rbzero.spi_registers.new_texadd2[14] ;
 wire \rbzero.spi_registers.new_texadd2[15] ;
 wire \rbzero.spi_registers.new_texadd2[16] ;
 wire \rbzero.spi_registers.new_texadd2[17] ;
 wire \rbzero.spi_registers.new_texadd2[18] ;
 wire \rbzero.spi_registers.new_texadd2[19] ;
 wire \rbzero.spi_registers.new_texadd2[1] ;
 wire \rbzero.spi_registers.new_texadd2[20] ;
 wire \rbzero.spi_registers.new_texadd2[21] ;
 wire \rbzero.spi_registers.new_texadd2[22] ;
 wire \rbzero.spi_registers.new_texadd2[23] ;
 wire \rbzero.spi_registers.new_texadd2[2] ;
 wire \rbzero.spi_registers.new_texadd2[3] ;
 wire \rbzero.spi_registers.new_texadd2[4] ;
 wire \rbzero.spi_registers.new_texadd2[5] ;
 wire \rbzero.spi_registers.new_texadd2[6] ;
 wire \rbzero.spi_registers.new_texadd2[7] ;
 wire \rbzero.spi_registers.new_texadd2[8] ;
 wire \rbzero.spi_registers.new_texadd2[9] ;
 wire \rbzero.spi_registers.new_texadd3[0] ;
 wire \rbzero.spi_registers.new_texadd3[10] ;
 wire \rbzero.spi_registers.new_texadd3[11] ;
 wire \rbzero.spi_registers.new_texadd3[12] ;
 wire \rbzero.spi_registers.new_texadd3[13] ;
 wire \rbzero.spi_registers.new_texadd3[14] ;
 wire \rbzero.spi_registers.new_texadd3[15] ;
 wire \rbzero.spi_registers.new_texadd3[16] ;
 wire \rbzero.spi_registers.new_texadd3[17] ;
 wire \rbzero.spi_registers.new_texadd3[18] ;
 wire \rbzero.spi_registers.new_texadd3[19] ;
 wire \rbzero.spi_registers.new_texadd3[1] ;
 wire \rbzero.spi_registers.new_texadd3[20] ;
 wire \rbzero.spi_registers.new_texadd3[21] ;
 wire \rbzero.spi_registers.new_texadd3[22] ;
 wire \rbzero.spi_registers.new_texadd3[23] ;
 wire \rbzero.spi_registers.new_texadd3[2] ;
 wire \rbzero.spi_registers.new_texadd3[3] ;
 wire \rbzero.spi_registers.new_texadd3[4] ;
 wire \rbzero.spi_registers.new_texadd3[5] ;
 wire \rbzero.spi_registers.new_texadd3[6] ;
 wire \rbzero.spi_registers.new_texadd3[7] ;
 wire \rbzero.spi_registers.new_texadd3[8] ;
 wire \rbzero.spi_registers.new_texadd3[9] ;
 wire \rbzero.spi_registers.new_vinf ;
 wire \rbzero.spi_registers.new_vshift[0] ;
 wire \rbzero.spi_registers.new_vshift[1] ;
 wire \rbzero.spi_registers.new_vshift[2] ;
 wire \rbzero.spi_registers.new_vshift[3] ;
 wire \rbzero.spi_registers.new_vshift[4] ;
 wire \rbzero.spi_registers.new_vshift[5] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[16] ;
 wire \rbzero.spi_registers.spi_buffer[17] ;
 wire \rbzero.spi_registers.spi_buffer[18] ;
 wire \rbzero.spi_registers.spi_buffer[19] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[20] ;
 wire \rbzero.spi_registers.spi_buffer[21] ;
 wire \rbzero.spi_registers.spi_buffer[22] ;
 wire \rbzero.spi_registers.spi_buffer[23] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.texadd0[0] ;
 wire \rbzero.spi_registers.texadd0[10] ;
 wire \rbzero.spi_registers.texadd0[11] ;
 wire \rbzero.spi_registers.texadd0[12] ;
 wire \rbzero.spi_registers.texadd0[13] ;
 wire \rbzero.spi_registers.texadd0[14] ;
 wire \rbzero.spi_registers.texadd0[15] ;
 wire \rbzero.spi_registers.texadd0[16] ;
 wire \rbzero.spi_registers.texadd0[17] ;
 wire \rbzero.spi_registers.texadd0[18] ;
 wire \rbzero.spi_registers.texadd0[19] ;
 wire \rbzero.spi_registers.texadd0[1] ;
 wire \rbzero.spi_registers.texadd0[20] ;
 wire \rbzero.spi_registers.texadd0[21] ;
 wire \rbzero.spi_registers.texadd0[22] ;
 wire \rbzero.spi_registers.texadd0[23] ;
 wire \rbzero.spi_registers.texadd0[2] ;
 wire \rbzero.spi_registers.texadd0[3] ;
 wire \rbzero.spi_registers.texadd0[4] ;
 wire \rbzero.spi_registers.texadd0[5] ;
 wire \rbzero.spi_registers.texadd0[6] ;
 wire \rbzero.spi_registers.texadd0[7] ;
 wire \rbzero.spi_registers.texadd0[8] ;
 wire \rbzero.spi_registers.texadd0[9] ;
 wire \rbzero.spi_registers.texadd1[0] ;
 wire \rbzero.spi_registers.texadd1[10] ;
 wire \rbzero.spi_registers.texadd1[11] ;
 wire \rbzero.spi_registers.texadd1[12] ;
 wire \rbzero.spi_registers.texadd1[13] ;
 wire \rbzero.spi_registers.texadd1[14] ;
 wire \rbzero.spi_registers.texadd1[15] ;
 wire \rbzero.spi_registers.texadd1[16] ;
 wire \rbzero.spi_registers.texadd1[17] ;
 wire \rbzero.spi_registers.texadd1[18] ;
 wire \rbzero.spi_registers.texadd1[19] ;
 wire \rbzero.spi_registers.texadd1[1] ;
 wire \rbzero.spi_registers.texadd1[20] ;
 wire \rbzero.spi_registers.texadd1[21] ;
 wire \rbzero.spi_registers.texadd1[22] ;
 wire \rbzero.spi_registers.texadd1[23] ;
 wire \rbzero.spi_registers.texadd1[2] ;
 wire \rbzero.spi_registers.texadd1[3] ;
 wire \rbzero.spi_registers.texadd1[4] ;
 wire \rbzero.spi_registers.texadd1[5] ;
 wire \rbzero.spi_registers.texadd1[6] ;
 wire \rbzero.spi_registers.texadd1[7] ;
 wire \rbzero.spi_registers.texadd1[8] ;
 wire \rbzero.spi_registers.texadd1[9] ;
 wire \rbzero.spi_registers.texadd2[0] ;
 wire \rbzero.spi_registers.texadd2[10] ;
 wire \rbzero.spi_registers.texadd2[11] ;
 wire \rbzero.spi_registers.texadd2[12] ;
 wire \rbzero.spi_registers.texadd2[13] ;
 wire \rbzero.spi_registers.texadd2[14] ;
 wire \rbzero.spi_registers.texadd2[15] ;
 wire \rbzero.spi_registers.texadd2[16] ;
 wire \rbzero.spi_registers.texadd2[17] ;
 wire \rbzero.spi_registers.texadd2[18] ;
 wire \rbzero.spi_registers.texadd2[19] ;
 wire \rbzero.spi_registers.texadd2[1] ;
 wire \rbzero.spi_registers.texadd2[20] ;
 wire \rbzero.spi_registers.texadd2[21] ;
 wire \rbzero.spi_registers.texadd2[22] ;
 wire \rbzero.spi_registers.texadd2[23] ;
 wire \rbzero.spi_registers.texadd2[2] ;
 wire \rbzero.spi_registers.texadd2[3] ;
 wire \rbzero.spi_registers.texadd2[4] ;
 wire \rbzero.spi_registers.texadd2[5] ;
 wire \rbzero.spi_registers.texadd2[6] ;
 wire \rbzero.spi_registers.texadd2[7] ;
 wire \rbzero.spi_registers.texadd2[8] ;
 wire \rbzero.spi_registers.texadd2[9] ;
 wire \rbzero.spi_registers.texadd3[0] ;
 wire \rbzero.spi_registers.texadd3[10] ;
 wire \rbzero.spi_registers.texadd3[11] ;
 wire \rbzero.spi_registers.texadd3[12] ;
 wire \rbzero.spi_registers.texadd3[13] ;
 wire \rbzero.spi_registers.texadd3[14] ;
 wire \rbzero.spi_registers.texadd3[15] ;
 wire \rbzero.spi_registers.texadd3[16] ;
 wire \rbzero.spi_registers.texadd3[17] ;
 wire \rbzero.spi_registers.texadd3[18] ;
 wire \rbzero.spi_registers.texadd3[19] ;
 wire \rbzero.spi_registers.texadd3[1] ;
 wire \rbzero.spi_registers.texadd3[20] ;
 wire \rbzero.spi_registers.texadd3[21] ;
 wire \rbzero.spi_registers.texadd3[22] ;
 wire \rbzero.spi_registers.texadd3[23] ;
 wire \rbzero.spi_registers.texadd3[2] ;
 wire \rbzero.spi_registers.texadd3[3] ;
 wire \rbzero.spi_registers.texadd3[4] ;
 wire \rbzero.spi_registers.texadd3[5] ;
 wire \rbzero.spi_registers.texadd3[6] ;
 wire \rbzero.spi_registers.texadd3[7] ;
 wire \rbzero.spi_registers.texadd3[8] ;
 wire \rbzero.spi_registers.texadd3[9] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.texu_hot[0] ;
 wire \rbzero.texu_hot[1] ;
 wire \rbzero.texu_hot[2] ;
 wire \rbzero.texu_hot[3] ;
 wire \rbzero.texu_hot[4] ;
 wire \rbzero.texu_hot[5] ;
 wire \rbzero.trace_state[0] ;
 wire \rbzero.trace_state[1] ;
 wire \rbzero.trace_state[2] ;
 wire \rbzero.trace_state[3] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_hot[0] ;
 wire \rbzero.wall_hot[1] ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \reg_gpout[0] ;
 wire \reg_gpout[1] ;
 wire \reg_gpout[2] ;
 wire \reg_gpout[3] ;
 wire \reg_gpout[4] ;
 wire \reg_gpout[5] ;
 wire reg_hsync;
 wire \reg_rgb[14] ;
 wire \reg_rgb[15] ;
 wire \reg_rgb[22] ;
 wire \reg_rgb[23] ;
 wire \reg_rgb[6] ;
 wire \reg_rgb[7] ;
 wire reg_vsync;
 wire net95;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net129;
 wire net75;
 wire net76;
 wire net127;
 wire net128;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_opt_2_0_i_clk;
 wire clknet_opt_3_0_i_clk;
 wire clknet_opt_4_0_i_clk;
 wire clknet_0__05795_;
 wire clknet_1_0__leaf__05795_;
 wire clknet_1_1__leaf__05795_;
 wire clknet_0__04767_;
 wire clknet_1_0__leaf__04767_;
 wire clknet_1_1__leaf__04767_;
 wire clknet_0__05854_;
 wire clknet_1_0__leaf__05854_;
 wire clknet_1_1__leaf__05854_;
 wire clknet_0__06092_;
 wire clknet_1_0__leaf__06092_;
 wire clknet_1_1__leaf__06092_;
 wire clknet_0__03944_;
 wire clknet_1_0__leaf__03944_;
 wire clknet_1_1__leaf__03944_;
 wire clknet_0__03943_;
 wire clknet_1_0__leaf__03943_;
 wire clknet_1_1__leaf__03943_;
 wire clknet_0__03932_;
 wire clknet_1_0__leaf__03932_;
 wire clknet_1_1__leaf__03932_;
 wire clknet_0__03942_;
 wire clknet_1_0__leaf__03942_;
 wire clknet_1_1__leaf__03942_;
 wire clknet_0__03941_;
 wire clknet_1_0__leaf__03941_;
 wire clknet_1_1__leaf__03941_;
 wire clknet_0__03940_;
 wire clknet_1_0__leaf__03940_;
 wire clknet_1_1__leaf__03940_;
 wire clknet_0__03939_;
 wire clknet_1_0__leaf__03939_;
 wire clknet_1_1__leaf__03939_;
 wire clknet_0__03938_;
 wire clknet_1_0__leaf__03938_;
 wire clknet_1_1__leaf__03938_;
 wire clknet_0__03937_;
 wire clknet_1_0__leaf__03937_;
 wire clknet_1_1__leaf__03937_;
 wire clknet_0__03936_;
 wire clknet_1_0__leaf__03936_;
 wire clknet_1_1__leaf__03936_;
 wire clknet_0__03935_;
 wire clknet_1_0__leaf__03935_;
 wire clknet_1_1__leaf__03935_;
 wire clknet_0__03934_;
 wire clknet_1_0__leaf__03934_;
 wire clknet_1_1__leaf__03934_;
 wire clknet_0__03933_;
 wire clknet_1_0__leaf__03933_;
 wire clknet_1_1__leaf__03933_;
 wire clknet_0__03921_;
 wire clknet_1_0__leaf__03921_;
 wire clknet_1_1__leaf__03921_;
 wire clknet_0__03931_;
 wire clknet_1_0__leaf__03931_;
 wire clknet_1_1__leaf__03931_;
 wire clknet_0__03930_;
 wire clknet_1_0__leaf__03930_;
 wire clknet_1_1__leaf__03930_;
 wire clknet_0__03929_;
 wire clknet_1_0__leaf__03929_;
 wire clknet_1_1__leaf__03929_;
 wire clknet_0__03928_;
 wire clknet_1_0__leaf__03928_;
 wire clknet_1_1__leaf__03928_;
 wire clknet_0__03927_;
 wire clknet_1_0__leaf__03927_;
 wire clknet_1_1__leaf__03927_;
 wire clknet_0__03926_;
 wire clknet_1_0__leaf__03926_;
 wire clknet_1_1__leaf__03926_;
 wire clknet_0__03925_;
 wire clknet_1_0__leaf__03925_;
 wire clknet_1_1__leaf__03925_;
 wire clknet_0__03924_;
 wire clknet_1_0__leaf__03924_;
 wire clknet_1_1__leaf__03924_;
 wire clknet_0__03923_;
 wire clknet_1_0__leaf__03923_;
 wire clknet_1_1__leaf__03923_;
 wire clknet_0__03922_;
 wire clknet_1_0__leaf__03922_;
 wire clknet_1_1__leaf__03922_;
 wire clknet_0__03711_;
 wire clknet_1_0__leaf__03711_;
 wire clknet_1_1__leaf__03711_;
 wire clknet_0__03920_;
 wire clknet_1_0__leaf__03920_;
 wire clknet_1_1__leaf__03920_;
 wire clknet_0__03919_;
 wire clknet_1_0__leaf__03919_;
 wire clknet_1_1__leaf__03919_;
 wire clknet_0__03918_;
 wire clknet_1_0__leaf__03918_;
 wire clknet_1_1__leaf__03918_;
 wire clknet_0__03917_;
 wire clknet_1_0__leaf__03917_;
 wire clknet_1_1__leaf__03917_;
 wire clknet_0__03916_;
 wire clknet_1_0__leaf__03916_;
 wire clknet_1_1__leaf__03916_;
 wire clknet_0__03915_;
 wire clknet_1_0__leaf__03915_;
 wire clknet_1_1__leaf__03915_;
 wire clknet_0__03914_;
 wire clknet_1_0__leaf__03914_;
 wire clknet_1_1__leaf__03914_;
 wire clknet_0__03913_;
 wire clknet_1_0__leaf__03913_;
 wire clknet_1_1__leaf__03913_;
 wire clknet_0__03912_;
 wire clknet_1_0__leaf__03912_;
 wire clknet_1_1__leaf__03912_;
 wire clknet_0__03712_;
 wire clknet_1_0__leaf__03712_;
 wire clknet_1_1__leaf__03712_;
 wire clknet_0__03704_;
 wire clknet_1_0__leaf__03704_;
 wire clknet_1_1__leaf__03704_;
 wire clknet_0__03710_;
 wire clknet_1_0__leaf__03710_;
 wire clknet_1_1__leaf__03710_;
 wire clknet_0__03709_;
 wire clknet_1_0__leaf__03709_;
 wire clknet_1_1__leaf__03709_;
 wire clknet_0__03708_;
 wire clknet_1_0__leaf__03708_;
 wire clknet_1_1__leaf__03708_;
 wire clknet_0__03707_;
 wire clknet_1_0__leaf__03707_;
 wire clknet_1_1__leaf__03707_;
 wire clknet_0__03706_;
 wire clknet_1_0__leaf__03706_;
 wire clknet_1_1__leaf__03706_;
 wire clknet_0__03705_;
 wire clknet_1_0__leaf__03705_;
 wire clknet_1_1__leaf__03705_;
 wire clknet_0__06036_;
 wire clknet_1_0__leaf__06036_;
 wire clknet_1_1__leaf__06036_;
 wire clknet_0__05977_;
 wire clknet_1_0__leaf__05977_;
 wire clknet_1_1__leaf__05977_;
 wire clknet_0__05916_;
 wire clknet_1_0__leaf__05916_;
 wire clknet_1_1__leaf__05916_;
 wire net74;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;

 sky130_fd_sc_hd__buf_4 _10521_ (.A(\gpout0.hpos[0] ),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_4 _10522_ (.A(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_4 _10523_ (.A(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__clkbuf_4 _10524_ (.A(\gpout0.hpos[7] ),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_4 _10525_ (.A(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__xor2_4 _10526_ (.A(net47),
    .B(net48),
    .X(_04108_));
 sky130_fd_sc_hd__buf_4 _10527_ (.A(\gpout0.hpos[8] ),
    .X(_04109_));
 sky130_fd_sc_hd__buf_4 _10528_ (.A(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__buf_4 _10529_ (.A(\gpout0.hpos[9] ),
    .X(_04111_));
 sky130_fd_sc_hd__and2b_1 _10530_ (.A_N(_04110_),
    .B(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__and4_4 _10531_ (.A(_04105_),
    .B(_04107_),
    .C(_04108_),
    .D(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__buf_4 _10532_ (.A(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_4 _10533_ (.A(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(\rbzero.tex_r1[63] ),
    .A1(net50),
    .S(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _10535_ (.A(_04116_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _10536_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[63] ),
    .S(_04115_),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _10537_ (.A(_04117_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_04115_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _10539_ (.A(_04118_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _10540_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(_04115_),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _10541_ (.A(_04119_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _10542_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_04115_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _10543_ (.A(_04120_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _10544_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_04115_),
    .X(_04121_));
 sky130_fd_sc_hd__clkbuf_1 _10545_ (.A(_04121_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_04115_),
    .X(_04122_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_04122_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(_04115_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _10549_ (.A(_04123_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_04115_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _10551_ (.A(_04124_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(_04115_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _10553_ (.A(_04125_),
    .X(_01588_));
 sky130_fd_sc_hd__clkbuf_4 _10554_ (.A(_04114_),
    .X(_04126_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__clkbuf_1 _10556_ (.A(_04127_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _10557_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(_04126_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _10558_ (.A(_04128_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _10559_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_04126_),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_1 _10560_ (.A(_04129_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _10561_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_04126_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _10562_ (.A(_04130_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _10563_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_04126_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _10564_ (.A(_04131_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _10565_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(_04126_),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _10566_ (.A(_04132_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_04126_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _10568_ (.A(_04133_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(_04126_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _10570_ (.A(_04134_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _10571_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_04126_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_1 _10572_ (.A(_04135_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(_04126_),
    .X(_04136_));
 sky130_fd_sc_hd__clkbuf_1 _10574_ (.A(_04136_),
    .X(_01578_));
 sky130_fd_sc_hd__clkbuf_4 _10575_ (.A(_04114_),
    .X(_04137_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__clkbuf_1 _10577_ (.A(_04138_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _10578_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(_04137_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _10579_ (.A(_04139_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _10580_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_04137_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_1 _10581_ (.A(_04140_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(_04137_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _10583_ (.A(_04141_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10584_ (.A0(\rbzero.tex_r1[39] ),
    .A1(net74),
    .S(_04137_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _10585_ (.A(_04142_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(_04137_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _10587_ (.A(_04143_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04137_),
    .X(_04144_));
 sky130_fd_sc_hd__clkbuf_1 _10589_ (.A(_04144_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_04137_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _10591_ (.A(_04145_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _10592_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_04137_),
    .X(_04146_));
 sky130_fd_sc_hd__clkbuf_1 _10593_ (.A(_04146_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(_04137_),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _10595_ (.A(_04147_),
    .X(_01568_));
 sky130_fd_sc_hd__clkbuf_4 _10596_ (.A(_04114_),
    .X(_04148_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_1 _10598_ (.A(_04149_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(_04148_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _10600_ (.A(_04150_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_04148_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_04151_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(_04148_),
    .X(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(_04152_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_04148_),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_04153_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(_04148_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(_04154_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_04148_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _10610_ (.A(_04155_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(_04148_),
    .X(_04156_));
 sky130_fd_sc_hd__clkbuf_1 _10612_ (.A(_04156_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_04148_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_04157_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(_04148_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _10616_ (.A(_04158_),
    .X(_01558_));
 sky130_fd_sc_hd__clkbuf_4 _10617_ (.A(_04114_),
    .X(_04159_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _10619_ (.A(_04160_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(_04159_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _10621_ (.A(_04161_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_04159_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_04162_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(_04159_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_04163_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_04159_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(_04164_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(_04159_),
    .X(_04165_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_04165_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_04159_),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_1 _10631_ (.A(_04166_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(_04159_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_04167_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_04159_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _10635_ (.A(_04168_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(_04159_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _10637_ (.A(_04169_),
    .X(_01548_));
 sky130_fd_sc_hd__clkbuf_4 _10638_ (.A(_04114_),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _10639_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _10640_ (.A(_04171_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_04170_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _10642_ (.A(_04172_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_04170_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(_04173_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(_04170_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(_04174_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_04170_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(_04175_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_04170_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(_04176_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04170_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _10652_ (.A(_04177_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(_04170_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _10654_ (.A(_04178_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04170_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _10656_ (.A(_04179_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(_04170_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _10658_ (.A(_04180_),
    .X(_01538_));
 sky130_fd_sc_hd__clkbuf_4 _10659_ (.A(_04114_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _10661_ (.A(_04182_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_04181_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(_04183_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_04181_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(_04184_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\rbzero.tex_r1[0] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(_04181_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(_04185_),
    .X(_01534_));
 sky130_fd_sc_hd__clkinv_2 _10668_ (.A(_04106_),
    .Y(_04186_));
 sky130_fd_sc_hd__clkinv_4 _10669_ (.A(_04108_),
    .Y(_04187_));
 sky130_fd_sc_hd__or2b_1 _10670_ (.A(_04109_),
    .B_N(\gpout0.hpos[9] ),
    .X(_04188_));
 sky130_fd_sc_hd__or4_4 _10671_ (.A(_04105_),
    .B(_04186_),
    .C(_04187_),
    .D(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__buf_4 _10672_ (.A(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_4 _10673_ (.A(_04190_),
    .X(_04191_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(net50),
    .A1(\rbzero.tex_r0[63] ),
    .S(_04191_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_04192_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04191_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _10677_ (.A(_04193_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_04191_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_04194_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04191_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_04195_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(_04191_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _10683_ (.A(_04196_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04191_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _10685_ (.A(_04197_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10686_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(_04191_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _10687_ (.A(_04198_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04191_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_04199_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(_04191_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _10691_ (.A(_04200_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04191_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _10693_ (.A(_04201_),
    .X(_01524_));
 sky130_fd_sc_hd__clkbuf_4 _10694_ (.A(_04190_),
    .X(_04202_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _10696_ (.A(_04203_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04202_),
    .X(_04204_));
 sky130_fd_sc_hd__clkbuf_1 _10698_ (.A(_04204_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_04202_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(_04205_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_04202_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _10702_ (.A(_04206_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(_04202_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _10704_ (.A(_04207_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10705_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04202_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _10706_ (.A(_04208_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10707_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(_04202_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _10708_ (.A(_04209_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10709_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04202_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _10710_ (.A(_04210_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_04202_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10712_ (.A(_04211_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10713_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04202_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _10714_ (.A(_04212_),
    .X(_01514_));
 sky130_fd_sc_hd__clkbuf_4 _10715_ (.A(_04190_),
    .X(_04213_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _10717_ (.A(_04214_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04213_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _10719_ (.A(_04215_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(_04213_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_04216_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04213_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _10723_ (.A(_04217_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(_04213_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _10725_ (.A(_04218_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04213_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _10727_ (.A(_04219_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10728_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(_04213_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _10729_ (.A(_04220_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04213_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _10731_ (.A(_04221_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(_04213_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _10733_ (.A(_04222_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04213_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _10735_ (.A(_04223_),
    .X(_01504_));
 sky130_fd_sc_hd__clkbuf_4 _10736_ (.A(_04190_),
    .X(_04224_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _10738_ (.A(_04225_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _10739_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _10740_ (.A(_04226_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(_04224_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _10742_ (.A(_04227_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04224_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _10744_ (.A(_04228_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(_04224_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _10746_ (.A(_04229_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10747_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04224_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _10748_ (.A(_04230_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_04224_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _10750_ (.A(_04231_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04224_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _10752_ (.A(_04232_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(_04224_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _10754_ (.A(_04233_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10755_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04224_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _10756_ (.A(_04234_),
    .X(_01494_));
 sky130_fd_sc_hd__clkbuf_4 _10757_ (.A(_04190_),
    .X(_04235_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_04236_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04235_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_04237_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(_04235_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_04238_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04235_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_04239_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(_04235_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(_04240_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04235_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_04241_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(_04235_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _10771_ (.A(_04242_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04235_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _10773_ (.A(_04243_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(_04235_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _10775_ (.A(_04244_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04235_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _10777_ (.A(_04245_),
    .X(_01484_));
 sky130_fd_sc_hd__clkbuf_4 _10778_ (.A(_04190_),
    .X(_04246_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(_04247_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04246_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(_04248_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(_04246_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(_04249_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04246_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_04250_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_04246_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(_04251_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04246_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(_04252_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(_04246_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_04253_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04246_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _10794_ (.A(_04254_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(_04246_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_04255_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04246_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _10798_ (.A(_04256_),
    .X(_01474_));
 sky130_fd_sc_hd__buf_4 _10799_ (.A(_04190_),
    .X(_04257_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _10801_ (.A(_04258_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_04257_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(_04259_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_04257_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(_04260_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04257_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(_04261_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(\rbzero.tex_g1[63] ),
    .A1(net51),
    .S(_04181_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10809_ (.A(_04262_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[63] ),
    .S(_04181_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(_04263_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_04181_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(_04264_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(_04181_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _10815_ (.A(_04265_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04181_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_04266_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_04181_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _10819_ (.A(_04267_),
    .X(_01464_));
 sky130_fd_sc_hd__clkbuf_4 _10820_ (.A(_04114_),
    .X(_04268_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(_04269_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(_04268_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(_04270_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_04268_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_04271_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(_04268_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _10828_ (.A(_04272_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_04268_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_04273_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(_04268_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(_04274_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04268_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_04275_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(_04268_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(_04276_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04268_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(_04277_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_04268_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(_04278_),
    .X(_01454_));
 sky130_fd_sc_hd__buf_4 _10841_ (.A(_04113_),
    .X(_04279_));
 sky130_fd_sc_hd__clkbuf_4 _10842_ (.A(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _10844_ (.A(_04281_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(_04280_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _10846_ (.A(_04282_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_04280_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _10848_ (.A(_04283_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(_04280_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_04284_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_04280_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _10852_ (.A(_04285_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(_04280_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(_04286_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_04280_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_04287_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_04280_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_04288_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_04280_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_04289_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(_04280_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(_04290_),
    .X(_01444_));
 sky130_fd_sc_hd__clkbuf_4 _10863_ (.A(_04279_),
    .X(_04291_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _10865_ (.A(_04292_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(_04291_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(_04293_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_04291_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(_04294_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(_04291_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _10871_ (.A(_04295_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_04291_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_04296_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(_04291_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(_04297_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_04291_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(_04298_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(_04291_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_04299_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_04291_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(_04300_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(_04291_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _10883_ (.A(_04301_),
    .X(_01434_));
 sky130_fd_sc_hd__clkbuf_4 _10884_ (.A(_04279_),
    .X(_04302_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(_04303_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(_04302_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_04304_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_04302_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_04305_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(_04302_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_04306_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04302_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_04307_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(_04302_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(_04308_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_04302_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_04309_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(_04302_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_04310_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04302_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_04311_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(_04302_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_04312_),
    .X(_01424_));
 sky130_fd_sc_hd__clkbuf_4 _10905_ (.A(_04279_),
    .X(_04313_));
 sky130_fd_sc_hd__mux2_1 _10906_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _10907_ (.A(_04314_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _10908_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(_04313_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _10909_ (.A(_04315_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10910_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_04313_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _10911_ (.A(_04316_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _10912_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(_04313_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _10913_ (.A(_04317_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_04313_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _10915_ (.A(_04318_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(_04313_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _10917_ (.A(_04319_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_04313_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _10919_ (.A(_04320_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(_04313_),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_1 _10921_ (.A(_04321_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_04313_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_04322_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(_04313_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_04323_),
    .X(_01414_));
 sky130_fd_sc_hd__buf_4 _10926_ (.A(_04279_),
    .X(_04324_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _10928_ (.A(_04325_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _10929_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(_04324_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _10930_ (.A(_04326_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_04324_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _10932_ (.A(_04327_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10933_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(_04324_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _10934_ (.A(_04328_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_04324_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _10936_ (.A(_04329_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(_04324_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _10938_ (.A(_04330_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10939_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_04324_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _10940_ (.A(_04331_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\rbzero.tex_g1[0] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_04324_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_1 _10942_ (.A(_04332_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(net51),
    .A1(\rbzero.tex_g0[63] ),
    .S(_04257_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(_04333_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_04257_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(_04334_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(_04257_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_04335_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04257_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_04336_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_04257_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _10952_ (.A(_04337_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _10953_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04257_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _10954_ (.A(_04338_),
    .X(_01400_));
 sky130_fd_sc_hd__clkbuf_4 _10955_ (.A(_04190_),
    .X(_04339_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _10957_ (.A(_04340_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_04339_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _10959_ (.A(_04341_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(_04339_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _10961_ (.A(_04342_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04339_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _10963_ (.A(_04343_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(_04339_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _10965_ (.A(_04344_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_04339_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _10967_ (.A(_04345_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(_04339_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_04346_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_04339_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(_04347_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(_04339_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(_04348_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04339_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _10975_ (.A(_04349_),
    .X(_01390_));
 sky130_fd_sc_hd__buf_4 _10976_ (.A(_04189_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_4 _10977_ (.A(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__mux2_1 _10978_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _10979_ (.A(_04352_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _10980_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04351_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _10981_ (.A(_04353_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(_04351_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _10983_ (.A(_04354_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_04351_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(_04355_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(_04351_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _10987_ (.A(_04356_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _10988_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04351_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _10989_ (.A(_04357_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_04351_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _10991_ (.A(_04358_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04351_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _10993_ (.A(_04359_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(_04351_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _10995_ (.A(_04360_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04351_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _10997_ (.A(_04361_),
    .X(_01380_));
 sky130_fd_sc_hd__clkbuf_4 _10998_ (.A(_04350_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _11000_ (.A(_04363_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04362_),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _11002_ (.A(_04364_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(_04362_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(_04365_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04362_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_04366_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(_04362_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _11008_ (.A(_04367_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04362_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _11010_ (.A(_04368_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(_04362_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _11012_ (.A(_04369_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_04362_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_1 _11014_ (.A(_04370_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _11015_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(_04362_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _11016_ (.A(_04371_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04362_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _11018_ (.A(_04372_),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_4 _11019_ (.A(_04350_),
    .X(_04373_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _11021_ (.A(_04374_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_04373_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _11023_ (.A(_04375_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(_04373_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _11025_ (.A(_04376_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_04373_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _11027_ (.A(_04377_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(_04373_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _11029_ (.A(_04378_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04373_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _11031_ (.A(_04379_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(_04373_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _11033_ (.A(_04380_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04373_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _11035_ (.A(_04381_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _11036_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(_04373_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _11037_ (.A(_04382_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_04373_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _11039_ (.A(_04383_),
    .X(_01360_));
 sky130_fd_sc_hd__clkbuf_4 _11040_ (.A(_04350_),
    .X(_04384_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _11042_ (.A(_04385_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04384_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _11044_ (.A(_04386_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(_04384_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _11046_ (.A(_04387_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_04384_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_04388_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(_04384_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _11050_ (.A(_04389_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04384_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _11052_ (.A(_04390_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _11053_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_04384_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _11054_ (.A(_04391_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _11055_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_04384_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _11056_ (.A(_04392_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _11057_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(_04384_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _11058_ (.A(_04393_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _11059_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04384_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _11060_ (.A(_04394_),
    .X(_01350_));
 sky130_fd_sc_hd__buf_4 _11061_ (.A(_04350_),
    .X(_04395_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(_04396_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04395_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(_04397_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(_04395_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(_04398_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04395_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(_04399_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(_04395_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _11071_ (.A(_04400_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_04395_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _11073_ (.A(_04401_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_04395_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _11075_ (.A(_04402_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _11076_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_04395_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _11077_ (.A(_04403_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _11078_ (.A0(\rbzero.tex_b1[63] ),
    .A1(net52),
    .S(_04324_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _11079_ (.A(_04404_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _11080_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[63] ),
    .S(_04324_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _11081_ (.A(_04405_),
    .X(_01340_));
 sky130_fd_sc_hd__clkbuf_4 _11082_ (.A(_04279_),
    .X(_04406_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _11084_ (.A(_04407_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(_04406_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _11086_ (.A(_04408_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04406_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _11088_ (.A(_04409_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(_04406_),
    .X(_04410_));
 sky130_fd_sc_hd__clkbuf_1 _11090_ (.A(_04410_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _11091_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_04406_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _11092_ (.A(_04411_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _11093_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(_04406_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _11094_ (.A(_04412_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _11095_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_04406_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _11096_ (.A(_04413_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _11097_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(_04406_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _11098_ (.A(_04414_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _11099_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04406_),
    .X(_04415_));
 sky130_fd_sc_hd__clkbuf_1 _11100_ (.A(_04415_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _11101_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(_04406_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _11102_ (.A(_04416_),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_4 _11103_ (.A(_04279_),
    .X(_04417_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _11105_ (.A(_04418_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(_04417_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _11107_ (.A(_04419_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04417_),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_1 _11109_ (.A(_04420_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(_04417_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_1 _11111_ (.A(_04421_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04417_),
    .X(_04422_));
 sky130_fd_sc_hd__clkbuf_1 _11113_ (.A(_04422_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _11114_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(_04417_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _11115_ (.A(_04423_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04417_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _11117_ (.A(_04424_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _11118_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(_04417_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _11119_ (.A(_04425_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _11120_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_04417_),
    .X(_04426_));
 sky130_fd_sc_hd__clkbuf_1 _11121_ (.A(_04426_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _11122_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(_04417_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _11123_ (.A(_04427_),
    .X(_01320_));
 sky130_fd_sc_hd__clkbuf_4 _11124_ (.A(_04279_),
    .X(_04428_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _11126_ (.A(_04429_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(_04428_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _11128_ (.A(_04430_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_04428_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(_04431_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _11131_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(_04428_),
    .X(_04432_));
 sky130_fd_sc_hd__clkbuf_1 _11132_ (.A(_04432_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _11133_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04428_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _11134_ (.A(_04433_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _11135_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(_04428_),
    .X(_04434_));
 sky130_fd_sc_hd__clkbuf_1 _11136_ (.A(_04434_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _11137_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_04428_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _11138_ (.A(_04435_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _11139_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(_04428_),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_1 _11140_ (.A(_04436_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _11141_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_04428_),
    .X(_04437_));
 sky130_fd_sc_hd__clkbuf_1 _11142_ (.A(_04437_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _11143_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(_04428_),
    .X(_04438_));
 sky130_fd_sc_hd__clkbuf_1 _11144_ (.A(_04438_),
    .X(_01310_));
 sky130_fd_sc_hd__clkbuf_4 _11145_ (.A(_04279_),
    .X(_04439_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__clkbuf_1 _11147_ (.A(_04440_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(_04439_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _11149_ (.A(_04441_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_04439_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _11151_ (.A(_04442_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_04439_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _11153_ (.A(_04443_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_04439_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(_04444_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(_04439_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _11157_ (.A(_04445_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _11158_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_04439_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _11159_ (.A(_04446_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(_04439_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _11161_ (.A(_04447_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_04439_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _11163_ (.A(_04448_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _11164_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_04439_),
    .X(_04449_));
 sky130_fd_sc_hd__clkbuf_1 _11165_ (.A(_04449_),
    .X(_01300_));
 sky130_fd_sc_hd__clkbuf_4 _11166_ (.A(_04279_),
    .X(_04450_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__clkbuf_1 _11168_ (.A(_04451_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(_04450_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(_04452_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04450_),
    .X(_04453_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(_04453_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(_04450_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _11174_ (.A(_04454_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_04450_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_1 _11176_ (.A(_04455_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _11177_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(_04450_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _11178_ (.A(_04456_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _11179_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04450_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _11180_ (.A(_04457_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _11181_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_04450_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _11182_ (.A(_04458_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04450_),
    .X(_04459_));
 sky130_fd_sc_hd__clkbuf_1 _11184_ (.A(_04459_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _11185_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(_04450_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _11186_ (.A(_04460_),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_4 _11187_ (.A(_04113_),
    .X(_04461_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(_04462_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(_04461_),
    .X(_04463_));
 sky130_fd_sc_hd__clkbuf_1 _11191_ (.A(_04463_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04461_),
    .X(_04464_));
 sky130_fd_sc_hd__clkbuf_1 _11193_ (.A(_04464_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_04461_),
    .X(_04465_));
 sky130_fd_sc_hd__clkbuf_1 _11195_ (.A(_04465_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _11196_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04461_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_1 _11197_ (.A(_04466_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(_04461_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _11199_ (.A(_04467_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04461_),
    .X(_04468_));
 sky130_fd_sc_hd__clkbuf_1 _11201_ (.A(_04468_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _11202_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_04461_),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_1 _11203_ (.A(_04469_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _11204_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04461_),
    .X(_04470_));
 sky130_fd_sc_hd__clkbuf_1 _11205_ (.A(_04470_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _11206_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_04461_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _11207_ (.A(_04471_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _11208_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_04114_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_1 _11209_ (.A(_04472_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _11210_ (.A0(\rbzero.tex_b1[0] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_04114_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _11211_ (.A(_04473_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(net52),
    .A1(\rbzero.tex_b0[63] ),
    .S(_04395_),
    .X(_04474_));
 sky130_fd_sc_hd__clkbuf_1 _11213_ (.A(_04474_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _11214_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_04395_),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_1 _11215_ (.A(_04475_),
    .X(_01185_));
 sky130_fd_sc_hd__clkbuf_4 _11216_ (.A(_04350_),
    .X(_04476_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _11218_ (.A(_04477_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_04476_),
    .X(_04478_));
 sky130_fd_sc_hd__clkbuf_1 _11220_ (.A(_04478_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _11221_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(_04476_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _11222_ (.A(_04479_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _11223_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_04476_),
    .X(_04480_));
 sky130_fd_sc_hd__clkbuf_1 _11224_ (.A(_04480_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _11225_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(_04476_),
    .X(_04481_));
 sky130_fd_sc_hd__clkbuf_1 _11226_ (.A(_04481_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _11227_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_04476_),
    .X(_04482_));
 sky130_fd_sc_hd__clkbuf_1 _11228_ (.A(_04482_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _11229_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(_04476_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _11230_ (.A(_04483_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _11231_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_04476_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _11232_ (.A(_04484_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _11233_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(_04476_),
    .X(_04485_));
 sky130_fd_sc_hd__clkbuf_1 _11234_ (.A(_04485_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _11235_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_04476_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_1 _11236_ (.A(_04486_),
    .X(_01175_));
 sky130_fd_sc_hd__clkbuf_4 _11237_ (.A(_04350_),
    .X(_04487_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__clkbuf_1 _11239_ (.A(_04488_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04487_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_1 _11241_ (.A(_04489_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _11242_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(_04487_),
    .X(_04490_));
 sky130_fd_sc_hd__clkbuf_1 _11243_ (.A(_04490_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_04487_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _11245_ (.A(_04491_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _11246_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(_04487_),
    .X(_04492_));
 sky130_fd_sc_hd__clkbuf_1 _11247_ (.A(_04492_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _11248_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_04487_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_1 _11249_ (.A(_04493_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _11250_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_04487_),
    .X(_04494_));
 sky130_fd_sc_hd__clkbuf_1 _11251_ (.A(_04494_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _11252_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_04487_),
    .X(_04495_));
 sky130_fd_sc_hd__clkbuf_1 _11253_ (.A(_04495_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _11254_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_04487_),
    .X(_04496_));
 sky130_fd_sc_hd__clkbuf_1 _11255_ (.A(_04496_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_04487_),
    .X(_04497_));
 sky130_fd_sc_hd__clkbuf_1 _11257_ (.A(_04497_),
    .X(_01165_));
 sky130_fd_sc_hd__clkbuf_4 _11258_ (.A(_04350_),
    .X(_04498_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__clkbuf_1 _11260_ (.A(_04499_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _11261_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_04498_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_1 _11262_ (.A(_04500_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _11263_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(_04498_),
    .X(_04501_));
 sky130_fd_sc_hd__clkbuf_1 _11264_ (.A(_04501_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _11265_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_04498_),
    .X(_04502_));
 sky130_fd_sc_hd__clkbuf_1 _11266_ (.A(_04502_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _11267_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(_04498_),
    .X(_04503_));
 sky130_fd_sc_hd__clkbuf_1 _11268_ (.A(_04503_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _11269_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04498_),
    .X(_04504_));
 sky130_fd_sc_hd__clkbuf_1 _11270_ (.A(_04504_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _11271_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_04498_),
    .X(_04505_));
 sky130_fd_sc_hd__clkbuf_1 _11272_ (.A(_04505_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _11273_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_04498_),
    .X(_04506_));
 sky130_fd_sc_hd__clkbuf_1 _11274_ (.A(_04506_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _11275_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(_04498_),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_1 _11276_ (.A(_04507_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _11277_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_04498_),
    .X(_04508_));
 sky130_fd_sc_hd__clkbuf_1 _11278_ (.A(_04508_),
    .X(_01155_));
 sky130_fd_sc_hd__clkbuf_4 _11279_ (.A(_04350_),
    .X(_04509_));
 sky130_fd_sc_hd__mux2_1 _11280_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_1 _11281_ (.A(_04510_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _11282_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_04509_),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_1 _11283_ (.A(_04511_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _11284_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(_04509_),
    .X(_04512_));
 sky130_fd_sc_hd__clkbuf_1 _11285_ (.A(_04512_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _11286_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_04509_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_1 _11287_ (.A(_04513_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _11288_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(_04509_),
    .X(_04514_));
 sky130_fd_sc_hd__clkbuf_1 _11289_ (.A(_04514_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _11290_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_04509_),
    .X(_04515_));
 sky130_fd_sc_hd__clkbuf_1 _11291_ (.A(_04515_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _11292_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(_04509_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _11293_ (.A(_04516_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _11294_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04509_),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_1 _11295_ (.A(_04517_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _11296_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(_04509_),
    .X(_04518_));
 sky130_fd_sc_hd__clkbuf_1 _11297_ (.A(_04518_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _11298_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_04509_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _11299_ (.A(_04519_),
    .X(_01145_));
 sky130_fd_sc_hd__clkbuf_4 _11300_ (.A(_04350_),
    .X(_04520_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_1 _11302_ (.A(_04521_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04520_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _11304_ (.A(_04522_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(_04520_),
    .X(_04523_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(_04523_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _11307_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_04520_),
    .X(_04524_));
 sky130_fd_sc_hd__clkbuf_1 _11308_ (.A(_04524_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(_04520_),
    .X(_04525_));
 sky130_fd_sc_hd__clkbuf_1 _11310_ (.A(_04525_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04520_),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_1 _11312_ (.A(_04526_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(_04520_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_1 _11314_ (.A(_04527_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_04520_),
    .X(_04528_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_04528_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _11317_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_04520_),
    .X(_04529_));
 sky130_fd_sc_hd__clkbuf_1 _11318_ (.A(_04529_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_04520_),
    .X(_04530_));
 sky130_fd_sc_hd__clkbuf_1 _11320_ (.A(_04530_),
    .X(_01135_));
 sky130_fd_sc_hd__clkbuf_4 _11321_ (.A(_04189_),
    .X(_04531_));
 sky130_fd_sc_hd__mux2_1 _11322_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__clkbuf_1 _11323_ (.A(_04532_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_04531_),
    .X(_04533_));
 sky130_fd_sc_hd__clkbuf_1 _11325_ (.A(_04533_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _11326_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(_04531_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_1 _11327_ (.A(_04534_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_04531_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _11329_ (.A(_04535_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _11330_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(_04531_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _11331_ (.A(_04536_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_04531_),
    .X(_04537_));
 sky130_fd_sc_hd__clkbuf_1 _11333_ (.A(_04537_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _11334_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(_04531_),
    .X(_04538_));
 sky130_fd_sc_hd__clkbuf_1 _11335_ (.A(_04538_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04531_),
    .X(_04539_));
 sky130_fd_sc_hd__clkbuf_1 _11337_ (.A(_04539_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(_04531_),
    .X(_04540_));
 sky130_fd_sc_hd__clkbuf_1 _11339_ (.A(_04540_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _11340_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_04531_),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_1 _11341_ (.A(_04541_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _11342_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_04190_),
    .X(_04542_));
 sky130_fd_sc_hd__clkbuf_1 _11343_ (.A(_04542_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _11344_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04190_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _11345_ (.A(_04543_),
    .X(_01123_));
 sky130_fd_sc_hd__buf_6 _11346_ (.A(_04187_),
    .X(_04544_));
 sky130_fd_sc_hd__buf_6 _11347_ (.A(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__buf_8 _11348_ (.A(_04545_),
    .X(net64));
 sky130_fd_sc_hd__inv_2 _11349_ (.A(\gpout0.hpos[6] ),
    .Y(_04546_));
 sky130_fd_sc_hd__clkbuf_4 _11350_ (.A(\gpout0.hpos[5] ),
    .X(_04547_));
 sky130_fd_sc_hd__clkinv_4 _11351_ (.A(\gpout0.hpos[3] ),
    .Y(_04548_));
 sky130_fd_sc_hd__clkinv_4 _11352_ (.A(\gpout0.hpos[4] ),
    .Y(_04549_));
 sky130_fd_sc_hd__nor2_2 _11353_ (.A(_04548_),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__nor2_1 _11354_ (.A(_04547_),
    .B(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__o21ai_4 _11355_ (.A1(_04546_),
    .A2(_04551_),
    .B1(_04186_),
    .Y(_04552_));
 sky130_fd_sc_hd__clkbuf_4 _11356_ (.A(\gpout0.hpos[6] ),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_4 _11357_ (.A(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__inv_2 _11358_ (.A(\gpout0.hpos[5] ),
    .Y(_04555_));
 sky130_fd_sc_hd__inv_2 _11359_ (.A(_04550_),
    .Y(_04556_));
 sky130_fd_sc_hd__nor2_1 _11360_ (.A(_04555_),
    .B(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__nor2_1 _11361_ (.A(_04551_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__and4_1 _11362_ (.A(_04186_),
    .B(_04554_),
    .C(\gpout0.hpos[9] ),
    .D(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__a21boi_4 _11363_ (.A1(_04110_),
    .A2(_04552_),
    .B1_N(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__clkinv_4 _11364_ (.A(_04560_),
    .Y(net72));
 sky130_fd_sc_hd__clkbuf_4 _11365_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_04561_));
 sky130_fd_sc_hd__buf_2 _11366_ (.A(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__buf_4 _11367_ (.A(\rbzero.trace_state[2] ),
    .X(_04563_));
 sky130_fd_sc_hd__or2_2 _11368_ (.A(\rbzero.trace_state[1] ),
    .B(\rbzero.trace_state[0] ),
    .X(_04564_));
 sky130_fd_sc_hd__clkinv_2 _11369_ (.A(\rbzero.vga_sync.vsync ),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_8 _11370_ (.A(_04565_),
    .B(_04108_),
    .Y(_04566_));
 sky130_fd_sc_hd__inv_2 _11371_ (.A(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__buf_4 _11372_ (.A(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__o31a_1 _11373_ (.A1(\rbzero.trace_state[3] ),
    .A2(_04563_),
    .A3(_04564_),
    .B1(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__buf_4 _11374_ (.A(\rbzero.trace_state[1] ),
    .X(_04570_));
 sky130_fd_sc_hd__clkbuf_2 _11375_ (.A(\rbzero.trace_state[0] ),
    .X(_04571_));
 sky130_fd_sc_hd__nor2_1 _11376_ (.A(\rbzero.trace_state[3] ),
    .B(_04563_),
    .Y(_04572_));
 sky130_fd_sc_hd__and3_1 _11377_ (.A(_04570_),
    .B(_04571_),
    .C(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__and4bb_1 _11378_ (.A_N(_04563_),
    .B_N(_04570_),
    .C(_04571_),
    .D(\rbzero.trace_state[3] ),
    .X(_04574_));
 sky130_fd_sc_hd__nor2_1 _11379_ (.A(_04573_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__buf_4 _11380_ (.A(_04568_),
    .X(_04576_));
 sky130_fd_sc_hd__a32o_1 _11381_ (.A1(_04562_),
    .A2(_04569_),
    .A3(_04575_),
    .B1(_04573_),
    .B2(_04576_),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_4 _11382_ (.A(_04112_),
    .B(_04552_),
    .Y(net71));
 sky130_fd_sc_hd__buf_2 _11383_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_04577_));
 sky130_fd_sc_hd__buf_2 _11384_ (.A(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__a21bo_1 _11385_ (.A1(_04578_),
    .A2(_04575_),
    .B1_N(_04569_),
    .X(_00000_));
 sky130_fd_sc_hd__inv_6 _11386_ (.A(\gpout0.hpos[2] ),
    .Y(_04579_));
 sky130_fd_sc_hd__nand2_2 _11387_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .Y(_04580_));
 sky130_fd_sc_hd__or2_1 _11388_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .X(_04581_));
 sky130_fd_sc_hd__inv_2 _11389_ (.A(\gpout0.hpos[1] ),
    .Y(_04582_));
 sky130_fd_sc_hd__clkbuf_8 _11390_ (.A(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__a21oi_1 _11391_ (.A1(_04583_),
    .A2(_04105_),
    .B1(_04579_),
    .Y(_04584_));
 sky130_fd_sc_hd__a31o_1 _11392_ (.A1(_04579_),
    .A2(_04580_),
    .A3(_04581_),
    .B1(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__buf_4 _11393_ (.A(\gpout0.hpos[3] ),
    .X(_04586_));
 sky130_fd_sc_hd__buf_2 _11394_ (.A(\gpout0.hpos[4] ),
    .X(_04587_));
 sky130_fd_sc_hd__clkbuf_4 _11395_ (.A(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__buf_4 _11396_ (.A(\gpout0.hpos[2] ),
    .X(_04589_));
 sky130_fd_sc_hd__inv_2 _11397_ (.A(\rbzero.wall_hot[1] ),
    .Y(_04590_));
 sky130_fd_sc_hd__clkbuf_4 _11398_ (.A(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__buf_4 _11399_ (.A(\rbzero.wall_hot[0] ),
    .X(_04592_));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(_04591_),
    .B(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__clkbuf_4 _11401_ (.A(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_4 _11402_ (.A(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__nor2_1 _11403_ (.A(_04590_),
    .B(_04592_),
    .Y(_04596_));
 sky130_fd_sc_hd__clkbuf_4 _11404_ (.A(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_4 _11405_ (.A(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__and2_1 _11406_ (.A(\rbzero.spi_registers.texadd1[23] ),
    .B(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__buf_4 _11407_ (.A(_04591_),
    .X(_04600_));
 sky130_fd_sc_hd__and2_2 _11408_ (.A(\rbzero.wall_hot[1] ),
    .B(\rbzero.wall_hot[0] ),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_4 _11409_ (.A(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__buf_4 _11410_ (.A(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__and2_1 _11411_ (.A(_04590_),
    .B(_04592_),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_4 _11412_ (.A(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__buf_4 _11413_ (.A(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__a221o_1 _11414_ (.A1(\rbzero.spi_registers.texadd3[23] ),
    .A2(_04600_),
    .B1(_04603_),
    .B2(\rbzero.spi_registers.texadd2[23] ),
    .C1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__o22a_1 _11415_ (.A1(\rbzero.spi_registers.texadd0[23] ),
    .A2(_04595_),
    .B1(_04599_),
    .B2(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__a221o_1 _11416_ (.A1(\rbzero.spi_registers.texadd2[22] ),
    .A2(_04592_),
    .B1(_04598_),
    .B2(\rbzero.spi_registers.texadd1[22] ),
    .C1(_04606_),
    .X(_04609_));
 sky130_fd_sc_hd__a21o_1 _11417_ (.A1(\rbzero.spi_registers.texadd3[22] ),
    .A2(_04600_),
    .B1(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__o21ai_1 _11418_ (.A1(\rbzero.spi_registers.texadd0[22] ),
    .A2(_04595_),
    .B1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_1 _11419_ (.A(_04104_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_4 _11420_ (.A(\rbzero.wall_hot[1] ),
    .B(_04592_),
    .Y(_04613_));
 sky130_fd_sc_hd__a22o_1 _11421_ (.A1(\rbzero.spi_registers.texadd2[14] ),
    .A2(_04603_),
    .B1(_04613_),
    .B2(\rbzero.spi_registers.texadd3[14] ),
    .X(_04614_));
 sky130_fd_sc_hd__a22o_1 _11422_ (.A1(\rbzero.spi_registers.texadd3[13] ),
    .A2(_04613_),
    .B1(_04597_),
    .B2(\rbzero.spi_registers.texadd1[13] ),
    .X(_04615_));
 sky130_fd_sc_hd__buf_2 _11423_ (.A(\rbzero.side_hot ),
    .X(_04616_));
 sky130_fd_sc_hd__clkbuf_4 _11424_ (.A(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__buf_4 _11425_ (.A(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__and2_1 _11426_ (.A(\rbzero.spi_registers.texadd1[12] ),
    .B(_04597_),
    .X(_04619_));
 sky130_fd_sc_hd__a221o_1 _11427_ (.A1(\rbzero.spi_registers.texadd3[12] ),
    .A2(_04591_),
    .B1(_04602_),
    .B2(\rbzero.spi_registers.texadd2[12] ),
    .C1(_04605_),
    .X(_04620_));
 sky130_fd_sc_hd__o22a_1 _11428_ (.A1(\rbzero.spi_registers.texadd0[12] ),
    .A2(_04594_),
    .B1(_04619_),
    .B2(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__nand2_1 _11429_ (.A(_04618_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__and2_1 _11430_ (.A(\rbzero.spi_registers.texadd1[11] ),
    .B(_04597_),
    .X(_04623_));
 sky130_fd_sc_hd__a221o_1 _11431_ (.A1(\rbzero.spi_registers.texadd3[11] ),
    .A2(_04591_),
    .B1(_04602_),
    .B2(\rbzero.spi_registers.texadd2[11] ),
    .C1(_04605_),
    .X(_04624_));
 sky130_fd_sc_hd__o22a_1 _11432_ (.A1(\rbzero.spi_registers.texadd0[11] ),
    .A2(_04594_),
    .B1(_04623_),
    .B2(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__nand2_1 _11433_ (.A(\rbzero.texu_hot[5] ),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__and2_1 _11434_ (.A(\rbzero.spi_registers.texadd1[10] ),
    .B(_04597_),
    .X(_04627_));
 sky130_fd_sc_hd__a221o_1 _11435_ (.A1(\rbzero.spi_registers.texadd3[10] ),
    .A2(_04591_),
    .B1(_04602_),
    .B2(\rbzero.spi_registers.texadd2[10] ),
    .C1(_04605_),
    .X(_04628_));
 sky130_fd_sc_hd__o22a_1 _11436_ (.A1(\rbzero.spi_registers.texadd0[10] ),
    .A2(_04594_),
    .B1(_04627_),
    .B2(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _11437_ (.A(\rbzero.texu_hot[4] ),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__and2_1 _11438_ (.A(\rbzero.spi_registers.texadd1[9] ),
    .B(_04596_),
    .X(_04631_));
 sky130_fd_sc_hd__a221o_1 _11439_ (.A1(\rbzero.spi_registers.texadd3[9] ),
    .A2(_04591_),
    .B1(_04601_),
    .B2(\rbzero.spi_registers.texadd2[9] ),
    .C1(_04605_),
    .X(_04632_));
 sky130_fd_sc_hd__o22a_1 _11440_ (.A1(\rbzero.spi_registers.texadd0[9] ),
    .A2(_04594_),
    .B1(_04631_),
    .B2(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__nand2_1 _11441_ (.A(\rbzero.texu_hot[3] ),
    .B(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__and2_1 _11442_ (.A(\rbzero.spi_registers.texadd1[8] ),
    .B(_04596_),
    .X(_04635_));
 sky130_fd_sc_hd__a221o_1 _11443_ (.A1(\rbzero.spi_registers.texadd3[8] ),
    .A2(_04591_),
    .B1(_04601_),
    .B2(\rbzero.spi_registers.texadd2[8] ),
    .C1(_04605_),
    .X(_04636_));
 sky130_fd_sc_hd__o22a_1 _11444_ (.A1(\rbzero.spi_registers.texadd0[8] ),
    .A2(_04593_),
    .B1(_04635_),
    .B2(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__nor2_1 _11445_ (.A(\rbzero.texu_hot[2] ),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__a22o_1 _11446_ (.A1(\rbzero.spi_registers.texadd3[7] ),
    .A2(_04590_),
    .B1(_04601_),
    .B2(\rbzero.spi_registers.texadd2[7] ),
    .X(_04639_));
 sky130_fd_sc_hd__a211o_1 _11447_ (.A1(\rbzero.spi_registers.texadd1[7] ),
    .A2(_04596_),
    .B1(_04604_),
    .C1(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__o21a_1 _11448_ (.A1(\rbzero.spi_registers.texadd0[7] ),
    .A2(_04593_),
    .B1(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__a22o_1 _11449_ (.A1(\rbzero.spi_registers.texadd3[6] ),
    .A2(_04591_),
    .B1(_04601_),
    .B2(\rbzero.spi_registers.texadd2[6] ),
    .X(_04642_));
 sky130_fd_sc_hd__a211o_1 _11450_ (.A1(\rbzero.spi_registers.texadd1[6] ),
    .A2(_04596_),
    .B1(_04605_),
    .C1(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__or2_1 _11451_ (.A(\rbzero.spi_registers.texadd0[6] ),
    .B(_04593_),
    .X(_04644_));
 sky130_fd_sc_hd__nand3_1 _11452_ (.A(\rbzero.texu_hot[0] ),
    .B(_04643_),
    .C(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__xnor2_1 _11453_ (.A(\rbzero.texu_hot[1] ),
    .B(_04641_),
    .Y(_04646_));
 sky130_fd_sc_hd__nor2_1 _11454_ (.A(_04645_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__a21oi_1 _11455_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_04641_),
    .B1(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__and2_1 _11456_ (.A(\rbzero.texu_hot[2] ),
    .B(_04637_),
    .X(_04649_));
 sky130_fd_sc_hd__o21ba_1 _11457_ (.A1(_04638_),
    .A2(_04648_),
    .B1_N(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__or2_1 _11458_ (.A(\rbzero.texu_hot[3] ),
    .B(_04633_),
    .X(_04651_));
 sky130_fd_sc_hd__nand2_1 _11459_ (.A(_04634_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__or2_1 _11460_ (.A(_04650_),
    .B(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__or2_1 _11461_ (.A(\rbzero.texu_hot[4] ),
    .B(_04629_),
    .X(_04654_));
 sky130_fd_sc_hd__nand2_1 _11462_ (.A(_04630_),
    .B(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a21o_1 _11463_ (.A1(_04634_),
    .A2(_04653_),
    .B1(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__or2_1 _11464_ (.A(\rbzero.texu_hot[5] ),
    .B(_04625_),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _11465_ (.A(_04626_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__a21o_1 _11466_ (.A1(_04630_),
    .A2(_04656_),
    .B1(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__or2_1 _11467_ (.A(_04618_),
    .B(_04621_),
    .X(_04660_));
 sky130_fd_sc_hd__nand2_1 _11468_ (.A(_04622_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__a21o_1 _11469_ (.A1(_04626_),
    .A2(_04659_),
    .B1(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__nor2_1 _11470_ (.A(\rbzero.spi_registers.texadd0[13] ),
    .B(_04594_),
    .Y(_04663_));
 sky130_fd_sc_hd__and2b_1 _11471_ (.A_N(\rbzero.spi_registers.texadd2[13] ),
    .B(_04602_),
    .X(_04664_));
 sky130_fd_sc_hd__a2111oi_2 _11472_ (.A1(_04622_),
    .A2(_04662_),
    .B1(_04663_),
    .C1(_04664_),
    .D1(_04615_),
    .Y(_04665_));
 sky130_fd_sc_hd__or2_1 _11473_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_04594_),
    .X(_04666_));
 sky130_fd_sc_hd__or3_1 _11474_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .B(_04591_),
    .C(_04592_),
    .X(_04667_));
 sky130_fd_sc_hd__a22oi_1 _11475_ (.A1(\rbzero.spi_registers.texadd2[14] ),
    .A2(_04602_),
    .B1(_04613_),
    .B2(\rbzero.spi_registers.texadd3[14] ),
    .Y(_04668_));
 sky130_fd_sc_hd__o2111a_1 _11476_ (.A1(_04615_),
    .A2(_04665_),
    .B1(_04666_),
    .C1(_04667_),
    .D1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__a22o_1 _11477_ (.A1(\rbzero.spi_registers.texadd3[15] ),
    .A2(_04591_),
    .B1(_04602_),
    .B2(\rbzero.spi_registers.texadd2[15] ),
    .X(_04670_));
 sky130_fd_sc_hd__a211o_1 _11478_ (.A1(\rbzero.spi_registers.texadd1[15] ),
    .A2(_04597_),
    .B1(_04605_),
    .C1(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__o21a_1 _11479_ (.A1(\rbzero.spi_registers.texadd0[15] ),
    .A2(_04594_),
    .B1(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__o21ai_1 _11480_ (.A1(_04614_),
    .A2(_04669_),
    .B1(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__a22o_1 _11481_ (.A1(\rbzero.spi_registers.texadd3[16] ),
    .A2(_04600_),
    .B1(_04602_),
    .B2(\rbzero.spi_registers.texadd2[16] ),
    .X(_04674_));
 sky130_fd_sc_hd__a211o_1 _11482_ (.A1(\rbzero.spi_registers.texadd1[16] ),
    .A2(_04597_),
    .B1(_04605_),
    .C1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__o21ai_1 _11483_ (.A1(\rbzero.spi_registers.texadd0[16] ),
    .A2(_04594_),
    .B1(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__nor2_1 _11484_ (.A(_04673_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__a22o_1 _11485_ (.A1(\rbzero.spi_registers.texadd3[17] ),
    .A2(_04600_),
    .B1(_04602_),
    .B2(\rbzero.spi_registers.texadd2[17] ),
    .X(_04678_));
 sky130_fd_sc_hd__a211o_1 _11486_ (.A1(\rbzero.spi_registers.texadd1[17] ),
    .A2(_04597_),
    .B1(_04605_),
    .C1(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__o21a_1 _11487_ (.A1(\rbzero.spi_registers.texadd0[17] ),
    .A2(_04594_),
    .B1(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__a22o_1 _11488_ (.A1(\rbzero.spi_registers.texadd3[18] ),
    .A2(_04600_),
    .B1(_04602_),
    .B2(\rbzero.spi_registers.texadd2[18] ),
    .X(_04681_));
 sky130_fd_sc_hd__a211o_1 _11489_ (.A1(\rbzero.spi_registers.texadd1[18] ),
    .A2(_04597_),
    .B1(_04606_),
    .C1(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__o21a_1 _11490_ (.A1(\rbzero.spi_registers.texadd0[18] ),
    .A2(_04595_),
    .B1(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__and3_1 _11491_ (.A(_04677_),
    .B(_04680_),
    .C(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(\rbzero.spi_registers.texadd3[19] ),
    .A2(_04600_),
    .B1(_04603_),
    .B2(\rbzero.spi_registers.texadd2[19] ),
    .X(_04685_));
 sky130_fd_sc_hd__a211o_1 _11493_ (.A1(\rbzero.spi_registers.texadd1[19] ),
    .A2(_04597_),
    .B1(_04606_),
    .C1(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__o21a_1 _11494_ (.A1(\rbzero.spi_registers.texadd0[19] ),
    .A2(_04595_),
    .B1(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__and2_1 _11495_ (.A(_04684_),
    .B(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__a22o_1 _11496_ (.A1(\rbzero.spi_registers.texadd3[20] ),
    .A2(_04600_),
    .B1(_04603_),
    .B2(\rbzero.spi_registers.texadd2[20] ),
    .X(_04689_));
 sky130_fd_sc_hd__a211o_1 _11497_ (.A1(\rbzero.spi_registers.texadd1[20] ),
    .A2(_04598_),
    .B1(_04606_),
    .C1(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__o21a_1 _11498_ (.A1(\rbzero.spi_registers.texadd0[20] ),
    .A2(_04595_),
    .B1(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__nand2_1 _11499_ (.A(_04688_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__a22o_1 _11500_ (.A1(\rbzero.spi_registers.texadd3[21] ),
    .A2(_04600_),
    .B1(_04603_),
    .B2(\rbzero.spi_registers.texadd2[21] ),
    .X(_04693_));
 sky130_fd_sc_hd__a211o_1 _11501_ (.A1(\rbzero.spi_registers.texadd1[21] ),
    .A2(_04598_),
    .B1(_04606_),
    .C1(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__o21a_1 _11502_ (.A1(\rbzero.spi_registers.texadd0[21] ),
    .A2(_04595_),
    .B1(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__or2b_1 _11503_ (.A(_04692_),
    .B_N(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__mux2_1 _11504_ (.A0(_04611_),
    .A1(_04612_),
    .S(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__o31a_1 _11505_ (.A1(_04105_),
    .A2(_04608_),
    .A3(_04697_),
    .B1(_04583_),
    .X(_04698_));
 sky130_fd_sc_hd__o21ai_1 _11506_ (.A1(_04105_),
    .A2(_04608_),
    .B1(_04697_),
    .Y(_04699_));
 sky130_fd_sc_hd__clkinv_4 _11507_ (.A(\gpout0.hpos[0] ),
    .Y(_04700_));
 sky130_fd_sc_hd__a31o_1 _11508_ (.A1(_04684_),
    .A2(_04687_),
    .A3(_04691_),
    .B1(_04695_),
    .X(_04701_));
 sky130_fd_sc_hd__a31o_1 _11509_ (.A1(_04700_),
    .A2(_04696_),
    .A3(_04701_),
    .B1(_04583_),
    .X(_04702_));
 sky130_fd_sc_hd__or2_1 _11510_ (.A(_04688_),
    .B(_04691_),
    .X(_04703_));
 sky130_fd_sc_hd__and3_1 _11511_ (.A(_04105_),
    .B(_04692_),
    .C(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__o2bb2a_1 _11512_ (.A1_N(_04698_),
    .A2_N(_04699_),
    .B1(_04702_),
    .B2(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__and2_1 _11513_ (.A(_04677_),
    .B(_04680_),
    .X(_04706_));
 sky130_fd_sc_hd__nor3_1 _11514_ (.A(_04700_),
    .B(_04706_),
    .C(_04683_),
    .Y(_04707_));
 sky130_fd_sc_hd__o22a_1 _11515_ (.A1(_04105_),
    .A2(_04687_),
    .B1(_04707_),
    .B2(_04684_),
    .X(_04708_));
 sky130_fd_sc_hd__o31ai_1 _11516_ (.A1(_04105_),
    .A2(_04684_),
    .A3(_04687_),
    .B1(_04583_),
    .Y(_04709_));
 sky130_fd_sc_hd__nor2_1 _11517_ (.A(_04708_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__buf_4 _11518_ (.A(\gpout0.hpos[1] ),
    .X(_04711_));
 sky130_fd_sc_hd__and3_1 _11519_ (.A(_04104_),
    .B(_04673_),
    .C(_04676_),
    .X(_04712_));
 sky130_fd_sc_hd__o22ai_1 _11520_ (.A1(_04105_),
    .A2(_04680_),
    .B1(_04712_),
    .B2(_04677_),
    .Y(_04713_));
 sky130_fd_sc_hd__or3_1 _11521_ (.A(_04104_),
    .B(_04677_),
    .C(_04680_),
    .X(_04714_));
 sky130_fd_sc_hd__a31o_1 _11522_ (.A1(_04711_),
    .A2(_04713_),
    .A3(_04714_),
    .B1(_04579_),
    .X(_04715_));
 sky130_fd_sc_hd__o221a_1 _11523_ (.A1(_04589_),
    .A2(_04705_),
    .B1(_04710_),
    .B2(_04715_),
    .C1(_04554_),
    .X(_04716_));
 sky130_fd_sc_hd__a22o_1 _11524_ (.A1(\rbzero.spi_registers.texadd2[5] ),
    .A2(_04603_),
    .B1(_04613_),
    .B2(\rbzero.spi_registers.texadd3[5] ),
    .X(_04717_));
 sky130_fd_sc_hd__a221o_1 _11525_ (.A1(\rbzero.spi_registers.texadd1[5] ),
    .A2(_04598_),
    .B1(_04606_),
    .B2(\rbzero.spi_registers.texadd0[5] ),
    .C1(_04104_),
    .X(_04718_));
 sky130_fd_sc_hd__a31o_1 _11526_ (.A1(\rbzero.spi_registers.texadd0[4] ),
    .A2(_04600_),
    .A3(_04592_),
    .B1(_04700_),
    .X(_04719_));
 sky130_fd_sc_hd__a22o_1 _11527_ (.A1(\rbzero.spi_registers.texadd2[4] ),
    .A2(_04603_),
    .B1(_04613_),
    .B2(\rbzero.spi_registers.texadd3[4] ),
    .X(_04720_));
 sky130_fd_sc_hd__a211o_1 _11528_ (.A1(\rbzero.spi_registers.texadd1[4] ),
    .A2(_04598_),
    .B1(_04719_),
    .C1(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__o21ai_1 _11529_ (.A1(_04717_),
    .A2(_04718_),
    .B1(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__and2_1 _11530_ (.A(_04645_),
    .B(_04646_),
    .X(_04723_));
 sky130_fd_sc_hd__a21oi_1 _11531_ (.A1(_04643_),
    .A2(_04644_),
    .B1(\rbzero.texu_hot[0] ),
    .Y(_04724_));
 sky130_fd_sc_hd__or3b_1 _11532_ (.A(_04724_),
    .B(_04700_),
    .C_N(_04645_),
    .X(_04725_));
 sky130_fd_sc_hd__o311a_1 _11533_ (.A1(_04104_),
    .A2(_04647_),
    .A3(_04723_),
    .B1(_04725_),
    .C1(_04583_),
    .X(_04726_));
 sky130_fd_sc_hd__a211oi_1 _11534_ (.A1(_04711_),
    .A2(_04722_),
    .B1(_04726_),
    .C1(_04589_),
    .Y(_04727_));
 sky130_fd_sc_hd__a22o_1 _11535_ (.A1(\rbzero.spi_registers.texadd2[1] ),
    .A2(_04603_),
    .B1(_04613_),
    .B2(\rbzero.spi_registers.texadd3[1] ),
    .X(_04728_));
 sky130_fd_sc_hd__a21o_1 _11536_ (.A1(\rbzero.spi_registers.texadd1[1] ),
    .A2(_04598_),
    .B1(_04606_),
    .X(_04729_));
 sky130_fd_sc_hd__o221a_1 _11537_ (.A1(\rbzero.spi_registers.texadd0[1] ),
    .A2(_04595_),
    .B1(_04728_),
    .B2(_04729_),
    .C1(_04700_),
    .X(_04730_));
 sky130_fd_sc_hd__a22o_1 _11538_ (.A1(\rbzero.spi_registers.texadd2[0] ),
    .A2(_04603_),
    .B1(_04613_),
    .B2(\rbzero.spi_registers.texadd3[0] ),
    .X(_04731_));
 sky130_fd_sc_hd__a211o_1 _11539_ (.A1(\rbzero.spi_registers.texadd1[0] ),
    .A2(_04598_),
    .B1(_04606_),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__o211a_1 _11540_ (.A1(\rbzero.spi_registers.texadd0[0] ),
    .A2(_04595_),
    .B1(_04732_),
    .C1(_04104_),
    .X(_04733_));
 sky130_fd_sc_hd__a22o_1 _11541_ (.A1(\rbzero.spi_registers.texadd2[2] ),
    .A2(_04603_),
    .B1(_04613_),
    .B2(\rbzero.spi_registers.texadd3[2] ),
    .X(_04734_));
 sky130_fd_sc_hd__a211o_1 _11542_ (.A1(\rbzero.spi_registers.texadd1[2] ),
    .A2(_04598_),
    .B1(_04606_),
    .C1(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__o211a_1 _11543_ (.A1(\rbzero.spi_registers.texadd0[2] ),
    .A2(_04595_),
    .B1(_04735_),
    .C1(_04103_),
    .X(_04736_));
 sky130_fd_sc_hd__a22o_1 _11544_ (.A1(\rbzero.spi_registers.texadd3[3] ),
    .A2(_04613_),
    .B1(_04598_),
    .B2(\rbzero.spi_registers.texadd1[3] ),
    .X(_04737_));
 sky130_fd_sc_hd__o21a_1 _11545_ (.A1(\rbzero.spi_registers.texadd2[3] ),
    .A2(_04600_),
    .B1(_04592_),
    .X(_04738_));
 sky130_fd_sc_hd__o221a_1 _11546_ (.A1(\rbzero.spi_registers.texadd0[3] ),
    .A2(_04595_),
    .B1(_04737_),
    .B2(_04738_),
    .C1(_04700_),
    .X(_04739_));
 sky130_fd_sc_hd__or3_1 _11547_ (.A(_04711_),
    .B(_04736_),
    .C(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__o311a_1 _11548_ (.A1(_04583_),
    .A2(_04730_),
    .A3(_04733_),
    .B1(_04740_),
    .C1(_04589_),
    .X(_04741_));
 sky130_fd_sc_hd__nand3_1 _11549_ (.A(_04655_),
    .B(_04634_),
    .C(_04653_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand3_1 _11550_ (.A(_04658_),
    .B(_04630_),
    .C(_04656_),
    .Y(_04743_));
 sky130_fd_sc_hd__and3_1 _11551_ (.A(_04700_),
    .B(_04659_),
    .C(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__a311o_1 _11552_ (.A1(_04104_),
    .A2(_04656_),
    .A3(_04742_),
    .B1(_04744_),
    .C1(_04711_),
    .X(_04745_));
 sky130_fd_sc_hd__xnor2_1 _11553_ (.A(_04650_),
    .B(_04652_),
    .Y(_04746_));
 sky130_fd_sc_hd__or2_1 _11554_ (.A(_04649_),
    .B(_04638_),
    .X(_04747_));
 sky130_fd_sc_hd__xnor2_1 _11555_ (.A(_04747_),
    .B(_04648_),
    .Y(_04748_));
 sky130_fd_sc_hd__mux2_1 _11556_ (.A0(_04746_),
    .A1(_04748_),
    .S(_04104_),
    .X(_04749_));
 sky130_fd_sc_hd__nand2_1 _11557_ (.A(_04711_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__a311o_1 _11558_ (.A1(_04668_),
    .A2(_04666_),
    .A3(_04667_),
    .B1(_04615_),
    .C1(_04665_),
    .X(_04751_));
 sky130_fd_sc_hd__or3b_1 _11559_ (.A(_04711_),
    .B(_04669_),
    .C_N(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__nand2_1 _11560_ (.A(_04711_),
    .B(_04662_),
    .Y(_04753_));
 sky130_fd_sc_hd__a31o_1 _11561_ (.A1(_04661_),
    .A2(_04626_),
    .A3(_04659_),
    .B1(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__a31o_1 _11562_ (.A1(_04104_),
    .A2(_04752_),
    .A3(_04754_),
    .B1(_04589_),
    .X(_04755_));
 sky130_fd_sc_hd__or3_1 _11563_ (.A(_04614_),
    .B(_04669_),
    .C(_04672_),
    .X(_04756_));
 sky130_fd_sc_hd__o311a_1 _11564_ (.A1(_04615_),
    .A2(_04663_),
    .A3(_04664_),
    .B1(_04622_),
    .C1(_04662_),
    .X(_04757_));
 sky130_fd_sc_hd__o31ai_1 _11565_ (.A1(_04583_),
    .A2(_04665_),
    .A3(_04757_),
    .B1(_04700_),
    .Y(_04758_));
 sky130_fd_sc_hd__a31o_1 _11566_ (.A1(_04583_),
    .A2(_04756_),
    .A3(_04673_),
    .B1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__and2b_1 _11567_ (.A_N(_04755_),
    .B(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__a311o_1 _11568_ (.A1(_04589_),
    .A2(_04745_),
    .A3(_04750_),
    .B1(_04588_),
    .C1(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__xnor2_2 _11569_ (.A(_04546_),
    .B(_04557_),
    .Y(_04762_));
 sky130_fd_sc_hd__o311a_1 _11570_ (.A1(_04586_),
    .A2(_04727_),
    .A3(_04741_),
    .B1(_04761_),
    .C1(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__nor2_1 _11571_ (.A(_04586_),
    .B(_04587_),
    .Y(_04764_));
 sky130_fd_sc_hd__o211a_1 _11572_ (.A1(_04763_),
    .A2(_04764_),
    .B1(_04556_),
    .C1(_04560_),
    .X(_04765_));
 sky130_fd_sc_hd__o31a_1 _11573_ (.A1(_04586_),
    .A2(_04588_),
    .A3(_04716_),
    .B1(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__a31o_4 _11574_ (.A1(_04550_),
    .A2(_04560_),
    .A3(_04585_),
    .B1(_04766_),
    .X(net73));
 sky130_fd_sc_hd__buf_1 _11575_ (.A(clknet_leaf_35_i_clk),
    .X(_04767_));
 sky130_fd_sc_hd__inv_2 _20835__4 (.A(clknet_1_1__leaf__03704_),
    .Y(net129));
 sky130_fd_sc_hd__clkinv_2 _11577_ (.A(net2),
    .Y(_04768_));
 sky130_fd_sc_hd__nor2_4 _11578_ (.A(_04579_),
    .B(_04580_),
    .Y(_04769_));
 sky130_fd_sc_hd__and2_1 _11579_ (.A(\gpout0.hpos[3] ),
    .B(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__or2_1 _11580_ (.A(\gpout0.hpos[4] ),
    .B(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__o21a_1 _11581_ (.A1(_04547_),
    .A2(_04771_),
    .B1(\gpout0.hpos[6] ),
    .X(_04772_));
 sky130_fd_sc_hd__and2_1 _11582_ (.A(\gpout0.hpos[7] ),
    .B(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__a21oi_2 _11583_ (.A1(\gpout0.hpos[8] ),
    .A2(_04773_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04774_));
 sky130_fd_sc_hd__clkbuf_4 _11584_ (.A(\gpout0.vpos[7] ),
    .X(_04775_));
 sky130_fd_sc_hd__clkinv_4 _11585_ (.A(net3),
    .Y(_04776_));
 sky130_fd_sc_hd__or4_2 _11586_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.vpos[8] ),
    .C(_04775_),
    .D(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__buf_4 _11587_ (.A(\gpout0.vpos[5] ),
    .X(_04778_));
 sky130_fd_sc_hd__or2_1 _11588_ (.A(_04778_),
    .B(\gpout0.vpos[4] ),
    .X(_04779_));
 sky130_fd_sc_hd__or2_1 _11589_ (.A(\gpout0.vpos[3] ),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__or3_2 _11590_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(\gpout0.vpos[0] ),
    .X(_04781_));
 sky130_fd_sc_hd__clkbuf_4 _11591_ (.A(\gpout0.vpos[6] ),
    .X(_04782_));
 sky130_fd_sc_hd__o21a_1 _11592_ (.A1(_04780_),
    .A2(_04781_),
    .B1(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__nor3_4 _11593_ (.A(_04774_),
    .B(_04777_),
    .C(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__or2_1 _11594_ (.A(\gpout0.vpos[4] ),
    .B(\gpout0.vpos[3] ),
    .X(_04785_));
 sky130_fd_sc_hd__nand2_1 _11595_ (.A(\gpout0.vpos[4] ),
    .B(\gpout0.vpos[3] ),
    .Y(_04786_));
 sky130_fd_sc_hd__clkbuf_4 _11596_ (.A(_04778_),
    .X(_04787_));
 sky130_fd_sc_hd__buf_4 _11597_ (.A(\gpout0.vpos[4] ),
    .X(_04788_));
 sky130_fd_sc_hd__nand2_1 _11598_ (.A(_04787_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__o21ai_1 _11599_ (.A1(_04579_),
    .A2(_04580_),
    .B1(_04781_),
    .Y(_04790_));
 sky130_fd_sc_hd__a41o_1 _11600_ (.A1(_04779_),
    .A2(_04785_),
    .A3(_04786_),
    .A4(_04789_),
    .B1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__and2_1 _11601_ (.A(_04784_),
    .B(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__clkbuf_4 _11602_ (.A(\gpout0.vpos[3] ),
    .X(_04793_));
 sky130_fd_sc_hd__nand2_1 _11603_ (.A(_04793_),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .Y(_04794_));
 sky130_fd_sc_hd__or2_1 _11604_ (.A(\gpout0.vpos[3] ),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .X(_04795_));
 sky130_fd_sc_hd__xor2_1 _11605_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_04106_),
    .X(_04796_));
 sky130_fd_sc_hd__a221o_1 _11606_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_04548_),
    .B1(_04546_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .C1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__xor2_1 _11607_ (.A(_04778_),
    .B(\rbzero.debug_overlay.playerY[2] ),
    .X(_04798_));
 sky130_fd_sc_hd__a211o_1 _11608_ (.A1(_04794_),
    .A2(_04795_),
    .B1(_04797_),
    .C1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__inv_2 _11609_ (.A(\gpout0.vpos[7] ),
    .Y(_04800_));
 sky130_fd_sc_hd__inv_2 _11610_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .Y(_04801_));
 sky130_fd_sc_hd__clkinv_2 _11611_ (.A(\gpout0.vpos[6] ),
    .Y(_04802_));
 sky130_fd_sc_hd__inv_2 _11612_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .Y(_04803_));
 sky130_fd_sc_hd__clkinv_2 _11613_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .Y(_04804_));
 sky130_fd_sc_hd__o22a_1 _11614_ (.A1(\gpout0.vpos[7] ),
    .A2(_04803_),
    .B1(_04804_),
    .B2(_04547_),
    .X(_04805_));
 sky130_fd_sc_hd__o221a_1 _11615_ (.A1(_04802_),
    .A2(\rbzero.debug_overlay.playerY[3] ),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .B2(_04555_),
    .C1(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__o221a_1 _11616_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_04546_),
    .B1(_04587_),
    .B2(_04801_),
    .C1(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__o221a_1 _11617_ (.A1(_04800_),
    .A2(\rbzero.debug_overlay.playerY[4] ),
    .B1(\rbzero.debug_overlay.playerX[1] ),
    .B2(_04549_),
    .C1(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__inv_2 _11618_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .Y(_04809_));
 sky130_fd_sc_hd__xnor2_1 _11619_ (.A(\gpout0.vpos[4] ),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .Y(_04810_));
 sky130_fd_sc_hd__o221a_1 _11620_ (.A1(\gpout0.vpos[6] ),
    .A2(_04809_),
    .B1(\rbzero.debug_overlay.playerX[0] ),
    .B2(_04548_),
    .C1(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__and3b_1 _11621_ (.A_N(_04799_),
    .B(_04808_),
    .C(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__or2_1 _11622_ (.A(\gpout0.hpos[2] ),
    .B(_04581_),
    .X(_04813_));
 sky130_fd_sc_hd__nand2_1 _11623_ (.A(_04813_),
    .B(_04781_),
    .Y(_04814_));
 sky130_fd_sc_hd__or2_1 _11624_ (.A(_04812_),
    .B(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__inv_2 _11625_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .Y(_04816_));
 sky130_fd_sc_hd__clkinv_4 _11626_ (.A(_04778_),
    .Y(_04817_));
 sky130_fd_sc_hd__xnor2_1 _11627_ (.A(_04788_),
    .B(\rbzero.map_overlay.i_mapdy[1] ),
    .Y(_04818_));
 sky130_fd_sc_hd__o221a_1 _11628_ (.A1(_04782_),
    .A2(_04816_),
    .B1(\rbzero.map_overlay.i_mapdy[2] ),
    .B2(_04817_),
    .C1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__inv_2 _11629_ (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .Y(_04820_));
 sky130_fd_sc_hd__o2bb2a_1 _11630_ (.A1_N(\rbzero.map_overlay.i_mapdy[2] ),
    .A2_N(_04817_),
    .B1(_04775_),
    .B2(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__clkinv_4 _11631_ (.A(\gpout0.vpos[3] ),
    .Y(_04822_));
 sky130_fd_sc_hd__or4_1 _11632_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_overlay.i_mapdy[2] ),
    .C(\rbzero.map_overlay.i_mapdy[1] ),
    .D(\rbzero.map_overlay.i_mapdy[0] ),
    .X(_04823_));
 sky130_fd_sc_hd__o21a_1 _11633_ (.A1(\rbzero.map_overlay.i_mapdy[5] ),
    .A2(_04823_),
    .B1(_04800_),
    .X(_04824_));
 sky130_fd_sc_hd__o2bb2a_1 _11634_ (.A1_N(_04822_),
    .A2_N(\rbzero.map_overlay.i_mapdy[0] ),
    .B1(\rbzero.map_overlay.i_mapdy[3] ),
    .B2(_04802_),
    .X(_04825_));
 sky130_fd_sc_hd__o221a_1 _11635_ (.A1(_04822_),
    .A2(\rbzero.map_overlay.i_mapdy[0] ),
    .B1(_04824_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__and3_1 _11636_ (.A(_04819_),
    .B(_04821_),
    .C(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__a22o_1 _11637_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04548_),
    .B1(_04549_),
    .B2(\rbzero.map_overlay.i_mapdx[1] ),
    .X(_04828_));
 sky130_fd_sc_hd__o22a_1 _11638_ (.A1(\rbzero.map_overlay.i_mapdx[4] ),
    .A2(_04186_),
    .B1(_04549_),
    .B2(\rbzero.map_overlay.i_mapdx[1] ),
    .X(_04829_));
 sky130_fd_sc_hd__or4_1 _11639_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(\rbzero.map_overlay.i_mapdx[2] ),
    .C(\rbzero.map_overlay.i_mapdx[1] ),
    .D(\rbzero.map_overlay.i_mapdx[0] ),
    .X(_04830_));
 sky130_fd_sc_hd__inv_2 _11640_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .Y(_04831_));
 sky130_fd_sc_hd__o21a_1 _11641_ (.A1(\rbzero.map_overlay.i_mapdx[5] ),
    .A2(_04830_),
    .B1(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__xnor2_1 _11642_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_04553_),
    .Y(_04833_));
 sky130_fd_sc_hd__o221a_1 _11643_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04548_),
    .B1(_04106_),
    .B2(_04832_),
    .C1(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__buf_4 _11644_ (.A(_04547_),
    .X(_04835_));
 sky130_fd_sc_hd__xnor2_1 _11645_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__and4b_1 _11646_ (.A_N(_04828_),
    .B(_04829_),
    .C(_04834_),
    .D(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__inv_2 _11647_ (.A(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__inv_2 _11648_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .Y(_04839_));
 sky130_fd_sc_hd__xnor2_1 _11649_ (.A(\gpout0.vpos[4] ),
    .B(\rbzero.map_overlay.i_othery[1] ),
    .Y(_04840_));
 sky130_fd_sc_hd__o221a_1 _11650_ (.A1(_04839_),
    .A2(_04554_),
    .B1(_04555_),
    .B2(\rbzero.map_overlay.i_otherx[2] ),
    .C1(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__inv_2 _11651_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .Y(_04842_));
 sky130_fd_sc_hd__xnor2_1 _11652_ (.A(_04778_),
    .B(\rbzero.map_overlay.i_othery[2] ),
    .Y(_04843_));
 sky130_fd_sc_hd__o221a_1 _11653_ (.A1(_04800_),
    .A2(\rbzero.map_overlay.i_othery[4] ),
    .B1(_04842_),
    .B2(_04587_),
    .C1(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__nand2_1 _11654_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_04106_),
    .Y(_04845_));
 sky130_fd_sc_hd__or2_1 _11655_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_04106_),
    .X(_04846_));
 sky130_fd_sc_hd__xor2_1 _11656_ (.A(_04793_),
    .B(\rbzero.map_overlay.i_othery[0] ),
    .X(_04847_));
 sky130_fd_sc_hd__xor2_1 _11657_ (.A(\gpout0.vpos[6] ),
    .B(\rbzero.map_overlay.i_othery[3] ),
    .X(_04848_));
 sky130_fd_sc_hd__a221o_1 _11658_ (.A1(_04800_),
    .A2(\rbzero.map_overlay.i_othery[4] ),
    .B1(_04842_),
    .B2(_04587_),
    .C1(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__xor2_1 _11659_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(\gpout0.hpos[3] ),
    .X(_04850_));
 sky130_fd_sc_hd__a221o_1 _11660_ (.A1(_04839_),
    .A2(_04553_),
    .B1(_04555_),
    .B2(\rbzero.map_overlay.i_otherx[2] ),
    .C1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__a2111oi_1 _11661_ (.A1(_04845_),
    .A2(_04846_),
    .B1(_04847_),
    .C1(_04849_),
    .D1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__and3_1 _11662_ (.A(_04841_),
    .B(_04844_),
    .C(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__a21oi_1 _11663_ (.A1(_04827_),
    .A2(_04838_),
    .B1(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__xnor2_1 _11664_ (.A(\gpout0.vpos[1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .Y(_04855_));
 sky130_fd_sc_hd__inv_2 _11665_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .Y(_04856_));
 sky130_fd_sc_hd__o22a_1 _11666_ (.A1(\gpout0.vpos[0] ),
    .A2(_04856_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .B2(_04579_),
    .X(_04857_));
 sky130_fd_sc_hd__and3_1 _11667_ (.A(_04812_),
    .B(_04855_),
    .C(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__inv_2 _11668_ (.A(\gpout0.vpos[0] ),
    .Y(_04859_));
 sky130_fd_sc_hd__xnor2_1 _11669_ (.A(\gpout0.vpos[2] ),
    .B(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_04860_));
 sky130_fd_sc_hd__o221a_1 _11670_ (.A1(_04859_),
    .A2(\rbzero.debug_overlay.playerY[-3] ),
    .B1(\rbzero.debug_overlay.playerX[-2] ),
    .B2(_04583_),
    .C1(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__inv_2 _11671_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_04862_));
 sky130_fd_sc_hd__inv_2 _11672_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .Y(_04863_));
 sky130_fd_sc_hd__xnor2_1 _11673_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_04103_),
    .Y(_04864_));
 sky130_fd_sc_hd__o221a_1 _11674_ (.A1(_04862_),
    .A2(\gpout0.hpos[2] ),
    .B1(\gpout0.hpos[1] ),
    .B2(_04863_),
    .C1(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__or3_1 _11675_ (.A(\gpout0.vpos[7] ),
    .B(\gpout0.vpos[6] ),
    .C(_04779_),
    .X(_04866_));
 sky130_fd_sc_hd__o31a_1 _11676_ (.A1(_04793_),
    .A2(_04781_),
    .A3(_04866_),
    .B1(\gpout0.vpos[8] ),
    .X(_04867_));
 sky130_fd_sc_hd__or3b_1 _11677_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.hpos[9] ),
    .C_N(net1),
    .X(_04868_));
 sky130_fd_sc_hd__or2_1 _11678_ (.A(\gpout0.hpos[6] ),
    .B(\gpout0.hpos[5] ),
    .X(_04869_));
 sky130_fd_sc_hd__or3_1 _11679_ (.A(\gpout0.hpos[3] ),
    .B(_04587_),
    .C(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__o31a_1 _11680_ (.A1(_04107_),
    .A2(_04813_),
    .A3(_04870_),
    .B1(_04109_),
    .X(_04871_));
 sky130_fd_sc_hd__or3_1 _11681_ (.A(_04867_),
    .B(_04868_),
    .C(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__a31o_1 _11682_ (.A1(_04858_),
    .A2(_04861_),
    .A3(_04865_),
    .B1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__o21ba_1 _11683_ (.A1(_04815_),
    .A2(_04854_),
    .B1_N(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _11684_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_04875_));
 sky130_fd_sc_hd__or2_1 _11685_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .X(_04876_));
 sky130_fd_sc_hd__nand2_1 _11686_ (.A(_04875_),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__or2_1 _11687_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _11688_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .Y(_04879_));
 sky130_fd_sc_hd__a21boi_1 _11689_ (.A1(\rbzero.texV[8] ),
    .A2(_04878_),
    .B1_N(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _11690_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .Y(_04881_));
 sky130_fd_sc_hd__or2_1 _11691_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .X(_04882_));
 sky130_fd_sc_hd__nand3_1 _11692_ (.A(\rbzero.texV[7] ),
    .B(_04881_),
    .C(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__a21o_1 _11693_ (.A1(_04881_),
    .A2(_04882_),
    .B1(\rbzero.texV[7] ),
    .X(_04884_));
 sky130_fd_sc_hd__nand2_1 _11694_ (.A(_04883_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_1 _11695_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .Y(_04886_));
 sky130_fd_sc_hd__or2_1 _11696_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .X(_04887_));
 sky130_fd_sc_hd__nand3_1 _11697_ (.A(\rbzero.texV[6] ),
    .B(_04886_),
    .C(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__nand3_1 _11698_ (.A(_04885_),
    .B(_04886_),
    .C(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__a21o_1 _11699_ (.A1(_04886_),
    .A2(_04887_),
    .B1(\rbzero.texV[6] ),
    .X(_04890_));
 sky130_fd_sc_hd__nand2_1 _11700_ (.A(_04888_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__and2_1 _11701_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .X(_04892_));
 sky130_fd_sc_hd__nor2_1 _11702_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .Y(_04893_));
 sky130_fd_sc_hd__nor2_1 _11703_ (.A(_04892_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__a21oi_1 _11704_ (.A1(\rbzero.texV[5] ),
    .A2(_04894_),
    .B1(_04892_),
    .Y(_04895_));
 sky130_fd_sc_hd__xnor2_1 _11705_ (.A(_04891_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__nand2_1 _11706_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .Y(_04897_));
 sky130_fd_sc_hd__or2_1 _11707_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .X(_04898_));
 sky130_fd_sc_hd__nand3_1 _11708_ (.A(\rbzero.texV[4] ),
    .B(_04897_),
    .C(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__xnor2_1 _11709_ (.A(\rbzero.texV[5] ),
    .B(_04894_),
    .Y(_04900_));
 sky130_fd_sc_hd__a21oi_1 _11710_ (.A1(_04897_),
    .A2(_04899_),
    .B1(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__a21o_1 _11711_ (.A1(_04897_),
    .A2(_04898_),
    .B1(\rbzero.texV[4] ),
    .X(_04902_));
 sky130_fd_sc_hd__nand2_1 _11712_ (.A(_04899_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__or2_1 _11713_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_1 _11714_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .Y(_04905_));
 sky130_fd_sc_hd__a21boi_1 _11715_ (.A1(\rbzero.texV[3] ),
    .A2(_04904_),
    .B1_N(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__nor2_1 _11716_ (.A(_04903_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__xnor2_1 _11717_ (.A(_04903_),
    .B(_04906_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand2_1 _11718_ (.A(_04905_),
    .B(_04904_),
    .Y(_04909_));
 sky130_fd_sc_hd__xor2_1 _11719_ (.A(\rbzero.texV[3] ),
    .B(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__o211a_1 _11720_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(\rbzero.texV[1] ),
    .B1(\rbzero.texV[0] ),
    .C1(\rbzero.traced_texVinit[0] ),
    .X(_04911_));
 sky130_fd_sc_hd__a221o_1 _11721_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(\rbzero.texV[1] ),
    .B2(\rbzero.traced_texVinit[1] ),
    .C1(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__o21ai_4 _11722_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__or2_1 _11723_ (.A(_04910_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__buf_4 _11724_ (.A(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__nor2_2 _11725_ (.A(_04908_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__and3_1 _11726_ (.A(_04900_),
    .B(_04897_),
    .C(_04899_),
    .X(_04917_));
 sky130_fd_sc_hd__or2_1 _11727_ (.A(_04901_),
    .B(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__inv_2 _11728_ (.A(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__o21a_1 _11729_ (.A1(_04907_),
    .A2(_04916_),
    .B1(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__nor2_1 _11730_ (.A(_04901_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__nor2_1 _11731_ (.A(_04896_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21bai_2 _11732_ (.A1(_04891_),
    .A2(_04895_),
    .B1_N(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__a21oi_1 _11733_ (.A1(_04886_),
    .A2(_04888_),
    .B1(_04885_),
    .Y(_04924_));
 sky130_fd_sc_hd__a21o_1 _11734_ (.A1(_04889_),
    .A2(_04923_),
    .B1(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__nand2_1 _11735_ (.A(_04879_),
    .B(_04878_),
    .Y(_04926_));
 sky130_fd_sc_hd__xor2_1 _11736_ (.A(\rbzero.texV[8] ),
    .B(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__nand3_1 _11737_ (.A(_04881_),
    .B(_04883_),
    .C(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _11738_ (.A(_04925_),
    .B(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__a21o_1 _11739_ (.A1(_04881_),
    .A2(_04883_),
    .B1(_04927_),
    .X(_04930_));
 sky130_fd_sc_hd__o21a_1 _11740_ (.A1(_04877_),
    .A2(_04880_),
    .B1(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__a22oi_2 _11741_ (.A1(_04877_),
    .A2(_04880_),
    .B1(_04929_),
    .B2(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__xor2_1 _11742_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .X(_04933_));
 sky130_fd_sc_hd__xnor2_1 _11743_ (.A(_04875_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__a21oi_1 _11744_ (.A1(_04932_),
    .A2(_04934_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04935_));
 sky130_fd_sc_hd__o21a_4 _11745_ (.A1(_04932_),
    .A2(_04934_),
    .B1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__inv_2 _11746_ (.A(_04889_),
    .Y(_04937_));
 sky130_fd_sc_hd__nor2_1 _11747_ (.A(_04937_),
    .B(_04924_),
    .Y(_04938_));
 sky130_fd_sc_hd__xnor2_2 _11748_ (.A(_04923_),
    .B(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__or2_4 _11749_ (.A(_04936_),
    .B(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__buf_6 _11750_ (.A(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__and3_1 _11751_ (.A(_04925_),
    .B(_04930_),
    .C(_04928_),
    .X(_04942_));
 sky130_fd_sc_hd__a21o_1 _11752_ (.A1(_04930_),
    .A2(_04928_),
    .B1(_04925_),
    .X(_04943_));
 sky130_fd_sc_hd__or3b_1 _11753_ (.A(_04936_),
    .B(_04942_),
    .C_N(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__buf_6 _11754_ (.A(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__and2_1 _11755_ (.A(_04896_),
    .B(_04921_),
    .X(_04946_));
 sky130_fd_sc_hd__or3_2 _11756_ (.A(_04922_),
    .B(_04936_),
    .C(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__buf_4 _11757_ (.A(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__nor3_2 _11758_ (.A(_04919_),
    .B(_04907_),
    .C(_04916_),
    .Y(_04949_));
 sky130_fd_sc_hd__or3_4 _11759_ (.A(_04920_),
    .B(_04936_),
    .C(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__buf_6 _11760_ (.A(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__nand2_1 _11761_ (.A(_04908_),
    .B(_04915_),
    .Y(_04952_));
 sky130_fd_sc_hd__or3b_1 _11762_ (.A(_04916_),
    .B(_04936_),
    .C_N(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__buf_4 _11763_ (.A(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__buf_4 _11764_ (.A(_04950_),
    .X(_04955_));
 sky130_fd_sc_hd__a21oi_4 _11765_ (.A1(_04910_),
    .A2(_04913_),
    .B1(_04936_),
    .Y(_04956_));
 sky130_fd_sc_hd__nand2_4 _11766_ (.A(_04915_),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__buf_6 _11767_ (.A(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__o211a_1 _11768_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_04954_),
    .B1(_04958_),
    .C1(\rbzero.floor_leak[0] ),
    .X(_04959_));
 sky130_fd_sc_hd__a221o_1 _11769_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_04954_),
    .B1(_04955_),
    .B2(\rbzero.floor_leak[2] ),
    .C1(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__o221a_1 _11770_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_04951_),
    .B1(_04947_),
    .B2(\rbzero.floor_leak[3] ),
    .C1(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__a221o_1 _11771_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04948_),
    .B1(_04940_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__o221a_1 _11772_ (.A1(\rbzero.floor_leak[4] ),
    .A2(_04941_),
    .B1(_04945_),
    .B2(\rbzero.floor_leak[5] ),
    .C1(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__nor3_4 _11773_ (.A(_04922_),
    .B(_04936_),
    .C(_04946_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand2_1 _11774_ (.A(_04954_),
    .B(_04950_),
    .Y(_04965_));
 sky130_fd_sc_hd__buf_4 _11775_ (.A(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__and2_2 _11776_ (.A(_04915_),
    .B(_04956_),
    .X(_04967_));
 sky130_fd_sc_hd__nand2_1 _11777_ (.A(_04940_),
    .B(_04945_),
    .Y(_04968_));
 sky130_fd_sc_hd__or2_1 _11778_ (.A(_04106_),
    .B(_04553_),
    .X(_04969_));
 sky130_fd_sc_hd__a21oi_4 _11779_ (.A1(_04109_),
    .A2(_04969_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04970_));
 sky130_fd_sc_hd__or3_1 _11780_ (.A(_04967_),
    .B(_04968_),
    .C(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__or3_1 _11781_ (.A(\rbzero.row_render.size[2] ),
    .B(\rbzero.row_render.size[1] ),
    .C(\rbzero.row_render.size[0] ),
    .X(_04972_));
 sky130_fd_sc_hd__or2_1 _11782_ (.A(\rbzero.row_render.size[3] ),
    .B(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__or3_1 _11783_ (.A(\rbzero.row_render.size[5] ),
    .B(\rbzero.row_render.size[4] ),
    .C(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__and2_1 _11784_ (.A(\rbzero.row_render.size[6] ),
    .B(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__or2_1 _11785_ (.A(\rbzero.row_render.size[7] ),
    .B(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__xor2_1 _11786_ (.A(\rbzero.row_render.size[8] ),
    .B(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__a21oi_1 _11787_ (.A1(\rbzero.row_render.size[8] ),
    .A2(_04976_),
    .B1(\rbzero.row_render.size[9] ),
    .Y(_04978_));
 sky130_fd_sc_hd__and3_1 _11788_ (.A(\rbzero.row_render.size[9] ),
    .B(\rbzero.row_render.size[8] ),
    .C(_04976_),
    .X(_04979_));
 sky130_fd_sc_hd__nand2_1 _11789_ (.A(\rbzero.row_render.size[7] ),
    .B(_04975_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2_1 _11790_ (.A(_04976_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__nor2_1 _11791_ (.A(\rbzero.row_render.size[6] ),
    .B(_04974_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_1 _11792_ (.A(_04975_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__o21ai_1 _11793_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_04973_),
    .B1(\rbzero.row_render.size[5] ),
    .Y(_04984_));
 sky130_fd_sc_hd__nand2_1 _11794_ (.A(_04974_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__xnor2_1 _11795_ (.A(\rbzero.row_render.size[4] ),
    .B(_04973_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_1 _11796_ (.A(\rbzero.row_render.size[3] ),
    .B(_04972_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand2_1 _11797_ (.A(_04973_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__o21ai_1 _11798_ (.A1(\rbzero.row_render.size[1] ),
    .A2(\rbzero.row_render.size[0] ),
    .B1(\rbzero.row_render.size[2] ),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_1 _11799_ (.A(_04972_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__o211a_1 _11800_ (.A1(\rbzero.row_render.size[0] ),
    .A2(\gpout0.hpos[1] ),
    .B1(_04581_),
    .C1(\rbzero.row_render.size[1] ),
    .X(_04991_));
 sky130_fd_sc_hd__nor2_1 _11801_ (.A(\rbzero.row_render.size[1] ),
    .B(\rbzero.row_render.size[0] ),
    .Y(_04992_));
 sky130_fd_sc_hd__a221o_1 _11802_ (.A1(\rbzero.row_render.size[2] ),
    .A2(\gpout0.hpos[2] ),
    .B1(\gpout0.hpos[1] ),
    .B2(_04103_),
    .C1(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__o22a_1 _11803_ (.A1(\gpout0.hpos[2] ),
    .A2(_04990_),
    .B1(_04991_),
    .B2(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__o21a_1 _11804_ (.A1(\gpout0.hpos[3] ),
    .A2(_04988_),
    .B1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__a221o_1 _11805_ (.A1(\gpout0.hpos[3] ),
    .A2(_04988_),
    .B1(_04986_),
    .B2(\gpout0.hpos[4] ),
    .C1(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__o221a_1 _11806_ (.A1(\gpout0.hpos[4] ),
    .A2(_04986_),
    .B1(_04985_),
    .B2(_04547_),
    .C1(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__a221o_1 _11807_ (.A1(_04547_),
    .A2(_04985_),
    .B1(_04983_),
    .B2(_04553_),
    .C1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__o221a_1 _11808_ (.A1(_04553_),
    .A2(_04983_),
    .B1(_04981_),
    .B2(\gpout0.hpos[7] ),
    .C1(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__a221o_1 _11809_ (.A1(\gpout0.hpos[7] ),
    .A2(_04981_),
    .B1(_04977_),
    .B2(_04109_),
    .C1(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__o221a_1 _11810_ (.A1(_04109_),
    .A2(_04977_),
    .B1(_04978_),
    .B2(_04979_),
    .C1(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__a21o_1 _11811_ (.A1(\rbzero.row_render.size[7] ),
    .A2(\rbzero.row_render.size[6] ),
    .B1(\rbzero.row_render.size[8] ),
    .X(_05002_));
 sky130_fd_sc_hd__nor2_1 _11812_ (.A(\rbzero.row_render.size[9] ),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__xnor2_1 _11813_ (.A(\rbzero.row_render.size[7] ),
    .B(\rbzero.row_render.size[6] ),
    .Y(_05004_));
 sky130_fd_sc_hd__nand3_1 _11814_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(\rbzero.row_render.size[6] ),
    .Y(_05005_));
 sky130_fd_sc_hd__and2_1 _11815_ (.A(_05002_),
    .B(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__a21o_1 _11816_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_04582_),
    .B1(_04700_),
    .X(_05007_));
 sky130_fd_sc_hd__o22a_1 _11817_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_04579_),
    .B1(_04582_),
    .B2(\rbzero.row_render.size[1] ),
    .X(_05008_));
 sky130_fd_sc_hd__o21a_1 _11818_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_05007_),
    .B1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__a221o_1 _11819_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_04548_),
    .B1(_04579_),
    .B2(\rbzero.row_render.size[2] ),
    .C1(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__o221a_1 _11820_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_04548_),
    .B1(_04549_),
    .B2(\rbzero.row_render.size[4] ),
    .C1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__a221o_1 _11821_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_04555_),
    .B1(_04549_),
    .B2(\rbzero.row_render.size[4] ),
    .C1(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__o2bb2a_1 _11822_ (.A1_N(\rbzero.row_render.size[6] ),
    .A2_N(\gpout0.hpos[6] ),
    .B1(_04555_),
    .B2(\rbzero.row_render.size[5] ),
    .X(_05013_));
 sky130_fd_sc_hd__nand2_1 _11823_ (.A(_05012_),
    .B(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__o221a_1 _11824_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_04553_),
    .B1(_05004_),
    .B2(\gpout0.hpos[7] ),
    .C1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__a221o_1 _11825_ (.A1(\gpout0.hpos[7] ),
    .A2(_05004_),
    .B1(_05006_),
    .B2(_04109_),
    .C1(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__o2bb2a_1 _11826_ (.A1_N(\rbzero.row_render.size[9] ),
    .A2_N(_05002_),
    .B1(_05006_),
    .B2(_04109_),
    .X(_05017_));
 sky130_fd_sc_hd__a22o_1 _11827_ (.A1(\gpout0.hpos[9] ),
    .A2(_05003_),
    .B1(_05016_),
    .B2(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__o21ai_1 _11828_ (.A1(\gpout0.hpos[9] ),
    .A2(_05003_),
    .B1(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__o21a_1 _11829_ (.A1(\gpout0.hpos[9] ),
    .A2(_05001_),
    .B1(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__or3b_4 _11830_ (.A(\rbzero.row_render.size[10] ),
    .B(_05020_),
    .C_N(_04978_),
    .X(_05021_));
 sky130_fd_sc_hd__o31a_1 _11831_ (.A1(_04964_),
    .A2(_04966_),
    .A3(_04971_),
    .B1(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__a2bb2o_1 _11832_ (.A1_N(\rbzero.row_render.vinf ),
    .A2_N(_05022_),
    .B1(_04945_),
    .B2(\rbzero.floor_leak[5] ),
    .X(_05023_));
 sky130_fd_sc_hd__nor2_1 _11833_ (.A(_04963_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__clkbuf_4 _11834_ (.A(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__mux2_1 _11835_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_04970_),
    .X(_05026_));
 sky130_fd_sc_hd__or2_1 _11836_ (.A(_05025_),
    .B(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__clkinv_2 _11837_ (.A(net42),
    .Y(_05028_));
 sky130_fd_sc_hd__nor2_4 _11838_ (.A(_04936_),
    .B(_04939_),
    .Y(_05029_));
 sky130_fd_sc_hd__buf_6 _11839_ (.A(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__nor3_4 _11840_ (.A(_04920_),
    .B(_04936_),
    .C(_04949_),
    .Y(_05031_));
 sky130_fd_sc_hd__buf_6 _11841_ (.A(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__buf_6 _11842_ (.A(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__buf_8 _11843_ (.A(_04958_),
    .X(_05034_));
 sky130_fd_sc_hd__buf_6 _11844_ (.A(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__mux2_1 _11845_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_05035_),
    .X(_05037_));
 sky130_fd_sc_hd__nor3b_4 _11847_ (.A(_04916_),
    .B(_04936_),
    .C_N(_04952_),
    .Y(_05038_));
 sky130_fd_sc_hd__buf_4 _11848_ (.A(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__buf_4 _11849_ (.A(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__clkbuf_8 _11850_ (.A(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__mux2_1 _11851_ (.A0(_05036_),
    .A1(_05037_),
    .S(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__buf_6 _11852_ (.A(_05038_),
    .X(_05043_));
 sky130_fd_sc_hd__buf_6 _11853_ (.A(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__buf_6 _11854_ (.A(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__buf_8 _11855_ (.A(_04957_),
    .X(_05046_));
 sky130_fd_sc_hd__buf_6 _11856_ (.A(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__buf_6 _11857_ (.A(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__buf_4 _11859_ (.A(_04915_),
    .X(_05050_));
 sky130_fd_sc_hd__buf_4 _11860_ (.A(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__buf_4 _11861_ (.A(_04956_),
    .X(_05052_));
 sky130_fd_sc_hd__buf_4 _11862_ (.A(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__and3_1 _11863_ (.A(\rbzero.tex_r0[51] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__buf_6 _11864_ (.A(_04957_),
    .X(_05055_));
 sky130_fd_sc_hd__buf_6 _11865_ (.A(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__buf_6 _11866_ (.A(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__buf_6 _11867_ (.A(_04954_),
    .X(_05058_));
 sky130_fd_sc_hd__buf_4 _11868_ (.A(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__a21o_1 _11869_ (.A1(\rbzero.tex_r0[50] ),
    .A2(_05057_),
    .B1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__buf_6 _11870_ (.A(_04951_),
    .X(_05061_));
 sky130_fd_sc_hd__buf_6 _11871_ (.A(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__o221a_1 _11872_ (.A1(_05045_),
    .A2(_05049_),
    .B1(_05054_),
    .B2(_05060_),
    .C1(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__buf_6 _11873_ (.A(_04964_),
    .X(_05064_));
 sky130_fd_sc_hd__a211o_1 _11874_ (.A1(_05033_),
    .A2(_05042_),
    .B1(_05063_),
    .C1(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_05035_),
    .X(_05066_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_05035_),
    .X(_05067_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(_05066_),
    .A1(_05067_),
    .S(_05041_),
    .X(_05068_));
 sky130_fd_sc_hd__buf_6 _11878_ (.A(_04958_),
    .X(_05069_));
 sky130_fd_sc_hd__buf_6 _11879_ (.A(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__mux2_1 _11881_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_05034_),
    .X(_05072_));
 sky130_fd_sc_hd__or2_1 _11882_ (.A(_05059_),
    .B(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__o211a_1 _11883_ (.A1(_05045_),
    .A2(_05071_),
    .B1(_05073_),
    .C1(_05033_),
    .X(_05074_));
 sky130_fd_sc_hd__buf_6 _11884_ (.A(_04948_),
    .X(_05075_));
 sky130_fd_sc_hd__a211o_1 _11885_ (.A1(_05062_),
    .A2(_05068_),
    .B1(_05074_),
    .C1(_05075_),
    .X(_05076_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_05048_),
    .X(_05077_));
 sky130_fd_sc_hd__buf_6 _11887_ (.A(_05046_),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__or2_1 _11889_ (.A(_05044_),
    .B(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__buf_6 _11890_ (.A(_05031_),
    .X(_05081_));
 sky130_fd_sc_hd__o211a_1 _11891_ (.A1(_05059_),
    .A2(_05077_),
    .B1(_05080_),
    .C1(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_1 _11892_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_05048_),
    .X(_05083_));
 sky130_fd_sc_hd__and3_1 _11893_ (.A(\rbzero.tex_r0[43] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05084_));
 sky130_fd_sc_hd__buf_6 _11894_ (.A(_05069_),
    .X(_05085_));
 sky130_fd_sc_hd__a21o_1 _11895_ (.A1(\rbzero.tex_r0[42] ),
    .A2(_05085_),
    .B1(_05059_),
    .X(_05086_));
 sky130_fd_sc_hd__buf_4 _11896_ (.A(_04951_),
    .X(_05087_));
 sky130_fd_sc_hd__o221a_1 _11897_ (.A1(_05045_),
    .A2(_05083_),
    .B1(_05084_),
    .B2(_05086_),
    .C1(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__buf_6 _11898_ (.A(_04958_),
    .X(_05089_));
 sky130_fd_sc_hd__mux2_1 _11899_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_05089_),
    .X(_05091_));
 sky130_fd_sc_hd__mux2_1 _11901_ (.A0(_05090_),
    .A1(_05091_),
    .S(_05044_),
    .X(_05092_));
 sky130_fd_sc_hd__buf_6 _11902_ (.A(_05043_),
    .X(_05093_));
 sky130_fd_sc_hd__mux2_1 _11903_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_05069_),
    .X(_05094_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04958_),
    .X(_05095_));
 sky130_fd_sc_hd__or2_1 _11905_ (.A(_05058_),
    .B(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__o211a_1 _11906_ (.A1(_05093_),
    .A2(_05094_),
    .B1(_05096_),
    .C1(_05032_),
    .X(_05097_));
 sky130_fd_sc_hd__a211o_1 _11907_ (.A1(_05062_),
    .A2(_05092_),
    .B1(_05097_),
    .C1(_05064_),
    .X(_05098_));
 sky130_fd_sc_hd__o311a_1 _11908_ (.A1(_05075_),
    .A2(_05082_),
    .A3(_05088_),
    .B1(_04941_),
    .C1(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__a31o_1 _11909_ (.A1(_05030_),
    .A2(_05065_),
    .A3(_05076_),
    .B1(_05099_),
    .X(_05100_));
 sky130_fd_sc_hd__and2_1 _11910_ (.A(\rbzero.tex_r0[22] ),
    .B(_05048_),
    .X(_05101_));
 sky130_fd_sc_hd__a31o_1 _11911_ (.A1(\rbzero.tex_r0[23] ),
    .A2(_05050_),
    .A3(_05052_),
    .B1(_05058_),
    .X(_05102_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_05056_),
    .X(_05103_));
 sky130_fd_sc_hd__o221a_1 _11913_ (.A1(_05101_),
    .A2(_05102_),
    .B1(_05103_),
    .B2(_05041_),
    .C1(_05081_),
    .X(_05104_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_05056_),
    .X(_05105_));
 sky130_fd_sc_hd__and3_1 _11915_ (.A(\rbzero.tex_r0[19] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05106_));
 sky130_fd_sc_hd__buf_6 _11916_ (.A(_04954_),
    .X(_05107_));
 sky130_fd_sc_hd__clkbuf_8 _11917_ (.A(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__a21o_1 _11918_ (.A1(\rbzero.tex_r0[18] ),
    .A2(_05070_),
    .B1(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__o221a_1 _11919_ (.A1(_05041_),
    .A2(_05105_),
    .B1(_05106_),
    .B2(_05109_),
    .C1(_05061_),
    .X(_05110_));
 sky130_fd_sc_hd__mux2_1 _11920_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_05048_),
    .X(_05111_));
 sky130_fd_sc_hd__and3_1 _11921_ (.A(\rbzero.tex_r0[27] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05112_));
 sky130_fd_sc_hd__a21o_1 _11922_ (.A1(\rbzero.tex_r0[26] ),
    .A2(_05057_),
    .B1(_05059_),
    .X(_05113_));
 sky130_fd_sc_hd__o221a_1 _11923_ (.A1(_05045_),
    .A2(_05111_),
    .B1(_05112_),
    .B2(_05113_),
    .C1(_05062_),
    .X(_05114_));
 sky130_fd_sc_hd__mux2_1 _11924_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_05034_),
    .X(_05115_));
 sky130_fd_sc_hd__mux2_1 _11925_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_05034_),
    .X(_05116_));
 sky130_fd_sc_hd__mux2_1 _11926_ (.A0(_05115_),
    .A1(_05116_),
    .S(_05108_),
    .X(_05117_));
 sky130_fd_sc_hd__buf_6 _11927_ (.A(_04948_),
    .X(_05118_));
 sky130_fd_sc_hd__a21o_1 _11928_ (.A1(_05033_),
    .A2(_05117_),
    .B1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__o32a_1 _11929_ (.A1(_05064_),
    .A2(_05104_),
    .A3(_05110_),
    .B1(_05114_),
    .B2(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__mux2_1 _11930_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_05070_),
    .X(_05121_));
 sky130_fd_sc_hd__a31o_1 _11931_ (.A1(_05045_),
    .A2(_05087_),
    .A3(_05121_),
    .B1(_05118_),
    .X(_05122_));
 sky130_fd_sc_hd__nor2_2 _11932_ (.A(_05093_),
    .B(_05032_),
    .Y(_05123_));
 sky130_fd_sc_hd__or2_1 _11933_ (.A(\rbzero.tex_r0[8] ),
    .B(_04967_),
    .X(_05124_));
 sky130_fd_sc_hd__or2_1 _11934_ (.A(\rbzero.tex_r0[9] ),
    .B(_05085_),
    .X(_05125_));
 sky130_fd_sc_hd__mux2_1 _11935_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_05047_),
    .X(_05126_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_05047_),
    .X(_05127_));
 sky130_fd_sc_hd__mux2_1 _11937_ (.A0(_05126_),
    .A1(_05127_),
    .S(_05040_),
    .X(_05128_));
 sky130_fd_sc_hd__a32o_1 _11938_ (.A1(_05123_),
    .A2(_05124_),
    .A3(_05125_),
    .B1(_05128_),
    .B2(_05081_),
    .X(_05129_));
 sky130_fd_sc_hd__mux2_1 _11939_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_05047_),
    .X(_05130_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_05047_),
    .X(_05131_));
 sky130_fd_sc_hd__mux2_1 _11941_ (.A0(_05130_),
    .A1(_05131_),
    .S(_05040_),
    .X(_05132_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_05034_),
    .X(_05133_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_05046_),
    .X(_05134_));
 sky130_fd_sc_hd__or2_1 _11944_ (.A(_05043_),
    .B(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__o211a_1 _11945_ (.A1(_05059_),
    .A2(_05133_),
    .B1(_05135_),
    .C1(_05032_),
    .X(_05136_));
 sky130_fd_sc_hd__buf_6 _11946_ (.A(_04964_),
    .X(_05137_));
 sky130_fd_sc_hd__a211o_1 _11947_ (.A1(_05062_),
    .A2(_05132_),
    .B1(_05136_),
    .C1(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__o21a_1 _11948_ (.A1(_05122_),
    .A2(_05129_),
    .B1(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(_05120_),
    .A1(_05139_),
    .S(_04941_),
    .X(_05140_));
 sky130_fd_sc_hd__mux2_1 _11950_ (.A0(_05100_),
    .A1(_05140_),
    .S(_04945_),
    .X(_05141_));
 sky130_fd_sc_hd__inv_2 _11951_ (.A(\rbzero.row_render.side ),
    .Y(_05142_));
 sky130_fd_sc_hd__inv_2 _11952_ (.A(\rbzero.row_render.wall[0] ),
    .Y(_05143_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(_05143_),
    .B(\rbzero.row_render.wall[1] ),
    .Y(_05144_));
 sky130_fd_sc_hd__a21o_1 _11954_ (.A1(_05142_),
    .A2(_05144_),
    .B1(_05028_),
    .X(_05145_));
 sky130_fd_sc_hd__a31o_1 _11955_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_05057_),
    .A3(_05123_),
    .B1(_05142_),
    .X(_05146_));
 sky130_fd_sc_hd__nand2_1 _11956_ (.A(_05143_),
    .B(\rbzero.row_render.wall[1] ),
    .Y(_05147_));
 sky130_fd_sc_hd__buf_4 _11957_ (.A(_04966_),
    .X(_05148_));
 sky130_fd_sc_hd__or4bb_1 _11958_ (.A(\rbzero.row_render.texu[4] ),
    .B(\rbzero.row_render.texu[3] ),
    .C_N(\rbzero.row_render.texu[2] ),
    .D_N(\rbzero.row_render.texu[1] ),
    .X(_05149_));
 sky130_fd_sc_hd__nand2_1 _11959_ (.A(\rbzero.row_render.texu[4] ),
    .B(\rbzero.row_render.texu[3] ),
    .Y(_05150_));
 sky130_fd_sc_hd__o31a_1 _11960_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(\rbzero.row_render.texu[1] ),
    .A3(_05150_),
    .B1(_04964_),
    .X(_05151_));
 sky130_fd_sc_hd__a211o_1 _11961_ (.A1(_04948_),
    .A2(_05149_),
    .B1(_05151_),
    .C1(\rbzero.row_render.texu[0] ),
    .X(_05152_));
 sky130_fd_sc_hd__o31ai_2 _11962_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04967_),
    .A3(_05148_),
    .B1(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__nor2_1 _11963_ (.A(\rbzero.row_render.side ),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__nor2_1 _11964_ (.A(_05147_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__a32o_1 _11965_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(\rbzero.row_render.texu[2] ),
    .A3(\rbzero.row_render.texu[1] ),
    .B1(_05118_),
    .B2(_05123_),
    .X(_05156_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(\rbzero.row_render.wall[1] ),
    .B(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2_1 _11967_ (.A(_05038_),
    .B(_05031_),
    .Y(_05158_));
 sky130_fd_sc_hd__buf_4 _11968_ (.A(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__buf_4 _11969_ (.A(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__o32a_1 _11970_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(\rbzero.row_render.texu[2] ),
    .A3(\rbzero.row_render.texu[1] ),
    .B1(_04948_),
    .B2(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__nand2_1 _11971_ (.A(\rbzero.row_render.wall[0] ),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__or2_1 _11972_ (.A(\rbzero.row_render.side ),
    .B(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__o21ai_1 _11973_ (.A1(_05157_),
    .A2(_05162_),
    .B1(\rbzero.row_render.side ),
    .Y(_05164_));
 sky130_fd_sc_hd__o21ai_1 _11974_ (.A1(_05157_),
    .A2(_05163_),
    .B1(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__a221oi_1 _11975_ (.A1(_05146_),
    .A2(_05155_),
    .B1(_05165_),
    .B2(_05147_),
    .C1(_05144_),
    .Y(_05166_));
 sky130_fd_sc_hd__o21ai_1 _11976_ (.A1(_05145_),
    .A2(_05166_),
    .B1(_05025_),
    .Y(_05167_));
 sky130_fd_sc_hd__a21o_1 _11977_ (.A1(_05028_),
    .A2(_05141_),
    .B1(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__nor3_4 _11978_ (.A(_04867_),
    .B(_04868_),
    .C(_04871_),
    .Y(_05169_));
 sky130_fd_sc_hd__a21oi_1 _11979_ (.A1(_05027_),
    .A2(_05168_),
    .B1(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__inv_2 _11980_ (.A(_04784_),
    .Y(_05171_));
 sky130_fd_sc_hd__o21a_1 _11981_ (.A1(_04874_),
    .A2(_05170_),
    .B1(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__and3_2 _11982_ (.A(\rbzero.trace_state[3] ),
    .B(_04563_),
    .C(_04570_),
    .X(_05173_));
 sky130_fd_sc_hd__a21o_1 _11983_ (.A1(\rbzero.trace_state[0] ),
    .A2(_05173_),
    .B1(_04768_),
    .X(_05174_));
 sky130_fd_sc_hd__o21ai_1 _11984_ (.A1(_04792_),
    .A2(_05172_),
    .B1(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__o21ai_4 _11985_ (.A1(_04107_),
    .A2(_04109_),
    .B1(_04111_),
    .Y(_05176_));
 sky130_fd_sc_hd__clkbuf_4 _11986_ (.A(\gpout0.vpos[8] ),
    .X(_05177_));
 sky130_fd_sc_hd__and3_2 _11987_ (.A(\gpout0.vpos[7] ),
    .B(\gpout0.vpos[6] ),
    .C(_04778_),
    .X(_05178_));
 sky130_fd_sc_hd__a21oi_4 _11988_ (.A1(_05177_),
    .A2(_05178_),
    .B1(\gpout0.vpos[9] ),
    .Y(_05179_));
 sky130_fd_sc_hd__and2_2 _11989_ (.A(_05176_),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__o211a_4 _11990_ (.A1(\rbzero.trace_state[0] ),
    .A2(_04768_),
    .B1(_05175_),
    .C1(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__buf_4 _11991_ (.A(net45),
    .X(_05182_));
 sky130_fd_sc_hd__mux2_2 _11992_ (.A0(\reg_rgb[6] ),
    .A1(_05181_),
    .S(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__clkbuf_1 _11993_ (.A(_05183_),
    .X(net69));
 sky130_fd_sc_hd__nor2_1 _11994_ (.A(\gpout0.hpos[7] ),
    .B(_04772_),
    .Y(_05184_));
 sky130_fd_sc_hd__or2_1 _11995_ (.A(_04773_),
    .B(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__mux2_1 _11996_ (.A0(\gpout0.hpos[6] ),
    .A1(_04762_),
    .S(_04769_),
    .X(_05186_));
 sky130_fd_sc_hd__nor2_1 _11997_ (.A(\gpout0.hpos[3] ),
    .B(_04769_),
    .Y(_05187_));
 sky130_fd_sc_hd__or2_1 _11998_ (.A(_04770_),
    .B(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__nor2_1 _11999_ (.A(\gpout0.hpos[4] ),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__o21ba_1 _12000_ (.A1(_04771_),
    .A2(_04869_),
    .B1_N(_04772_),
    .X(_05190_));
 sky130_fd_sc_hd__or3_1 _12001_ (.A(_05186_),
    .B(_05189_),
    .C(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__or2_1 _12002_ (.A(_05185_),
    .B(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__a2bb2o_1 _12003_ (.A1_N(_05189_),
    .A2_N(_05190_),
    .B1(\gpout0.hpos[6] ),
    .B2(_04547_),
    .X(_05193_));
 sky130_fd_sc_hd__o21bai_1 _12004_ (.A1(_05185_),
    .A2(_05193_),
    .B1_N(_04773_),
    .Y(_05194_));
 sky130_fd_sc_hd__xnor2_1 _12005_ (.A(_04109_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__or2_1 _12006_ (.A(_05192_),
    .B(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__nand2_1 _12007_ (.A(_05192_),
    .B(_05195_),
    .Y(_05197_));
 sky130_fd_sc_hd__a21o_4 _12008_ (.A1(_05196_),
    .A2(_05197_),
    .B1(_05186_),
    .X(_05198_));
 sky130_fd_sc_hd__mux2_2 _12009_ (.A0(_04547_),
    .A1(_04558_),
    .S(_04769_),
    .X(_05199_));
 sky130_fd_sc_hd__o21a_4 _12010_ (.A1(\gpout0.hpos[7] ),
    .A2(\gpout0.hpos[8] ),
    .B1(\gpout0.hpos[9] ),
    .X(_05200_));
 sky130_fd_sc_hd__or3b_2 _12011_ (.A(_04774_),
    .B(_05200_),
    .C_N(_05192_),
    .X(_05201_));
 sky130_fd_sc_hd__nor2_1 _12012_ (.A(_05188_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__and2_1 _12013_ (.A(\gpout0.hpos[4] ),
    .B(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__nand2_1 _12014_ (.A(_05199_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__nor2_4 _12015_ (.A(_05198_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__or2b_1 _12016_ (.A(_05201_),
    .B_N(_05188_),
    .X(_05206_));
 sky130_fd_sc_hd__a21bo_1 _12017_ (.A1(_04550_),
    .A2(_04769_),
    .B1_N(_04771_),
    .X(_05207_));
 sky130_fd_sc_hd__and2b_1 _12018_ (.A_N(_05206_),
    .B(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__nand2_2 _12019_ (.A(_05199_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__nor2_4 _12020_ (.A(_05198_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__or2_1 _12021_ (.A(_04551_),
    .B(_04557_),
    .X(_05211_));
 sky130_fd_sc_hd__mux2_2 _12022_ (.A0(_04555_),
    .A1(_05211_),
    .S(_04769_),
    .X(_05212_));
 sky130_fd_sc_hd__or2_1 _12023_ (.A(_05207_),
    .B(_05206_),
    .X(_05213_));
 sky130_fd_sc_hd__or2_1 _12024_ (.A(_05212_),
    .B(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__nor2_4 _12025_ (.A(_05198_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__a22o_1 _12026_ (.A1(\rbzero.debug_overlay.vplaneY[0] ),
    .A2(_05210_),
    .B1(_05215_),
    .B2(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_05216_));
 sky130_fd_sc_hd__nand2_2 _12027_ (.A(_05212_),
    .B(_05203_),
    .Y(_05217_));
 sky130_fd_sc_hd__nand2_1 _12028_ (.A(_04549_),
    .B(_05202_),
    .Y(_05218_));
 sky130_fd_sc_hd__or2_2 _12029_ (.A(_05212_),
    .B(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__nand2_2 _12030_ (.A(_05186_),
    .B(_05195_),
    .Y(_05220_));
 sky130_fd_sc_hd__a41o_1 _12031_ (.A1(_05209_),
    .A2(_05213_),
    .A3(_05217_),
    .A4(_05219_),
    .B1(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__nand2_1 _12032_ (.A(_05191_),
    .B(_05193_),
    .Y(_05222_));
 sky130_fd_sc_hd__xnor2_1 _12033_ (.A(_05185_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__a31o_1 _12034_ (.A1(_05221_),
    .A2(_05204_),
    .A3(_05214_),
    .B1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__o31ai_4 _12035_ (.A1(_05198_),
    .A2(_05199_),
    .A3(_05201_),
    .B1(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__clkbuf_4 _12036_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_05226_));
 sky130_fd_sc_hd__or2_1 _12037_ (.A(_05199_),
    .B(_05218_),
    .X(_05227_));
 sky130_fd_sc_hd__nor2_2 _12038_ (.A(_05220_),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__nand2_1 _12039_ (.A(_05212_),
    .B(_05208_),
    .Y(_05229_));
 sky130_fd_sc_hd__nor2_2 _12040_ (.A(_05220_),
    .B(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__a221o_1 _12041_ (.A1(_05226_),
    .A2(_05228_),
    .B1(_05230_),
    .B2(\rbzero.debug_overlay.vplaneY[-4] ),
    .C1(_04822_),
    .X(_05231_));
 sky130_fd_sc_hd__nor2_4 _12042_ (.A(_05198_),
    .B(_05219_),
    .Y(_05232_));
 sky130_fd_sc_hd__or2_1 _12043_ (.A(_04547_),
    .B(_05213_),
    .X(_05233_));
 sky130_fd_sc_hd__or2b_4 _12044_ (.A(_05220_),
    .B_N(_05223_),
    .X(_05234_));
 sky130_fd_sc_hd__nor2_4 _12045_ (.A(_05233_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__nor2_4 _12046_ (.A(_05219_),
    .B(_05234_),
    .Y(_05236_));
 sky130_fd_sc_hd__a22o_1 _12047_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(_05235_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_05237_));
 sky130_fd_sc_hd__nor2_4 _12048_ (.A(_05217_),
    .B(_05234_),
    .Y(_05238_));
 sky130_fd_sc_hd__nor2_4 _12049_ (.A(_05209_),
    .B(_05234_),
    .Y(_05239_));
 sky130_fd_sc_hd__a22o_1 _12050_ (.A1(\rbzero.debug_overlay.vplaneY[-7] ),
    .A2(_05238_),
    .B1(_05239_),
    .B2(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_05240_));
 sky130_fd_sc_hd__a211o_1 _12051_ (.A1(\rbzero.debug_overlay.vplaneY[-1] ),
    .A2(_05232_),
    .B1(_05237_),
    .C1(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__a211o_1 _12052_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(_05225_),
    .B1(_05231_),
    .C1(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__a211o_1 _12053_ (.A1(\rbzero.debug_overlay.vplaneY[-3] ),
    .A2(_05205_),
    .B1(_05216_),
    .C1(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__a22o_1 _12054_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_05210_),
    .B1(_05215_),
    .B2(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_05244_));
 sky130_fd_sc_hd__a21o_1 _12055_ (.A1(\rbzero.debug_overlay.vplaneX[-3] ),
    .A2(_05205_),
    .B1(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__buf_2 _12056_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_05246_));
 sky130_fd_sc_hd__a22o_1 _12057_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(_05235_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_05247_));
 sky130_fd_sc_hd__a221o_1 _12058_ (.A1(\rbzero.debug_overlay.vplaneX[-7] ),
    .A2(_05238_),
    .B1(_05239_),
    .B2(_05246_),
    .C1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__clkbuf_4 _12059_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_05249_));
 sky130_fd_sc_hd__a221o_1 _12060_ (.A1(_05249_),
    .A2(_05228_),
    .B1(_05230_),
    .B2(\rbzero.debug_overlay.vplaneX[-4] ),
    .C1(\gpout0.vpos[3] ),
    .X(_05250_));
 sky130_fd_sc_hd__a211o_1 _12061_ (.A1(\rbzero.debug_overlay.vplaneX[-1] ),
    .A2(_05232_),
    .B1(_05248_),
    .C1(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__a211o_1 _12062_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_05225_),
    .B1(_05245_),
    .C1(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__and3b_1 _12063_ (.A_N(_04789_),
    .B(_05243_),
    .C(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__a22o_1 _12064_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_05235_),
    .B1(_05238_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .X(_05254_));
 sky130_fd_sc_hd__a22o_1 _12065_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_05228_),
    .B1(_05230_),
    .B2(\rbzero.debug_overlay.facingY[-4] ),
    .X(_05255_));
 sky130_fd_sc_hd__a221o_1 _12066_ (.A1(\rbzero.debug_overlay.facingY[-1] ),
    .A2(_05232_),
    .B1(_05239_),
    .B2(\rbzero.debug_overlay.facingY[-8] ),
    .C1(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__a22o_1 _12067_ (.A1(\rbzero.debug_overlay.facingY[-3] ),
    .A2(_05205_),
    .B1(_05215_),
    .B2(\rbzero.debug_overlay.facingY[-2] ),
    .X(_05257_));
 sky130_fd_sc_hd__a221o_1 _12068_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_05225_),
    .B1(_05210_),
    .B2(\rbzero.debug_overlay.facingY[0] ),
    .C1(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__or2_1 _12069_ (.A(_05256_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__a211o_1 _12070_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(_05236_),
    .B1(_05254_),
    .C1(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__nor2_2 _12071_ (.A(_04817_),
    .B(\gpout0.vpos[4] ),
    .Y(_05261_));
 sky130_fd_sc_hd__and3_1 _12072_ (.A(_04822_),
    .B(_05260_),
    .C(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__nor2_1 _12073_ (.A(_04778_),
    .B(_04786_),
    .Y(_05263_));
 sky130_fd_sc_hd__a22o_1 _12074_ (.A1(\rbzero.debug_overlay.facingX[-6] ),
    .A2(_05235_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.facingX[-9] ),
    .X(_05264_));
 sky130_fd_sc_hd__a22o_1 _12075_ (.A1(\rbzero.debug_overlay.facingX[-7] ),
    .A2(_05238_),
    .B1(_05239_),
    .B2(\rbzero.debug_overlay.facingX[-8] ),
    .X(_05265_));
 sky130_fd_sc_hd__a21bo_1 _12076_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_05230_),
    .B1_N(_05263_),
    .X(_05266_));
 sky130_fd_sc_hd__a221o_1 _12077_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(_05215_),
    .B1(_05228_),
    .B2(\rbzero.debug_overlay.facingX[-5] ),
    .C1(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__or3_1 _12078_ (.A(_05264_),
    .B(_05265_),
    .C(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__a22o_1 _12079_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(_05232_),
    .B1(_05205_),
    .B2(\rbzero.debug_overlay.facingX[-3] ),
    .X(_05269_));
 sky130_fd_sc_hd__a221o_1 _12080_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_05225_),
    .B1(_05210_),
    .B2(\rbzero.debug_overlay.facingX[0] ),
    .C1(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__o32a_1 _12081_ (.A1(_05253_),
    .A2(_05262_),
    .A3(_05263_),
    .B1(_05268_),
    .B2(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__o21ba_1 _12082_ (.A1(_04787_),
    .A2(_04788_),
    .B1_N(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__nor2_1 _12083_ (.A(_05198_),
    .B(_05227_),
    .Y(_05273_));
 sky130_fd_sc_hd__a22o_1 _12084_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_05232_),
    .B1(_05215_),
    .B2(\rbzero.debug_overlay.playerX[-2] ),
    .X(_05274_));
 sky130_fd_sc_hd__a221o_1 _12085_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_05273_),
    .B1(_05210_),
    .B2(\rbzero.debug_overlay.playerX[0] ),
    .C1(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__nor2_1 _12086_ (.A(_05198_),
    .B(_05217_),
    .Y(_05276_));
 sky130_fd_sc_hd__nor2_1 _12087_ (.A(_05198_),
    .B(_05233_),
    .Y(_05277_));
 sky130_fd_sc_hd__nor2_1 _12088_ (.A(_05198_),
    .B(_05229_),
    .Y(_05278_));
 sky130_fd_sc_hd__nor2_1 _12089_ (.A(_05223_),
    .B(_05204_),
    .Y(_05279_));
 sky130_fd_sc_hd__a221o_1 _12090_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_05230_),
    .B1(_05279_),
    .B2(\rbzero.debug_overlay.playerX[5] ),
    .C1(_04780_),
    .X(_05280_));
 sky130_fd_sc_hd__a221o_1 _12091_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_05278_),
    .B1(_05228_),
    .B2(\rbzero.debug_overlay.playerX[-5] ),
    .C1(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__a221o_1 _12092_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_05277_),
    .B1(_05205_),
    .B2(\rbzero.debug_overlay.playerX[-3] ),
    .C1(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__a22o_1 _12093_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_05235_),
    .B1(_05238_),
    .B2(\rbzero.debug_overlay.playerX[-7] ),
    .X(_05283_));
 sky130_fd_sc_hd__a221o_1 _12094_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(_05236_),
    .B1(_05239_),
    .B2(\rbzero.debug_overlay.playerX[-8] ),
    .C1(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__a211o_1 _12095_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_05276_),
    .B1(_05282_),
    .C1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__nor2_1 _12096_ (.A(_05275_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__a22o_1 _12097_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_05232_),
    .B1(_05205_),
    .B2(\rbzero.debug_overlay.playerY[-3] ),
    .X(_05287_));
 sky130_fd_sc_hd__a221o_1 _12098_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_05273_),
    .B1(_05210_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .C1(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__a22o_1 _12099_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_05230_),
    .B1(_05279_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .X(_05289_));
 sky130_fd_sc_hd__or3_1 _12100_ (.A(_04822_),
    .B(_04779_),
    .C(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__a221o_1 _12101_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_05278_),
    .B1(_05228_),
    .B2(\rbzero.debug_overlay.playerY[-5] ),
    .C1(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__a221o_1 _12102_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_05277_),
    .B1(_05215_),
    .B2(\rbzero.debug_overlay.playerY[-2] ),
    .C1(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__a22o_1 _12103_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_05235_),
    .B1(_05239_),
    .B2(\rbzero.debug_overlay.playerY[-8] ),
    .X(_05293_));
 sky130_fd_sc_hd__a221o_1 _12104_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_05238_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .C1(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__a211o_1 _12105_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_05276_),
    .B1(_05292_),
    .C1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__nor2_1 _12106_ (.A(_05288_),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__or4_1 _12107_ (.A(_04790_),
    .B(_05272_),
    .C(_05286_),
    .D(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__or4b_1 _12108_ (.A(_04586_),
    .B(_04588_),
    .C(_04969_),
    .D_N(_04769_),
    .X(_05298_));
 sky130_fd_sc_hd__or3_1 _12109_ (.A(_04188_),
    .B(_05211_),
    .C(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__and3_2 _12110_ (.A(_04784_),
    .B(_05297_),
    .C(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_1 _12111_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_05048_),
    .X(_05301_));
 sky130_fd_sc_hd__buf_6 _12112_ (.A(_04957_),
    .X(_05302_));
 sky130_fd_sc_hd__buf_6 _12113_ (.A(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__mux2_1 _12114_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__buf_8 _12115_ (.A(_05302_),
    .X(_05305_));
 sky130_fd_sc_hd__mux2_1 _12116_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__nand2_4 _12117_ (.A(_05038_),
    .B(_04950_),
    .Y(_05307_));
 sky130_fd_sc_hd__mux2_1 _12118_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_05302_),
    .X(_05308_));
 sky130_fd_sc_hd__or3_1 _12119_ (.A(_05039_),
    .B(_04955_),
    .C(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__o221a_1 _12120_ (.A1(_05159_),
    .A2(_05304_),
    .B1(_05306_),
    .B2(_05307_),
    .C1(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__o211a_1 _12121_ (.A1(_04966_),
    .A2(_05301_),
    .B1(_05310_),
    .C1(_05118_),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _12122_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_05035_),
    .X(_05312_));
 sky130_fd_sc_hd__mux2_1 _12123_ (.A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_05305_),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_05078_),
    .X(_05314_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_05302_),
    .X(_05315_));
 sky130_fd_sc_hd__or3_1 _12126_ (.A(_05039_),
    .B(_04955_),
    .C(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__o221a_1 _12127_ (.A1(_05159_),
    .A2(_05313_),
    .B1(_05314_),
    .B2(_05307_),
    .C1(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__o211a_1 _12128_ (.A1(_05148_),
    .A2(_05312_),
    .B1(_05317_),
    .C1(_05137_),
    .X(_05318_));
 sky130_fd_sc_hd__mux2_1 _12129_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_05085_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _12130_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_05089_),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _12131_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_05089_),
    .X(_05321_));
 sky130_fd_sc_hd__buf_4 _12132_ (.A(_05307_),
    .X(_05322_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_05046_),
    .X(_05323_));
 sky130_fd_sc_hd__or3_1 _12134_ (.A(_05043_),
    .B(_04955_),
    .C(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__o221a_1 _12135_ (.A1(_05159_),
    .A2(_05320_),
    .B1(_05321_),
    .B2(_05322_),
    .C1(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__o211a_1 _12136_ (.A1(_05148_),
    .A2(_05319_),
    .B1(_05325_),
    .C1(_05075_),
    .X(_05326_));
 sky130_fd_sc_hd__mux2_1 _12137_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(_05069_),
    .X(_05327_));
 sky130_fd_sc_hd__or2_1 _12138_ (.A(_04966_),
    .B(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_05034_),
    .X(_05329_));
 sky130_fd_sc_hd__mux2_1 _12140_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_05089_),
    .X(_05330_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_05046_),
    .X(_05331_));
 sky130_fd_sc_hd__or3_1 _12142_ (.A(_05043_),
    .B(_04955_),
    .C(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__o221a_1 _12143_ (.A1(_05159_),
    .A2(_05329_),
    .B1(_05330_),
    .B2(_05322_),
    .C1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__a31o_1 _12144_ (.A1(_05137_),
    .A2(_05328_),
    .A3(_05333_),
    .B1(_05029_),
    .X(_05334_));
 sky130_fd_sc_hd__o32a_1 _12145_ (.A1(_04941_),
    .A2(_05311_),
    .A3(_05318_),
    .B1(_05326_),
    .B2(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__mux2_1 _12146_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_05047_),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _12147_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_05078_),
    .X(_05337_));
 sky130_fd_sc_hd__mux2_1 _12148_ (.A0(_05336_),
    .A1(_05337_),
    .S(_05040_),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _12149_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_05078_),
    .X(_05339_));
 sky130_fd_sc_hd__a31o_1 _12150_ (.A1(\rbzero.tex_r1[23] ),
    .A2(_05050_),
    .A3(_05052_),
    .B1(_05107_),
    .X(_05340_));
 sky130_fd_sc_hd__and2_1 _12151_ (.A(\rbzero.tex_r1[22] ),
    .B(_05069_),
    .X(_05341_));
 sky130_fd_sc_hd__o221a_1 _12152_ (.A1(_05044_),
    .A2(_05339_),
    .B1(_05340_),
    .B2(_05341_),
    .C1(_05032_),
    .X(_05342_));
 sky130_fd_sc_hd__a211o_1 _12153_ (.A1(_05087_),
    .A2(_05338_),
    .B1(_05342_),
    .C1(_05137_),
    .X(_05343_));
 sky130_fd_sc_hd__mux2_1 _12154_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_05078_),
    .X(_05344_));
 sky130_fd_sc_hd__or2_1 _12155_ (.A(_05108_),
    .B(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__buf_6 _12156_ (.A(_05046_),
    .X(_05346_));
 sky130_fd_sc_hd__mux2_1 _12157_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__o21a_1 _12158_ (.A1(_05044_),
    .A2(_05347_),
    .B1(_05032_),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _12159_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_05305_),
    .X(_05349_));
 sky130_fd_sc_hd__mux2_1 _12160_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_05305_),
    .X(_05350_));
 sky130_fd_sc_hd__buf_6 _12161_ (.A(_05039_),
    .X(_05351_));
 sky130_fd_sc_hd__mux2_1 _12162_ (.A0(_05349_),
    .A1(_05350_),
    .S(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__a221o_1 _12163_ (.A1(_05345_),
    .A2(_05348_),
    .B1(_05352_),
    .B2(_05087_),
    .C1(_05118_),
    .X(_05353_));
 sky130_fd_sc_hd__mux2_1 _12164_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_05303_),
    .X(_05354_));
 sky130_fd_sc_hd__and2_1 _12165_ (.A(\rbzero.tex_r1[4] ),
    .B(_05069_),
    .X(_05355_));
 sky130_fd_sc_hd__a31o_1 _12166_ (.A1(\rbzero.tex_r1[5] ),
    .A2(_05050_),
    .A3(_05052_),
    .B1(_05043_),
    .X(_05356_));
 sky130_fd_sc_hd__o221a_1 _12167_ (.A1(_05108_),
    .A2(_05354_),
    .B1(_05355_),
    .B2(_05356_),
    .C1(_05031_),
    .X(_05357_));
 sky130_fd_sc_hd__mux2_1 _12168_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[0] ),
    .S(_05305_),
    .X(_05358_));
 sky130_fd_sc_hd__and3_1 _12169_ (.A(\rbzero.tex_r1[3] ),
    .B(_05050_),
    .C(_05052_),
    .X(_05359_));
 sky130_fd_sc_hd__a21o_1 _12170_ (.A1(\rbzero.tex_r1[2] ),
    .A2(_05069_),
    .B1(_05107_),
    .X(_05360_));
 sky130_fd_sc_hd__o221a_1 _12171_ (.A1(_05044_),
    .A2(_05358_),
    .B1(_05359_),
    .B2(_05360_),
    .C1(_05061_),
    .X(_05361_));
 sky130_fd_sc_hd__mux2_1 _12172_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04958_),
    .X(_05362_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_04958_),
    .X(_05363_));
 sky130_fd_sc_hd__mux2_1 _12174_ (.A0(_05362_),
    .A1(_05363_),
    .S(_05043_),
    .X(_05364_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_04958_),
    .X(_05365_));
 sky130_fd_sc_hd__a21o_1 _12176_ (.A1(\rbzero.tex_r1[14] ),
    .A2(_05055_),
    .B1(_04954_),
    .X(_05366_));
 sky130_fd_sc_hd__and3_1 _12177_ (.A(\rbzero.tex_r1[15] ),
    .B(_04915_),
    .C(_04956_),
    .X(_05367_));
 sky130_fd_sc_hd__o221a_1 _12178_ (.A1(_05043_),
    .A2(_05365_),
    .B1(_05366_),
    .B2(_05367_),
    .C1(_05031_),
    .X(_05368_));
 sky130_fd_sc_hd__a211o_1 _12179_ (.A1(_05061_),
    .A2(_05364_),
    .B1(_05368_),
    .C1(_04948_),
    .X(_05369_));
 sky130_fd_sc_hd__o311a_1 _12180_ (.A1(_04964_),
    .A2(_05357_),
    .A3(_05361_),
    .B1(_04940_),
    .C1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__a31o_1 _12181_ (.A1(_05030_),
    .A2(_05343_),
    .A3(_05353_),
    .B1(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _12182_ (.A0(_05335_),
    .A1(_05371_),
    .S(_04945_),
    .X(_05372_));
 sky130_fd_sc_hd__a21o_1 _12183_ (.A1(\rbzero.row_render.side ),
    .A2(_05153_),
    .B1(_05147_),
    .X(_05373_));
 sky130_fd_sc_hd__or2_1 _12184_ (.A(_05143_),
    .B(\rbzero.row_render.wall[1] ),
    .X(_05374_));
 sky130_fd_sc_hd__o211a_1 _12185_ (.A1(_05157_),
    .A2(_05163_),
    .B1(_05373_),
    .C1(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__nand2_1 _12186_ (.A(\rbzero.row_render.texu[4] ),
    .B(_05030_),
    .Y(_05376_));
 sky130_fd_sc_hd__or2_1 _12187_ (.A(\rbzero.row_render.texu[4] ),
    .B(_05030_),
    .X(_05377_));
 sky130_fd_sc_hd__a31o_1 _12188_ (.A1(_05144_),
    .A2(_05376_),
    .A3(_05377_),
    .B1(_05028_),
    .X(_05378_));
 sky130_fd_sc_hd__o221a_1 _12189_ (.A1(net42),
    .A2(_05372_),
    .B1(_05375_),
    .B2(_05378_),
    .C1(_05025_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _12190_ (.A0(\rbzero.color_sky[1] ),
    .A1(\rbzero.color_floor[1] ),
    .S(_04970_),
    .X(_05380_));
 sky130_fd_sc_hd__and2b_1 _12191_ (.A_N(_05025_),
    .B(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__or2_1 _12192_ (.A(_04853_),
    .B(_04837_),
    .X(_05382_));
 sky130_fd_sc_hd__xnor2_1 _12193_ (.A(_04787_),
    .B(_04586_),
    .Y(_05383_));
 sky130_fd_sc_hd__a22o_1 _12194_ (.A1(\gpout0.vpos[4] ),
    .A2(_04553_),
    .B1(_04587_),
    .B2(_04793_),
    .X(_05384_));
 sky130_fd_sc_hd__a221o_1 _12195_ (.A1(_04802_),
    .A2(_04555_),
    .B1(_04549_),
    .B2(_04822_),
    .C1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__a2bb2o_1 _12196_ (.A1_N(_04788_),
    .A2_N(_04554_),
    .B1(_04835_),
    .B2(\gpout0.vpos[6] ),
    .X(_05386_));
 sky130_fd_sc_hd__or3_1 _12197_ (.A(_05383_),
    .B(_05385_),
    .C(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__or3b_1 _12198_ (.A(_04106_),
    .B(_04546_),
    .C_N(_04764_),
    .X(_05388_));
 sky130_fd_sc_hd__or4b_1 _12199_ (.A(\gpout0.vpos[7] ),
    .B(_04778_),
    .C(_04793_),
    .D_N(\gpout0.vpos[4] ),
    .X(_05389_));
 sky130_fd_sc_hd__or4_1 _12200_ (.A(_04802_),
    .B(_04835_),
    .C(_05388_),
    .D(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__nand2_1 _12201_ (.A(_05387_),
    .B(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__and3_1 _12202_ (.A(_04106_),
    .B(_04553_),
    .C(_04547_),
    .X(_05392_));
 sky130_fd_sc_hd__a2bb2o_1 _12203_ (.A1_N(_04106_),
    .A2_N(_04870_),
    .B1(_05392_),
    .B2(_04550_),
    .X(_05393_));
 sky130_fd_sc_hd__xnor2_1 _12204_ (.A(_04778_),
    .B(_04835_),
    .Y(_05394_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(_04785_),
    .B(_04786_),
    .Y(_05395_));
 sky130_fd_sc_hd__nor2_1 _12206_ (.A(\gpout0.vpos[3] ),
    .B(\gpout0.hpos[3] ),
    .Y(_05396_));
 sky130_fd_sc_hd__a31o_1 _12207_ (.A1(_04778_),
    .A2(_04587_),
    .A3(_05395_),
    .B1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__a2bb2o_1 _12208_ (.A1_N(_04793_),
    .A2_N(_04866_),
    .B1(_05394_),
    .B2(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__and3_1 _12209_ (.A(_04788_),
    .B(_04793_),
    .C(_05178_),
    .X(_05399_));
 sky130_fd_sc_hd__a2bb2o_1 _12210_ (.A1_N(\gpout0.vpos[4] ),
    .A2_N(_04587_),
    .B1(\gpout0.hpos[3] ),
    .B2(\gpout0.vpos[3] ),
    .X(_05400_));
 sky130_fd_sc_hd__or4_1 _12211_ (.A(\gpout0.vpos[6] ),
    .B(_04553_),
    .C(_05396_),
    .D(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__a211o_1 _12212_ (.A1(_04788_),
    .A2(_04587_),
    .B1(_05394_),
    .C1(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__or4b_2 _12213_ (.A(_05393_),
    .B(_05398_),
    .C(_05399_),
    .D_N(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__and3b_1 _12214_ (.A_N(_04827_),
    .B(_05391_),
    .C(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__o21ba_1 _12215_ (.A1(_05382_),
    .A2(_05404_),
    .B1_N(_04815_),
    .X(_05405_));
 sky130_fd_sc_hd__o32a_1 _12216_ (.A1(_05169_),
    .A2(_05379_),
    .A3(_05381_),
    .B1(_05405_),
    .B2(_04873_),
    .X(_05406_));
 sky130_fd_sc_hd__nor2_1 _12217_ (.A(_04784_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__o21ai_1 _12218_ (.A1(_05300_),
    .A2(_05407_),
    .B1(_05174_),
    .Y(_05408_));
 sky130_fd_sc_hd__o211ai_4 _12219_ (.A1(_04570_),
    .A2(_04768_),
    .B1(_05180_),
    .C1(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__inv_2 _12220_ (.A(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__mux2_2 _12221_ (.A0(\reg_rgb[7] ),
    .A1(_05410_),
    .S(_05182_),
    .X(_05411_));
 sky130_fd_sc_hd__clkbuf_1 _12222_ (.A(_05411_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_05048_),
    .X(_05412_));
 sky130_fd_sc_hd__buf_4 _12224_ (.A(_05078_),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _12225_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(_05412_),
    .A1(_05414_),
    .S(_05093_),
    .X(_05415_));
 sky130_fd_sc_hd__mux2_1 _12227_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_05413_),
    .X(_05416_));
 sky130_fd_sc_hd__and3_1 _12228_ (.A(\rbzero.tex_g0[51] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05417_));
 sky130_fd_sc_hd__a21o_1 _12229_ (.A1(\rbzero.tex_g0[50] ),
    .A2(_05085_),
    .B1(_05059_),
    .X(_05418_));
 sky130_fd_sc_hd__o221a_1 _12230_ (.A1(_05045_),
    .A2(_05416_),
    .B1(_05417_),
    .B2(_05418_),
    .C1(_05087_),
    .X(_05419_));
 sky130_fd_sc_hd__a211o_1 _12231_ (.A1(_05033_),
    .A2(_05415_),
    .B1(_05419_),
    .C1(_05064_),
    .X(_05420_));
 sky130_fd_sc_hd__mux2_1 _12232_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_05413_),
    .X(_05421_));
 sky130_fd_sc_hd__mux2_1 _12233_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_05413_),
    .X(_05422_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(_05421_),
    .A1(_05422_),
    .S(_05093_),
    .X(_05423_));
 sky130_fd_sc_hd__mux2_1 _12235_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_05035_),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _12236_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_05047_),
    .X(_05425_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(_05108_),
    .B(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__o211a_1 _12238_ (.A1(_05045_),
    .A2(_05424_),
    .B1(_05426_),
    .C1(_05081_),
    .X(_05427_));
 sky130_fd_sc_hd__a211o_1 _12239_ (.A1(_05062_),
    .A2(_05423_),
    .B1(_05427_),
    .C1(_05075_),
    .X(_05428_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_05413_),
    .X(_05429_));
 sky130_fd_sc_hd__mux2_1 _12241_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_05303_),
    .X(_05430_));
 sky130_fd_sc_hd__or2_1 _12242_ (.A(_05040_),
    .B(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__o211a_1 _12243_ (.A1(_05059_),
    .A2(_05429_),
    .B1(_05431_),
    .C1(_05081_),
    .X(_05432_));
 sky130_fd_sc_hd__buf_6 _12244_ (.A(_05303_),
    .X(_05433_));
 sky130_fd_sc_hd__mux2_1 _12245_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__and3_1 _12246_ (.A(\rbzero.tex_g0[43] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05435_));
 sky130_fd_sc_hd__a21o_1 _12247_ (.A1(\rbzero.tex_g0[42] ),
    .A2(_05085_),
    .B1(_05108_),
    .X(_05436_));
 sky130_fd_sc_hd__o221a_1 _12248_ (.A1(_05041_),
    .A2(_05434_),
    .B1(_05435_),
    .B2(_05436_),
    .C1(_05087_),
    .X(_05437_));
 sky130_fd_sc_hd__mux2_1 _12249_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_05034_),
    .X(_05438_));
 sky130_fd_sc_hd__mux2_1 _12250_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_05346_),
    .X(_05439_));
 sky130_fd_sc_hd__mux2_1 _12251_ (.A0(_05438_),
    .A1(_05439_),
    .S(_05040_),
    .X(_05440_));
 sky130_fd_sc_hd__mux2_1 _12252_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_05089_),
    .X(_05441_));
 sky130_fd_sc_hd__mux2_1 _12253_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04958_),
    .X(_05442_));
 sky130_fd_sc_hd__or2_1 _12254_ (.A(_05107_),
    .B(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__o211a_1 _12255_ (.A1(_05093_),
    .A2(_05441_),
    .B1(_05443_),
    .C1(_05032_),
    .X(_05444_));
 sky130_fd_sc_hd__a211o_1 _12256_ (.A1(_05062_),
    .A2(_05440_),
    .B1(_05444_),
    .C1(_05137_),
    .X(_05445_));
 sky130_fd_sc_hd__o311a_1 _12257_ (.A1(_05075_),
    .A2(_05432_),
    .A3(_05437_),
    .B1(_04941_),
    .C1(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__a31o_1 _12258_ (.A1(_05030_),
    .A2(_05420_),
    .A3(_05428_),
    .B1(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__and2_1 _12259_ (.A(\rbzero.tex_g0[22] ),
    .B(_05413_),
    .X(_05448_));
 sky130_fd_sc_hd__a31o_1 _12260_ (.A1(\rbzero.tex_g0[23] ),
    .A2(_05050_),
    .A3(_05052_),
    .B1(_05058_),
    .X(_05449_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_05056_),
    .X(_05450_));
 sky130_fd_sc_hd__o221a_1 _12262_ (.A1(_05448_),
    .A2(_05449_),
    .B1(_05450_),
    .B2(_05093_),
    .C1(_05081_),
    .X(_05451_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_05056_),
    .X(_05452_));
 sky130_fd_sc_hd__and3_1 _12264_ (.A(\rbzero.tex_g0[19] ),
    .B(_05050_),
    .C(_05052_),
    .X(_05453_));
 sky130_fd_sc_hd__a21o_1 _12265_ (.A1(\rbzero.tex_g0[18] ),
    .A2(_05070_),
    .B1(_05108_),
    .X(_05454_));
 sky130_fd_sc_hd__o221a_1 _12266_ (.A1(_05093_),
    .A2(_05452_),
    .B1(_05453_),
    .B2(_05454_),
    .C1(_05061_),
    .X(_05455_));
 sky130_fd_sc_hd__mux2_1 _12267_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_05413_),
    .X(_05456_));
 sky130_fd_sc_hd__and3_1 _12268_ (.A(\rbzero.tex_g0[27] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05457_));
 sky130_fd_sc_hd__a21o_1 _12269_ (.A1(\rbzero.tex_g0[26] ),
    .A2(_05085_),
    .B1(_05059_),
    .X(_05458_));
 sky130_fd_sc_hd__o221a_1 _12270_ (.A1(_05041_),
    .A2(_05456_),
    .B1(_05457_),
    .B2(_05458_),
    .C1(_05087_),
    .X(_05459_));
 sky130_fd_sc_hd__mux2_1 _12271_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_05078_),
    .X(_05460_));
 sky130_fd_sc_hd__mux2_1 _12272_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_05078_),
    .X(_05461_));
 sky130_fd_sc_hd__mux2_1 _12273_ (.A0(_05460_),
    .A1(_05461_),
    .S(_05058_),
    .X(_05462_));
 sky130_fd_sc_hd__a21o_1 _12274_ (.A1(_05033_),
    .A2(_05462_),
    .B1(_05118_),
    .X(_05463_));
 sky130_fd_sc_hd__o32a_1 _12275_ (.A1(_05064_),
    .A2(_05451_),
    .A3(_05455_),
    .B1(_05459_),
    .B2(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__and2_1 _12276_ (.A(\rbzero.tex_g0[14] ),
    .B(_05070_),
    .X(_05465_));
 sky130_fd_sc_hd__a31o_1 _12277_ (.A1(\rbzero.tex_g0[15] ),
    .A2(_05051_),
    .A3(_05053_),
    .B1(_05058_),
    .X(_05466_));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_05433_),
    .X(_05467_));
 sky130_fd_sc_hd__o221a_1 _12279_ (.A1(_05465_),
    .A2(_05466_),
    .B1(_05467_),
    .B2(_05041_),
    .C1(_05081_),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _12280_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_05303_),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_1 _12281_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_05303_),
    .X(_05470_));
 sky130_fd_sc_hd__mux2_1 _12282_ (.A0(_05469_),
    .A1(_05470_),
    .S(_05351_),
    .X(_05471_));
 sky130_fd_sc_hd__a21o_1 _12283_ (.A1(_05087_),
    .A2(_05471_),
    .B1(_04948_),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_05055_),
    .X(_05473_));
 sky130_fd_sc_hd__mux2_1 _12285_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_05055_),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_1 _12286_ (.A0(_05473_),
    .A1(_05474_),
    .S(_05351_),
    .X(_05475_));
 sky130_fd_sc_hd__mux2_1 _12287_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_05055_),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_05055_),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _12289_ (.A0(_05476_),
    .A1(_05477_),
    .S(_05058_),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(_05475_),
    .A1(_05478_),
    .S(_05081_),
    .X(_05479_));
 sky130_fd_sc_hd__o22a_1 _12291_ (.A1(_05468_),
    .A2(_05472_),
    .B1(_05479_),
    .B2(_05064_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(_05464_),
    .A1(_05480_),
    .S(_04941_),
    .X(_05481_));
 sky130_fd_sc_hd__mux2_1 _12293_ (.A0(_05447_),
    .A1(_05481_),
    .S(_04945_),
    .X(_05482_));
 sky130_fd_sc_hd__a41o_1 _12294_ (.A1(_05045_),
    .A2(_04967_),
    .A3(_05033_),
    .A4(_05152_),
    .B1(_05146_),
    .X(_05483_));
 sky130_fd_sc_hd__o31a_1 _12295_ (.A1(_05142_),
    .A2(_05143_),
    .A3(_05161_),
    .B1(_05374_),
    .X(_05484_));
 sky130_fd_sc_hd__a21boi_1 _12296_ (.A1(_05155_),
    .A2(_05483_),
    .B1_N(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__o21ai_1 _12297_ (.A1(_05145_),
    .A2(_05485_),
    .B1(_05025_),
    .Y(_05486_));
 sky130_fd_sc_hd__a21oi_1 _12298_ (.A1(_05028_),
    .A2(_05482_),
    .B1(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_04970_),
    .X(_05488_));
 sky130_fd_sc_hd__nor2_1 _12300_ (.A(_05025_),
    .B(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__nand2_1 _12301_ (.A(_05169_),
    .B(_04812_),
    .Y(_05490_));
 sky130_fd_sc_hd__o311a_1 _12302_ (.A1(_05169_),
    .A2(_05487_),
    .A3(_05489_),
    .B1(_05490_),
    .C1(_05171_),
    .X(_05491_));
 sky130_fd_sc_hd__o21ai_1 _12303_ (.A1(_04792_),
    .A2(_05491_),
    .B1(_05174_),
    .Y(_05492_));
 sky130_fd_sc_hd__o211a_2 _12304_ (.A1(_04563_),
    .A2(_04768_),
    .B1(_05180_),
    .C1(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_2 _12305_ (.A0(\reg_rgb[14] ),
    .A1(_05493_),
    .S(_05182_),
    .X(_05494_));
 sky130_fd_sc_hd__clkbuf_1 _12306_ (.A(_05494_),
    .X(net65));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_05433_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _12308_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_05055_),
    .X(_05496_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_05055_),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _12310_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04957_),
    .X(_05498_));
 sky130_fd_sc_hd__or3_1 _12311_ (.A(_05039_),
    .B(_04950_),
    .C(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__o221a_1 _12312_ (.A1(_05158_),
    .A2(_05496_),
    .B1(_05497_),
    .B2(_05307_),
    .C1(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__o211a_1 _12313_ (.A1(_04966_),
    .A2(_05495_),
    .B1(_05500_),
    .C1(_04948_),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _12314_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_05413_),
    .X(_05502_));
 sky130_fd_sc_hd__buf_6 _12315_ (.A(_05302_),
    .X(_05503_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(\rbzero.tex_g1[63] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__mux2_1 _12317_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_05503_),
    .X(_05505_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04957_),
    .X(_05506_));
 sky130_fd_sc_hd__or3_1 _12319_ (.A(_05039_),
    .B(_04950_),
    .C(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__o221a_1 _12320_ (.A1(_05159_),
    .A2(_05504_),
    .B1(_05505_),
    .B2(_05307_),
    .C1(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__o211a_1 _12321_ (.A1(_04966_),
    .A2(_05502_),
    .B1(_05508_),
    .C1(_04964_),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_05070_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _12323_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_05078_),
    .X(_05511_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_05346_),
    .X(_05512_));
 sky130_fd_sc_hd__mux2_1 _12325_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_05302_),
    .X(_05513_));
 sky130_fd_sc_hd__or3_1 _12326_ (.A(_05039_),
    .B(_04955_),
    .C(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__o221a_1 _12327_ (.A1(_05159_),
    .A2(_05511_),
    .B1(_05512_),
    .B2(_05307_),
    .C1(_05514_),
    .X(_05515_));
 sky130_fd_sc_hd__o211a_1 _12328_ (.A1(_05148_),
    .A2(_05510_),
    .B1(_05515_),
    .C1(_05118_),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_1 _12329_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_05034_),
    .X(_05517_));
 sky130_fd_sc_hd__or2_1 _12330_ (.A(_04965_),
    .B(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__mux2_1 _12331_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_05305_),
    .X(_05519_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_05047_),
    .X(_05520_));
 sky130_fd_sc_hd__mux2_1 _12333_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_05302_),
    .X(_05521_));
 sky130_fd_sc_hd__or3_1 _12334_ (.A(_05039_),
    .B(_04955_),
    .C(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__o221a_1 _12335_ (.A1(_05159_),
    .A2(_05519_),
    .B1(_05520_),
    .B2(_05307_),
    .C1(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__a31o_1 _12336_ (.A1(_05137_),
    .A2(_05518_),
    .A3(_05523_),
    .B1(_05029_),
    .X(_05524_));
 sky130_fd_sc_hd__o32a_1 _12337_ (.A1(_04941_),
    .A2(_05501_),
    .A3(_05509_),
    .B1(_05516_),
    .B2(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__mux2_1 _12338_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_05303_),
    .X(_05526_));
 sky130_fd_sc_hd__mux2_1 _12339_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_05303_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(_05526_),
    .A1(_05527_),
    .S(_05351_),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _12341_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_05503_),
    .X(_05529_));
 sky130_fd_sc_hd__a31o_1 _12342_ (.A1(\rbzero.tex_g1[23] ),
    .A2(_05050_),
    .A3(_05052_),
    .B1(_05107_),
    .X(_05530_));
 sky130_fd_sc_hd__and2_1 _12343_ (.A(\rbzero.tex_g1[22] ),
    .B(_05089_),
    .X(_05531_));
 sky130_fd_sc_hd__o221a_1 _12344_ (.A1(_05040_),
    .A2(_05529_),
    .B1(_05530_),
    .B2(_05531_),
    .C1(_05031_),
    .X(_05532_));
 sky130_fd_sc_hd__a211o_1 _12345_ (.A1(_05087_),
    .A2(_05528_),
    .B1(_05532_),
    .C1(_05137_),
    .X(_05533_));
 sky130_fd_sc_hd__mux2_1 _12346_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_05503_),
    .X(_05534_));
 sky130_fd_sc_hd__or2_1 _12347_ (.A(_05058_),
    .B(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__mux2_1 _12348_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_05305_),
    .X(_05536_));
 sky130_fd_sc_hd__o21a_1 _12349_ (.A1(_05040_),
    .A2(_05536_),
    .B1(_05031_),
    .X(_05537_));
 sky130_fd_sc_hd__mux2_1 _12350_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_05503_),
    .X(_05538_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_05503_),
    .X(_05539_));
 sky130_fd_sc_hd__mux2_1 _12352_ (.A0(_05538_),
    .A1(_05539_),
    .S(_05351_),
    .X(_05540_));
 sky130_fd_sc_hd__a221o_1 _12353_ (.A1(_05535_),
    .A2(_05537_),
    .B1(_05540_),
    .B2(_05061_),
    .C1(_04948_),
    .X(_05541_));
 sky130_fd_sc_hd__mux2_1 _12354_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[0] ),
    .S(_05055_),
    .X(_05542_));
 sky130_fd_sc_hd__and2_1 _12355_ (.A(\rbzero.tex_g1[2] ),
    .B(_05346_),
    .X(_05543_));
 sky130_fd_sc_hd__a31o_1 _12356_ (.A1(\rbzero.tex_g1[3] ),
    .A2(_04915_),
    .A3(_04956_),
    .B1(_04954_),
    .X(_05544_));
 sky130_fd_sc_hd__o221a_1 _12357_ (.A1(_05351_),
    .A2(_05542_),
    .B1(_05543_),
    .B2(_05544_),
    .C1(_04951_),
    .X(_05545_));
 sky130_fd_sc_hd__mux2_1 _12358_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_05503_),
    .X(_05546_));
 sky130_fd_sc_hd__a21o_1 _12359_ (.A1(\rbzero.tex_g1[6] ),
    .A2(_05069_),
    .B1(_05107_),
    .X(_05547_));
 sky130_fd_sc_hd__and3_1 _12360_ (.A(\rbzero.tex_g1[7] ),
    .B(_04915_),
    .C(_04956_),
    .X(_05548_));
 sky130_fd_sc_hd__o221a_1 _12361_ (.A1(_05040_),
    .A2(_05546_),
    .B1(_05547_),
    .B2(_05548_),
    .C1(_05031_),
    .X(_05549_));
 sky130_fd_sc_hd__mux2_1 _12362_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_05046_),
    .X(_05550_));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_05046_),
    .X(_05551_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(_05550_),
    .A1(_05551_),
    .S(_05107_),
    .X(_05552_));
 sky130_fd_sc_hd__mux2_1 _12365_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_05302_),
    .X(_05553_));
 sky130_fd_sc_hd__and3_1 _12366_ (.A(\rbzero.tex_g1[11] ),
    .B(_04915_),
    .C(_04956_),
    .X(_05554_));
 sky130_fd_sc_hd__a21o_1 _12367_ (.A1(\rbzero.tex_g1[10] ),
    .A2(_04958_),
    .B1(_04954_),
    .X(_05555_));
 sky130_fd_sc_hd__o221a_1 _12368_ (.A1(_05043_),
    .A2(_05553_),
    .B1(_05554_),
    .B2(_05555_),
    .C1(_04951_),
    .X(_05556_));
 sky130_fd_sc_hd__a211o_1 _12369_ (.A1(_05032_),
    .A2(_05552_),
    .B1(_05556_),
    .C1(_04948_),
    .X(_05557_));
 sky130_fd_sc_hd__o311a_1 _12370_ (.A1(_04964_),
    .A2(_05545_),
    .A3(_05549_),
    .B1(_04940_),
    .C1(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__a31o_1 _12371_ (.A1(_05030_),
    .A2(_05533_),
    .A3(_05541_),
    .B1(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(_05525_),
    .A1(_05559_),
    .S(_04945_),
    .X(_05560_));
 sky130_fd_sc_hd__a21oi_1 _12373_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_05033_),
    .B1(_05374_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21a_1 _12374_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_05033_),
    .B1(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__a41o_1 _12375_ (.A1(\rbzero.row_render.side ),
    .A2(_05143_),
    .A3(\rbzero.row_render.wall[1] ),
    .A4(_05153_),
    .B1(_05028_),
    .X(_05563_));
 sky130_fd_sc_hd__o221a_1 _12376_ (.A1(net42),
    .A2(_05560_),
    .B1(_05562_),
    .B2(_05563_),
    .C1(_05025_),
    .X(_05564_));
 sky130_fd_sc_hd__mux2_1 _12377_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_04970_),
    .X(_05565_));
 sky130_fd_sc_hd__and2b_1 _12378_ (.A_N(_05024_),
    .B(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__and2b_1 _12379_ (.A_N(_04815_),
    .B(_05403_),
    .X(_05567_));
 sky130_fd_sc_hd__nor2_1 _12380_ (.A(_04827_),
    .B(_05382_),
    .Y(_05568_));
 sky130_fd_sc_hd__and3b_1 _12381_ (.A_N(_05391_),
    .B(_05567_),
    .C(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__o32a_1 _12382_ (.A1(_05169_),
    .A2(_05564_),
    .A3(_05566_),
    .B1(_04873_),
    .B2(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__nor2_1 _12383_ (.A(_04784_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__o21ai_1 _12384_ (.A1(_05300_),
    .A2(_05571_),
    .B1(_05174_),
    .Y(_05572_));
 sky130_fd_sc_hd__o211a_4 _12385_ (.A1(\rbzero.trace_state[3] ),
    .A2(_04768_),
    .B1(_05180_),
    .C1(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__mux2_2 _12386_ (.A0(\reg_rgb[15] ),
    .A1(_05573_),
    .S(_05182_),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_1 _12387_ (.A(_05574_),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_04970_),
    .X(_05575_));
 sky130_fd_sc_hd__o21a_1 _12389_ (.A1(_05057_),
    .A2(_05160_),
    .B1(_05154_),
    .X(_05576_));
 sky130_fd_sc_hd__o211a_1 _12390_ (.A1(_05373_),
    .A2(_05576_),
    .B1(_05484_),
    .C1(_05163_),
    .X(_05577_));
 sky130_fd_sc_hd__mux2_1 _12391_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_05057_),
    .X(_05578_));
 sky130_fd_sc_hd__mux2_1 _12392_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_05035_),
    .X(_05579_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_05070_),
    .X(_05580_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_05346_),
    .X(_05581_));
 sky130_fd_sc_hd__or3_1 _12395_ (.A(_05044_),
    .B(_04951_),
    .C(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__o221a_1 _12396_ (.A1(_05160_),
    .A2(_05579_),
    .B1(_05580_),
    .B2(_05322_),
    .C1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__o211a_1 _12397_ (.A1(_05148_),
    .A2(_05578_),
    .B1(_05583_),
    .C1(_05075_),
    .X(_05584_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_05057_),
    .X(_05585_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_05085_),
    .X(_05586_));
 sky130_fd_sc_hd__mux2_1 _12400_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_05085_),
    .X(_05587_));
 sky130_fd_sc_hd__o22a_1 _12401_ (.A1(_05148_),
    .A2(_05586_),
    .B1(_05587_),
    .B2(_05322_),
    .X(_05588_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_05085_),
    .X(_05589_));
 sky130_fd_sc_hd__o31a_1 _12403_ (.A1(_05045_),
    .A2(_05062_),
    .A3(_05589_),
    .B1(_05064_),
    .X(_05590_));
 sky130_fd_sc_hd__o211a_1 _12404_ (.A1(_05160_),
    .A2(_05585_),
    .B1(_05588_),
    .C1(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__nor2_1 _12405_ (.A(_05584_),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__mux2_1 _12406_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_05048_),
    .X(_05593_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_05303_),
    .X(_05594_));
 sky130_fd_sc_hd__mux2_1 _12408_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_05305_),
    .X(_05595_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_05302_),
    .X(_05596_));
 sky130_fd_sc_hd__or3_1 _12410_ (.A(_05039_),
    .B(_04955_),
    .C(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__o221a_1 _12411_ (.A1(_05307_),
    .A2(_05594_),
    .B1(_05595_),
    .B2(_05159_),
    .C1(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__o211a_1 _12412_ (.A1(_04966_),
    .A2(_05593_),
    .B1(_05598_),
    .C1(_05118_),
    .X(_05599_));
 sky130_fd_sc_hd__mux2_1 _12413_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_05035_),
    .X(_05600_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_05034_),
    .X(_05601_));
 sky130_fd_sc_hd__mux2_1 _12415_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_05089_),
    .X(_05602_));
 sky130_fd_sc_hd__o22a_1 _12416_ (.A1(_04965_),
    .A2(_05601_),
    .B1(_05602_),
    .B2(_05322_),
    .X(_05603_));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_05089_),
    .X(_05604_));
 sky130_fd_sc_hd__o31a_1 _12418_ (.A1(_05093_),
    .A2(_04951_),
    .A3(_05604_),
    .B1(_04964_),
    .X(_05605_));
 sky130_fd_sc_hd__o211a_1 _12419_ (.A1(_05160_),
    .A2(_05600_),
    .B1(_05603_),
    .C1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__nor2_1 _12420_ (.A(_05599_),
    .B(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hd__or3b_1 _12421_ (.A(_05607_),
    .B(_04941_),
    .C_N(_04945_),
    .X(_05608_));
 sky130_fd_sc_hd__mux2_1 _12422_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_05057_),
    .X(_05609_));
 sky130_fd_sc_hd__mux2_1 _12423_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_05413_),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_05048_),
    .X(_05611_));
 sky130_fd_sc_hd__mux2_1 _12425_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_05503_),
    .X(_05612_));
 sky130_fd_sc_hd__or3_1 _12426_ (.A(_05040_),
    .B(_04951_),
    .C(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__o221a_1 _12427_ (.A1(_05160_),
    .A2(_05610_),
    .B1(_05611_),
    .B2(_04966_),
    .C1(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__o211ai_1 _12428_ (.A1(_05322_),
    .A2(_05609_),
    .B1(_05614_),
    .C1(_05064_),
    .Y(_05615_));
 sky130_fd_sc_hd__mux2_1 _12429_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_05057_),
    .X(_05616_));
 sky130_fd_sc_hd__mux2_1 _12430_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_05433_),
    .X(_05617_));
 sky130_fd_sc_hd__mux2_1 _12431_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_05413_),
    .X(_05618_));
 sky130_fd_sc_hd__mux2_1 _12432_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_05503_),
    .X(_05619_));
 sky130_fd_sc_hd__or3_1 _12433_ (.A(_05351_),
    .B(_04951_),
    .C(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__o221a_1 _12434_ (.A1(_05160_),
    .A2(_05617_),
    .B1(_05618_),
    .B2(_05322_),
    .C1(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__o211ai_1 _12435_ (.A1(_05148_),
    .A2(_05616_),
    .B1(_05621_),
    .C1(_05075_),
    .Y(_05622_));
 sky130_fd_sc_hd__mux2_1 _12436_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_05070_),
    .X(_05623_));
 sky130_fd_sc_hd__mux2_1 _12437_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_05346_),
    .X(_05624_));
 sky130_fd_sc_hd__mux2_1 _12438_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_05034_),
    .X(_05625_));
 sky130_fd_sc_hd__mux2_1 _12439_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_05302_),
    .X(_05626_));
 sky130_fd_sc_hd__or3_1 _12440_ (.A(_05039_),
    .B(_04955_),
    .C(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__o221a_1 _12441_ (.A1(_05307_),
    .A2(_05624_),
    .B1(_05625_),
    .B2(_05159_),
    .C1(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__o211a_1 _12442_ (.A1(_05148_),
    .A2(_05623_),
    .B1(_05628_),
    .C1(_05118_),
    .X(_05629_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_05085_),
    .X(_05630_));
 sky130_fd_sc_hd__mux2_1 _12444_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_05089_),
    .X(_05631_));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_05069_),
    .X(_05632_));
 sky130_fd_sc_hd__mux2_1 _12446_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_05046_),
    .X(_05633_));
 sky130_fd_sc_hd__or3_1 _12447_ (.A(_05043_),
    .B(_04955_),
    .C(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__o221a_1 _12448_ (.A1(_04966_),
    .A2(_05631_),
    .B1(_05632_),
    .B2(_05322_),
    .C1(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__o211a_1 _12449_ (.A1(_05160_),
    .A2(_05630_),
    .B1(_05635_),
    .C1(_05064_),
    .X(_05636_));
 sky130_fd_sc_hd__nor3_1 _12450_ (.A(_05030_),
    .B(_05629_),
    .C(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__a311o_1 _12451_ (.A1(_05030_),
    .A2(_05615_),
    .A3(_05622_),
    .B1(_04945_),
    .C1(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__o211ai_2 _12452_ (.A1(_04968_),
    .A2(_05592_),
    .B1(_05608_),
    .C1(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a2bb2o_1 _12453_ (.A1_N(_05145_),
    .A2_N(_05577_),
    .B1(_05639_),
    .B2(_05028_),
    .X(_05640_));
 sky130_fd_sc_hd__mux2_1 _12454_ (.A0(_05575_),
    .A1(_05640_),
    .S(_05025_),
    .X(_05641_));
 sky130_fd_sc_hd__o21ai_1 _12455_ (.A1(_05391_),
    .A2(_05403_),
    .B1(_05568_),
    .Y(_05642_));
 sky130_fd_sc_hd__or3b_1 _12456_ (.A(_04872_),
    .B(_04814_),
    .C_N(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__o211a_1 _12457_ (.A1(_05169_),
    .A2(_05641_),
    .B1(_05643_),
    .C1(_05490_),
    .X(_05644_));
 sky130_fd_sc_hd__nand2_1 _12458_ (.A(_05174_),
    .B(_05180_),
    .Y(_05645_));
 sky130_fd_sc_hd__nor2_1 _12459_ (.A(_04792_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__o21a_2 _12460_ (.A1(_04784_),
    .A2(_05644_),
    .B1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__mux2_2 _12461_ (.A0(\reg_rgb[22] ),
    .A1(_05647_),
    .S(_05182_),
    .X(_05648_));
 sky130_fd_sc_hd__clkbuf_1 _12462_ (.A(_05648_),
    .X(net67));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_05433_),
    .X(_05649_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_05433_),
    .X(_05650_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(_05649_),
    .A1(_05650_),
    .S(_05093_),
    .X(_05651_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_05056_),
    .X(_05652_));
 sky130_fd_sc_hd__and3_1 _12467_ (.A(\rbzero.tex_b1[35] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05653_));
 sky130_fd_sc_hd__a21o_1 _12468_ (.A1(\rbzero.tex_b1[34] ),
    .A2(_05070_),
    .B1(_05108_),
    .X(_05654_));
 sky130_fd_sc_hd__o221a_1 _12469_ (.A1(_05041_),
    .A2(_05652_),
    .B1(_05653_),
    .B2(_05654_),
    .C1(_05061_),
    .X(_05655_));
 sky130_fd_sc_hd__a211o_1 _12470_ (.A1(_05033_),
    .A2(_05651_),
    .B1(_05655_),
    .C1(_05064_),
    .X(_05656_));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_05433_),
    .X(_05657_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_05433_),
    .X(_05658_));
 sky130_fd_sc_hd__mux2_1 _12473_ (.A0(_05657_),
    .A1(_05658_),
    .S(_05093_),
    .X(_05659_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_05433_),
    .X(_05660_));
 sky130_fd_sc_hd__mux2_1 _12475_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_05303_),
    .X(_05661_));
 sky130_fd_sc_hd__or2_1 _12476_ (.A(_05108_),
    .B(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__o211a_1 _12477_ (.A1(_05041_),
    .A2(_05660_),
    .B1(_05662_),
    .C1(_05081_),
    .X(_05663_));
 sky130_fd_sc_hd__a211o_1 _12478_ (.A1(_05062_),
    .A2(_05659_),
    .B1(_05663_),
    .C1(_05075_),
    .X(_05664_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_05056_),
    .X(_05665_));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_05503_),
    .X(_05666_));
 sky130_fd_sc_hd__or2_1 _12481_ (.A(_05351_),
    .B(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__o211a_1 _12482_ (.A1(_05059_),
    .A2(_05665_),
    .B1(_05667_),
    .C1(_05081_),
    .X(_05668_));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_05056_),
    .X(_05669_));
 sky130_fd_sc_hd__and3_1 _12484_ (.A(\rbzero.tex_b1[59] ),
    .B(_05051_),
    .C(_05053_),
    .X(_05670_));
 sky130_fd_sc_hd__a21o_1 _12485_ (.A1(\rbzero.tex_b1[58] ),
    .A2(_05070_),
    .B1(_05108_),
    .X(_05671_));
 sky130_fd_sc_hd__o221a_1 _12486_ (.A1(_05041_),
    .A2(_05669_),
    .B1(_05670_),
    .B2(_05671_),
    .C1(_05061_),
    .X(_05672_));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_05305_),
    .X(_05673_));
 sky130_fd_sc_hd__mux2_1 _12488_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_05305_),
    .X(_05674_));
 sky130_fd_sc_hd__mux2_1 _12489_ (.A0(_05673_),
    .A1(_05674_),
    .S(_05351_),
    .X(_05675_));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_05346_),
    .X(_05676_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_05046_),
    .X(_05677_));
 sky130_fd_sc_hd__or2_1 _12492_ (.A(_05107_),
    .B(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__o211a_1 _12493_ (.A1(_05044_),
    .A2(_05676_),
    .B1(_05678_),
    .C1(_05032_),
    .X(_05679_));
 sky130_fd_sc_hd__a211o_1 _12494_ (.A1(_05087_),
    .A2(_05675_),
    .B1(_05679_),
    .C1(_05137_),
    .X(_05680_));
 sky130_fd_sc_hd__o311a_1 _12495_ (.A1(_05075_),
    .A2(_05668_),
    .A3(_05672_),
    .B1(_05030_),
    .C1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__a31o_1 _12496_ (.A1(_04941_),
    .A2(_05656_),
    .A3(_05664_),
    .B1(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_05057_),
    .X(_05683_));
 sky130_fd_sc_hd__mux2_1 _12498_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_05056_),
    .X(_05684_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_05433_),
    .X(_05685_));
 sky130_fd_sc_hd__mux2_1 _12500_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_05055_),
    .X(_05686_));
 sky130_fd_sc_hd__or3_1 _12501_ (.A(_05351_),
    .B(_04951_),
    .C(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__o221a_1 _12502_ (.A1(_05322_),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05160_),
    .C1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__o211a_1 _12503_ (.A1(_05148_),
    .A2(_05683_),
    .B1(_05688_),
    .C1(_05075_),
    .X(_05689_));
 sky130_fd_sc_hd__mux2_1 _12504_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_05057_),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_05048_),
    .X(_05691_));
 sky130_fd_sc_hd__mux2_1 _12506_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_05035_),
    .X(_05692_));
 sky130_fd_sc_hd__o22a_1 _12507_ (.A1(_04966_),
    .A2(_05691_),
    .B1(_05692_),
    .B2(_05322_),
    .X(_05693_));
 sky130_fd_sc_hd__mux2_1 _12508_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_05035_),
    .X(_05694_));
 sky130_fd_sc_hd__o31a_1 _12509_ (.A1(_05045_),
    .A2(_05061_),
    .A3(_05694_),
    .B1(_05137_),
    .X(_05695_));
 sky130_fd_sc_hd__o211a_1 _12510_ (.A1(_05160_),
    .A2(_05690_),
    .B1(_05693_),
    .C1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__mux2_1 _12511_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_05346_),
    .X(_05697_));
 sky130_fd_sc_hd__mux2_1 _12512_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_05346_),
    .X(_05698_));
 sky130_fd_sc_hd__mux2_1 _12513_ (.A0(_05697_),
    .A1(_05698_),
    .S(_05058_),
    .X(_05699_));
 sky130_fd_sc_hd__mux2_1 _12514_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_05346_),
    .X(_05700_));
 sky130_fd_sc_hd__and2_1 _12515_ (.A(\rbzero.tex_b1[22] ),
    .B(_05069_),
    .X(_05701_));
 sky130_fd_sc_hd__a31o_1 _12516_ (.A1(\rbzero.tex_b1[23] ),
    .A2(_05050_),
    .A3(_05052_),
    .B1(_05107_),
    .X(_05702_));
 sky130_fd_sc_hd__o221a_1 _12517_ (.A1(_05044_),
    .A2(_05700_),
    .B1(_05701_),
    .B2(_05702_),
    .C1(_05032_),
    .X(_05703_));
 sky130_fd_sc_hd__a211o_1 _12518_ (.A1(_05062_),
    .A2(_05699_),
    .B1(_05703_),
    .C1(_05137_),
    .X(_05704_));
 sky130_fd_sc_hd__mux2_1 _12519_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_05047_),
    .X(_05705_));
 sky130_fd_sc_hd__mux2_1 _12520_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_05047_),
    .X(_05706_));
 sky130_fd_sc_hd__mux2_1 _12521_ (.A0(_05705_),
    .A1(_05706_),
    .S(_05058_),
    .X(_05707_));
 sky130_fd_sc_hd__mux2_1 _12522_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_05078_),
    .X(_05708_));
 sky130_fd_sc_hd__and3_1 _12523_ (.A(\rbzero.tex_b1[27] ),
    .B(_05050_),
    .C(_05052_),
    .X(_05709_));
 sky130_fd_sc_hd__a21o_1 _12524_ (.A1(\rbzero.tex_b1[26] ),
    .A2(_05056_),
    .B1(_05107_),
    .X(_05710_));
 sky130_fd_sc_hd__o221a_1 _12525_ (.A1(_05044_),
    .A2(_05708_),
    .B1(_05709_),
    .B2(_05710_),
    .C1(_05061_),
    .X(_05711_));
 sky130_fd_sc_hd__a211o_1 _12526_ (.A1(_05033_),
    .A2(_05707_),
    .B1(_05711_),
    .C1(_05118_),
    .X(_05712_));
 sky130_fd_sc_hd__a21o_1 _12527_ (.A1(_05704_),
    .A2(_05712_),
    .B1(_04941_),
    .X(_05713_));
 sky130_fd_sc_hd__o31a_1 _12528_ (.A1(_05030_),
    .A2(_05689_),
    .A3(_05696_),
    .B1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__mux2_2 _12529_ (.A0(_05682_),
    .A1(_05714_),
    .S(_04945_),
    .X(_05715_));
 sky130_fd_sc_hd__a21oi_1 _12530_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04967_),
    .B1(_05374_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21a_1 _12531_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04967_),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__a21o_1 _12532_ (.A1(_05148_),
    .A2(_05152_),
    .B1(_05373_),
    .X(_05718_));
 sky130_fd_sc_hd__a31o_1 _12533_ (.A1(\rbzero.row_render.wall[1] ),
    .A2(_05163_),
    .A3(_05718_),
    .B1(_05028_),
    .X(_05719_));
 sky130_fd_sc_hd__o22ai_2 _12534_ (.A1(net42),
    .A2(_05715_),
    .B1(_05717_),
    .B2(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_04970_),
    .X(_05721_));
 sky130_fd_sc_hd__nor2_1 _12536_ (.A(_05025_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__a211o_1 _12537_ (.A1(_05025_),
    .A2(_05720_),
    .B1(_05722_),
    .C1(_05169_),
    .X(_05723_));
 sky130_fd_sc_hd__o311a_1 _12538_ (.A1(_04872_),
    .A2(_04815_),
    .A3(_05642_),
    .B1(_05723_),
    .C1(_05171_),
    .X(_05724_));
 sky130_fd_sc_hd__nor3_4 _12539_ (.A(_05300_),
    .B(_05645_),
    .C(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__mux2_2 _12540_ (.A0(\reg_rgb[23] ),
    .A1(_05725_),
    .S(_05182_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_1 _12541_ (.A(_05726_),
    .X(net68));
 sky130_fd_sc_hd__mux2_4 _12542_ (.A0(reg_vsync),
    .A1(_04565_),
    .S(_05182_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_1 _12543_ (.A(_05727_),
    .X(net75));
 sky130_fd_sc_hd__clkinv_2 _12544_ (.A(\rbzero.hsync ),
    .Y(_05728_));
 sky130_fd_sc_hd__mux2_2 _12545_ (.A0(reg_hsync),
    .A1(_05728_),
    .S(_05182_),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_1 _12546_ (.A(_05729_),
    .X(net63));
 sky130_fd_sc_hd__nor2_1 _12547_ (.A(net5),
    .B(net4),
    .Y(_05730_));
 sky130_fd_sc_hd__nor2_2 _12548_ (.A(net7),
    .B(net6),
    .Y(_05731_));
 sky130_fd_sc_hd__nor2_1 _12549_ (.A(net9),
    .B(net8),
    .Y(_05732_));
 sky130_fd_sc_hd__nand3_1 _12550_ (.A(_05730_),
    .B(_05731_),
    .C(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__buf_2 _12551_ (.A(net6),
    .X(_05734_));
 sky130_fd_sc_hd__buf_2 _12552_ (.A(net7),
    .X(_05735_));
 sky130_fd_sc_hd__a21o_1 _12553_ (.A1(net5),
    .A2(_05734_),
    .B1(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__nand2_1 _12554_ (.A(net8),
    .B(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__inv_2 _12555_ (.A(net5),
    .Y(_05738_));
 sky130_fd_sc_hd__clkbuf_4 _12556_ (.A(_04793_),
    .X(_05739_));
 sky130_fd_sc_hd__clkbuf_4 _12557_ (.A(net4),
    .X(_05740_));
 sky130_fd_sc_hd__mux4_1 _12558_ (.A0(\gpout0.vpos[2] ),
    .A1(_05739_),
    .A2(_04782_),
    .A3(_04775_),
    .S0(_05740_),
    .S1(_05734_),
    .X(_05741_));
 sky130_fd_sc_hd__clkbuf_4 _12559_ (.A(_04788_),
    .X(_05742_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(_05742_),
    .A1(_04787_),
    .S(_05740_),
    .X(_05743_));
 sky130_fd_sc_hd__clkbuf_4 _12561_ (.A(\gpout0.vpos[0] ),
    .X(_05744_));
 sky130_fd_sc_hd__buf_2 _12562_ (.A(\gpout0.vpos[1] ),
    .X(_05745_));
 sky130_fd_sc_hd__buf_2 _12563_ (.A(\gpout0.vpos[9] ),
    .X(_05746_));
 sky130_fd_sc_hd__mux4_1 _12564_ (.A0(_05744_),
    .A1(_05745_),
    .A2(_05177_),
    .A3(_05746_),
    .S0(_05740_),
    .S1(_05735_),
    .X(_05747_));
 sky130_fd_sc_hd__or2b_1 _12565_ (.A(_05747_),
    .B_N(_05734_),
    .X(_05748_));
 sky130_fd_sc_hd__o211a_1 _12566_ (.A1(_05734_),
    .A2(_05743_),
    .B1(_05748_),
    .C1(net5),
    .X(_05749_));
 sky130_fd_sc_hd__a21oi_1 _12567_ (.A1(_05738_),
    .A2(_05741_),
    .B1(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__nor2_1 _12568_ (.A(_05738_),
    .B(_05740_),
    .Y(_05751_));
 sky130_fd_sc_hd__inv_2 _12569_ (.A(net4),
    .Y(_05752_));
 sky130_fd_sc_hd__nor2_1 _12570_ (.A(_05738_),
    .B(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__and3_1 _12571_ (.A(_05200_),
    .B(_05731_),
    .C(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__a31o_1 _12572_ (.A1(net44),
    .A2(_05731_),
    .A3(_05751_),
    .B1(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__nor2_1 _12573_ (.A(net5),
    .B(_05752_),
    .Y(_05756_));
 sky130_fd_sc_hd__inv_2 _12574_ (.A(_05735_),
    .Y(_05757_));
 sky130_fd_sc_hd__a21o_1 _12575_ (.A1(net55),
    .A2(_05732_),
    .B1(net51),
    .X(_05758_));
 sky130_fd_sc_hd__a22o_1 _12576_ (.A1(net50),
    .A2(_05751_),
    .B1(_05758_),
    .B2(_05753_),
    .X(_05759_));
 sky130_fd_sc_hd__a22o_1 _12577_ (.A1(net52),
    .A2(_05730_),
    .B1(_05756_),
    .B2(net40),
    .X(_05760_));
 sky130_fd_sc_hd__a221o_1 _12578_ (.A1(net42),
    .A2(_05753_),
    .B1(_05751_),
    .B2(net41),
    .C1(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__and3b_1 _12579_ (.A_N(net6),
    .B(_05761_),
    .C(net7),
    .X(_05762_));
 sky130_fd_sc_hd__a31o_1 _12580_ (.A1(net43),
    .A2(_05730_),
    .A3(_05731_),
    .B1(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__a31o_1 _12581_ (.A1(_05757_),
    .A2(net6),
    .A3(_05759_),
    .B1(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__a31o_1 _12582_ (.A1(net46),
    .A2(_05756_),
    .A3(_05731_),
    .B1(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__or3_1 _12583_ (.A(net5),
    .B(_05740_),
    .C(_05179_),
    .X(_05766_));
 sky130_fd_sc_hd__o31a_1 _12584_ (.A1(net5),
    .A2(_05752_),
    .A3(_04560_),
    .B1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__or3b_1 _12585_ (.A(_05735_),
    .B(_05767_),
    .C_N(_05734_),
    .X(_05768_));
 sky130_fd_sc_hd__or3b_1 _12586_ (.A(_05755_),
    .B(_05765_),
    .C_N(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__inv_2 _12587_ (.A(net8),
    .Y(_05770_));
 sky130_fd_sc_hd__a2bb2o_1 _12588_ (.A1_N(_05737_),
    .A2_N(_05750_),
    .B1(_05769_),
    .B2(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__buf_6 _12589_ (.A(net55),
    .X(_05772_));
 sky130_fd_sc_hd__and3b_1 _12590_ (.A_N(_05735_),
    .B(_05734_),
    .C(_05753_),
    .X(_05773_));
 sky130_fd_sc_hd__a21o_1 _12591_ (.A1(_05735_),
    .A2(_05734_),
    .B1(net8),
    .X(_05774_));
 sky130_fd_sc_hd__mux4_1 _12592_ (.A0(_04588_),
    .A1(_04835_),
    .A2(_04554_),
    .A3(_04107_),
    .S0(_05740_),
    .S1(net5),
    .X(_05775_));
 sky130_fd_sc_hd__mux2_1 _12593_ (.A0(_04110_),
    .A1(_04111_),
    .S(_05740_),
    .X(_05776_));
 sky130_fd_sc_hd__mux4_1 _12594_ (.A0(_04103_),
    .A1(\gpout0.hpos[1] ),
    .A2(_04589_),
    .A3(_04586_),
    .S0(_05740_),
    .S1(net5),
    .X(_05777_));
 sky130_fd_sc_hd__mux2_1 _12595_ (.A0(_05776_),
    .A1(_05777_),
    .S(_05735_),
    .X(_05778_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(_05775_),
    .A1(_05778_),
    .S(_05734_),
    .X(_05779_));
 sky130_fd_sc_hd__and2_1 _12597_ (.A(net53),
    .B(_05730_),
    .X(_05780_));
 sky130_fd_sc_hd__a221o_1 _12598_ (.A1(net54),
    .A2(_05756_),
    .B1(_05751_),
    .B2(net56),
    .C1(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__and3b_1 _12599_ (.A_N(_05735_),
    .B(_05734_),
    .C(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__o211a_1 _12600_ (.A1(_05752_),
    .A2(_04187_),
    .B1(_05731_),
    .C1(_05738_),
    .X(_05783_));
 sky130_fd_sc_hd__and3_2 _12601_ (.A(clknet_leaf_41_i_clk),
    .B(_05731_),
    .C(_05751_),
    .X(_05784_));
 sky130_fd_sc_hd__a31o_2 _12602_ (.A1(\gpout0.clk_div[1] ),
    .A2(_05731_),
    .A3(_05753_),
    .B1(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__o31a_2 _12603_ (.A1(_05782_),
    .A2(_05783_),
    .A3(_05785_),
    .B1(_05732_),
    .X(_05786_));
 sky130_fd_sc_hd__a41o_2 _12604_ (.A1(net9),
    .A2(_05737_),
    .A3(_05774_),
    .A4(_05779_),
    .B1(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__a31o_2 _12605_ (.A1(_05772_),
    .A2(_05732_),
    .A3(_05773_),
    .B1(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(_05181_),
    .A1(_05410_),
    .S(_05740_),
    .X(_05789_));
 sky130_fd_sc_hd__mux4_1 _12607_ (.A0(_05493_),
    .A1(_05573_),
    .A2(_05647_),
    .A3(_05725_),
    .S0(_05740_),
    .S1(_05735_),
    .X(_05790_));
 sky130_fd_sc_hd__and2_1 _12608_ (.A(net8),
    .B(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__a31o_1 _12609_ (.A1(_05735_),
    .A2(_05770_),
    .A3(_05789_),
    .B1(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__and4b_1 _12610_ (.A_N(net9),
    .B(_05792_),
    .C(net5),
    .D(_05734_),
    .X(_05793_));
 sky130_fd_sc_hd__a211o_2 _12611_ (.A1(net9),
    .A2(_05771_),
    .B1(_05788_),
    .C1(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__o21a_2 _12612_ (.A1(_05493_),
    .A2(_05733_),
    .B1(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__mux2_2 _12613_ (.A0(\reg_gpout[0] ),
    .A1(clknet_1_0__leaf__05795_),
    .S(_05182_),
    .X(_05796_));
 sky130_fd_sc_hd__buf_1 _12614_ (.A(_05796_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 _12615_ (.A(net10),
    .X(_05797_));
 sky130_fd_sc_hd__or2_1 _12616_ (.A(_05797_),
    .B(_05181_),
    .X(_05798_));
 sky130_fd_sc_hd__inv_2 _12617_ (.A(net13),
    .Y(_05799_));
 sky130_fd_sc_hd__nor2_1 _12618_ (.A(_05799_),
    .B(net14),
    .Y(_05800_));
 sky130_fd_sc_hd__nand2_1 _12619_ (.A(_05797_),
    .B(_05409_),
    .Y(_05801_));
 sky130_fd_sc_hd__mux4_1 _12620_ (.A0(_05493_),
    .A1(_05573_),
    .A2(_05647_),
    .A3(_05725_),
    .S0(_05797_),
    .S1(net13),
    .X(_05802_));
 sky130_fd_sc_hd__a32o_1 _12621_ (.A1(_05798_),
    .A2(_05800_),
    .A3(_05801_),
    .B1(_05802_),
    .B2(net14),
    .X(_05803_));
 sky130_fd_sc_hd__buf_2 _12622_ (.A(net11),
    .X(_05804_));
 sky130_fd_sc_hd__buf_2 _12623_ (.A(net12),
    .X(_05805_));
 sky130_fd_sc_hd__and4b_1 _12624_ (.A_N(net15),
    .B(_05803_),
    .C(_05804_),
    .D(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__mux4_1 _12625_ (.A0(\gpout0.vpos[2] ),
    .A1(_05739_),
    .A2(_04782_),
    .A3(_04775_),
    .S0(_05797_),
    .S1(_05805_),
    .X(_05807_));
 sky130_fd_sc_hd__a21o_1 _12626_ (.A1(net13),
    .A2(_05807_),
    .B1(_05804_),
    .X(_05808_));
 sky130_fd_sc_hd__or2b_1 _12627_ (.A(_05746_),
    .B_N(net10),
    .X(_05809_));
 sky130_fd_sc_hd__o2111a_1 _12628_ (.A1(_05177_),
    .A2(_05797_),
    .B1(net13),
    .C1(_05805_),
    .D1(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__a211o_1 _12629_ (.A1(_04817_),
    .A2(net10),
    .B1(_05799_),
    .C1(_05805_),
    .X(_05811_));
 sky130_fd_sc_hd__o21ba_1 _12630_ (.A1(_05742_),
    .A2(_05797_),
    .B1_N(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__or2b_1 _12631_ (.A(_05745_),
    .B_N(net10),
    .X(_05813_));
 sky130_fd_sc_hd__o2111a_1 _12632_ (.A1(_05744_),
    .A2(_05797_),
    .B1(_05799_),
    .C1(_05805_),
    .D1(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__or4b_1 _12633_ (.A(_05810_),
    .B(_05812_),
    .C(_05814_),
    .D_N(_05804_),
    .X(_05815_));
 sky130_fd_sc_hd__inv_2 _12634_ (.A(_05805_),
    .Y(_05816_));
 sky130_fd_sc_hd__nor2b_2 _12635_ (.A(_05804_),
    .B_N(net10),
    .Y(_05817_));
 sky130_fd_sc_hd__or2_1 _12636_ (.A(_05804_),
    .B(net10),
    .X(_05818_));
 sky130_fd_sc_hd__o2bb2a_1 _12637_ (.A1_N(net72),
    .A2_N(_05817_),
    .B1(_05179_),
    .B2(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__or3_1 _12638_ (.A(net13),
    .B(_05816_),
    .C(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__nor2_2 _12639_ (.A(net13),
    .B(net12),
    .Y(_05821_));
 sky130_fd_sc_hd__and2_1 _12640_ (.A(_05804_),
    .B(net10),
    .X(_05822_));
 sky130_fd_sc_hd__and2b_1 _12641_ (.A_N(net10),
    .B(_05804_),
    .X(_05823_));
 sky130_fd_sc_hd__a22o_1 _12642_ (.A1(_05200_),
    .A2(_05822_),
    .B1(_05823_),
    .B2(net44),
    .X(_05824_));
 sky130_fd_sc_hd__nor2_2 _12643_ (.A(net11),
    .B(net10),
    .Y(_05825_));
 sky130_fd_sc_hd__a22o_1 _12644_ (.A1(net42),
    .A2(_05822_),
    .B1(_05823_),
    .B2(net41),
    .X(_05826_));
 sky130_fd_sc_hd__a221o_1 _12645_ (.A1(net52),
    .A2(_05825_),
    .B1(_05817_),
    .B2(net40),
    .C1(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__a22o_1 _12646_ (.A1(net51),
    .A2(_05822_),
    .B1(_05823_),
    .B2(net50),
    .X(_05828_));
 sky130_fd_sc_hd__and3_1 _12647_ (.A(net43),
    .B(_05825_),
    .C(_05821_),
    .X(_05829_));
 sky130_fd_sc_hd__a31o_1 _12648_ (.A1(net46),
    .A2(_05817_),
    .A3(_05821_),
    .B1(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__a31o_1 _12649_ (.A1(_05799_),
    .A2(_05805_),
    .A3(_05828_),
    .B1(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__a31o_1 _12650_ (.A1(net13),
    .A2(_05816_),
    .A3(_05827_),
    .B1(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__a21oi_1 _12651_ (.A1(_05821_),
    .A2(_05824_),
    .B1(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__a21oi_1 _12652_ (.A1(_05820_),
    .A2(_05833_),
    .B1(net14),
    .Y(_05834_));
 sky130_fd_sc_hd__mux4_1 _12653_ (.A0(_04588_),
    .A1(_04835_),
    .A2(_04554_),
    .A3(_04107_),
    .S0(_05797_),
    .S1(_05804_),
    .X(_05835_));
 sky130_fd_sc_hd__nand2_1 _12654_ (.A(_04583_),
    .B(_05817_),
    .Y(_05836_));
 sky130_fd_sc_hd__nor2_1 _12655_ (.A(_04103_),
    .B(_05818_),
    .Y(_05837_));
 sky130_fd_sc_hd__a221oi_1 _12656_ (.A1(_04548_),
    .A2(_05822_),
    .B1(_05823_),
    .B2(_04579_),
    .C1(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__a221o_1 _12657_ (.A1(_04110_),
    .A2(_05825_),
    .B1(_05817_),
    .B2(_04111_),
    .C1(_05816_),
    .X(_05839_));
 sky130_fd_sc_hd__and3_1 _12658_ (.A(_05799_),
    .B(net14),
    .C(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__a41o_1 _12659_ (.A1(_05805_),
    .A2(_05800_),
    .A3(_05836_),
    .A4(_05838_),
    .B1(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__o21a_1 _12660_ (.A1(_05805_),
    .A2(_05835_),
    .B1(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__a311o_1 _12661_ (.A1(net14),
    .A2(_05808_),
    .A3(_05815_),
    .B1(_05834_),
    .C1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__nor2_1 _12662_ (.A(net14),
    .B(net15),
    .Y(_05844_));
 sky130_fd_sc_hd__a21oi_2 _12663_ (.A1(_05804_),
    .A2(net128),
    .B1(_05797_),
    .Y(_05845_));
 sky130_fd_sc_hd__a221o_2 _12664_ (.A1(net49),
    .A2(_05817_),
    .B1(_05822_),
    .B2(\gpout1.clk_div[1] ),
    .C1(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__and2_1 _12665_ (.A(net56),
    .B(_05823_),
    .X(_05847_));
 sky130_fd_sc_hd__a22o_1 _12666_ (.A1(net53),
    .A2(_05825_),
    .B1(_05817_),
    .B2(net54),
    .X(_05848_));
 sky130_fd_sc_hd__and3_1 _12667_ (.A(_05804_),
    .B(_05797_),
    .C(_05772_),
    .X(_05849_));
 sky130_fd_sc_hd__o311a_1 _12668_ (.A1(_05847_),
    .A2(_05848_),
    .A3(_05849_),
    .B1(_05805_),
    .C1(_05799_),
    .X(_05850_));
 sky130_fd_sc_hd__a21o_2 _12669_ (.A1(_05821_),
    .A2(_05846_),
    .B1(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__a22o_2 _12670_ (.A1(net15),
    .A2(_05843_),
    .B1(_05844_),
    .B2(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__nand3_1 _12671_ (.A(_05825_),
    .B(_05821_),
    .C(_05844_),
    .Y(_05853_));
 sky130_fd_sc_hd__o22a_2 _12672_ (.A1(_05806_),
    .A2(_05852_),
    .B1(_05853_),
    .B2(_05573_),
    .X(_05854_));
 sky130_fd_sc_hd__mux2_2 _12673_ (.A0(\reg_gpout[1] ),
    .A1(clknet_1_1__leaf__05854_),
    .S(_05182_),
    .X(_05855_));
 sky130_fd_sc_hd__buf_1 _12674_ (.A(_05855_),
    .X(net58));
 sky130_fd_sc_hd__buf_2 _12675_ (.A(net17),
    .X(_05856_));
 sky130_fd_sc_hd__clkbuf_4 _12676_ (.A(net16),
    .X(_05857_));
 sky130_fd_sc_hd__or2_1 _12677_ (.A(_05856_),
    .B(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__or2_1 _12678_ (.A(net19),
    .B(net18),
    .X(_05859_));
 sky130_fd_sc_hd__or3_1 _12679_ (.A(net21),
    .B(net20),
    .C(_05181_),
    .X(_05860_));
 sky130_fd_sc_hd__or2_1 _12680_ (.A(_05857_),
    .B(_05181_),
    .X(_05861_));
 sky130_fd_sc_hd__inv_2 _12681_ (.A(net19),
    .Y(_05862_));
 sky130_fd_sc_hd__nor2_1 _12682_ (.A(_05862_),
    .B(net20),
    .Y(_05863_));
 sky130_fd_sc_hd__nand2_1 _12683_ (.A(_05857_),
    .B(_05409_),
    .Y(_05864_));
 sky130_fd_sc_hd__mux4_1 _12684_ (.A0(_05493_),
    .A1(_05573_),
    .A2(_05647_),
    .A3(_05725_),
    .S0(_05857_),
    .S1(net19),
    .X(_05865_));
 sky130_fd_sc_hd__a32o_1 _12685_ (.A1(_05861_),
    .A2(_05863_),
    .A3(_05864_),
    .B1(_05865_),
    .B2(net20),
    .X(_05866_));
 sky130_fd_sc_hd__buf_2 _12686_ (.A(net18),
    .X(_05867_));
 sky130_fd_sc_hd__and4b_1 _12687_ (.A_N(net21),
    .B(_05866_),
    .C(_05856_),
    .D(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__a21o_1 _12688_ (.A1(_05856_),
    .A2(_05867_),
    .B1(net19),
    .X(_05869_));
 sky130_fd_sc_hd__a21oi_1 _12689_ (.A1(net19),
    .A2(_05867_),
    .B1(net20),
    .Y(_05870_));
 sky130_fd_sc_hd__a21oi_1 _12690_ (.A1(net20),
    .A2(_05869_),
    .B1(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__mux4_1 _12691_ (.A0(_04588_),
    .A1(_04835_),
    .A2(_04554_),
    .A3(_04107_),
    .S0(_05857_),
    .S1(_05856_),
    .X(_05872_));
 sky130_fd_sc_hd__mux4_1 _12692_ (.A0(_04103_),
    .A1(\gpout0.hpos[1] ),
    .A2(_04589_),
    .A3(_04586_),
    .S0(net16),
    .S1(_05856_),
    .X(_05873_));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(_04110_),
    .A1(_04111_),
    .S(_05857_),
    .X(_05874_));
 sky130_fd_sc_hd__mux2_1 _12694_ (.A0(_05873_),
    .A1(_05874_),
    .S(_05862_),
    .X(_05875_));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(_05872_),
    .A1(_05875_),
    .S(_05867_),
    .X(_05876_));
 sky130_fd_sc_hd__and3_1 _12696_ (.A(net21),
    .B(_05871_),
    .C(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__inv_2 _12697_ (.A(net17),
    .Y(_05878_));
 sky130_fd_sc_hd__mux4_1 _12698_ (.A0(\gpout0.vpos[2] ),
    .A1(_05739_),
    .A2(_04782_),
    .A3(_04775_),
    .S0(_05857_),
    .S1(_05867_),
    .X(_05879_));
 sky130_fd_sc_hd__inv_2 _12699_ (.A(_05867_),
    .Y(_05880_));
 sky130_fd_sc_hd__mux4_1 _12700_ (.A0(_05744_),
    .A1(_05745_),
    .A2(_05177_),
    .A3(_05746_),
    .S0(net16),
    .S1(net19),
    .X(_05881_));
 sky130_fd_sc_hd__or2_1 _12701_ (.A(_05880_),
    .B(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__mux2_1 _12702_ (.A0(_04788_),
    .A1(_04787_),
    .S(_05857_),
    .X(_05883_));
 sky130_fd_sc_hd__o21a_1 _12703_ (.A1(_05867_),
    .A2(_05883_),
    .B1(_05856_),
    .X(_05884_));
 sky130_fd_sc_hd__a22o_1 _12704_ (.A1(_05878_),
    .A2(_05879_),
    .B1(_05882_),
    .B2(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__mux4_1 _12705_ (.A0(net52),
    .A1(net41),
    .A2(net40),
    .A3(net42),
    .S0(_05856_),
    .S1(_05857_),
    .X(_05886_));
 sky130_fd_sc_hd__nor2_1 _12706_ (.A(net19),
    .B(net18),
    .Y(_05887_));
 sky130_fd_sc_hd__nor2_1 _12707_ (.A(_05878_),
    .B(net16),
    .Y(_05888_));
 sky130_fd_sc_hd__nand2_1 _12708_ (.A(_05856_),
    .B(net16),
    .Y(_05889_));
 sky130_fd_sc_hd__nor2_1 _12709_ (.A(net21),
    .B(net20),
    .Y(_05890_));
 sky130_fd_sc_hd__a21oi_1 _12710_ (.A1(_05772_),
    .A2(_05890_),
    .B1(net51),
    .Y(_05891_));
 sky130_fd_sc_hd__o2bb2a_1 _12711_ (.A1_N(net50),
    .A2_N(_05888_),
    .B1(_05889_),
    .B2(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__nor2_1 _12712_ (.A(net19),
    .B(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__a211o_1 _12713_ (.A1(_05880_),
    .A2(_05886_),
    .B1(_05887_),
    .C1(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__and3b_1 _12714_ (.A_N(_05889_),
    .B(_05862_),
    .C(_05867_),
    .X(_05895_));
 sky130_fd_sc_hd__and2b_1 _12715_ (.A_N(net20),
    .B(net21),
    .X(_05896_));
 sky130_fd_sc_hd__a31o_1 _12716_ (.A1(_05772_),
    .A2(_05890_),
    .A3(_05895_),
    .B1(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__nor2_1 _12717_ (.A(net17),
    .B(net16),
    .Y(_05898_));
 sky130_fd_sc_hd__inv_2 _12718_ (.A(net16),
    .Y(_05899_));
 sky130_fd_sc_hd__nor2_1 _12719_ (.A(_05856_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__a221o_1 _12720_ (.A1(net43),
    .A2(_05898_),
    .B1(_05900_),
    .B2(net46),
    .C1(_05859_),
    .X(_05901_));
 sky130_fd_sc_hd__and2_1 _12721_ (.A(net53),
    .B(_05898_),
    .X(_05902_));
 sky130_fd_sc_hd__a221o_1 _12722_ (.A1(net56),
    .A2(_05888_),
    .B1(_05900_),
    .B2(net54),
    .C1(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__o211a_1 _12723_ (.A1(net47),
    .A2(_05899_),
    .B1(_05887_),
    .C1(_05878_),
    .X(_05904_));
 sky130_fd_sc_hd__a41o_1 _12724_ (.A1(_05856_),
    .A2(_05857_),
    .A3(\gpout2.clk_div[1] ),
    .A4(_05887_),
    .B1(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__a31o_2 _12725_ (.A1(clknet_1_0__leaf__04767_),
    .A2(_05888_),
    .A3(_05887_),
    .B1(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__a31o_2 _12726_ (.A1(_05862_),
    .A2(_05867_),
    .A3(_05903_),
    .B1(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__a32o_2 _12727_ (.A1(_05894_),
    .A2(_05897_),
    .A3(_05901_),
    .B1(_05907_),
    .B2(_05890_),
    .X(_05908_));
 sky130_fd_sc_hd__a41o_2 _12728_ (.A1(net21),
    .A2(net20),
    .A3(_05869_),
    .A4(_05885_),
    .B1(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__o2bb2a_1 _12729_ (.A1_N(net72),
    .A2_N(_05900_),
    .B1(_05179_),
    .B2(_05858_),
    .X(_05910_));
 sky130_fd_sc_hd__nor3b_1 _12730_ (.A(net19),
    .B(_05910_),
    .C_N(_05867_),
    .Y(_05911_));
 sky130_fd_sc_hd__nor3_1 _12731_ (.A(_05176_),
    .B(_05889_),
    .C(_05859_),
    .Y(_05912_));
 sky130_fd_sc_hd__a31o_1 _12732_ (.A1(net44),
    .A2(_05888_),
    .A3(_05887_),
    .B1(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__o21a_1 _12733_ (.A1(_05911_),
    .A2(_05913_),
    .B1(_05896_),
    .X(_05914_));
 sky130_fd_sc_hd__or4_2 _12734_ (.A(_05868_),
    .B(_05877_),
    .C(_05909_),
    .D(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__o31a_2 _12735_ (.A1(_05858_),
    .A2(_05859_),
    .A3(_05860_),
    .B1(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__mux2_2 _12736_ (.A0(\reg_gpout[2] ),
    .A1(clknet_1_1__leaf__05916_),
    .S(net45),
    .X(_05917_));
 sky130_fd_sc_hd__buf_1 _12737_ (.A(_05917_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 _12738_ (.A(net22),
    .X(_05918_));
 sky130_fd_sc_hd__or2_1 _12739_ (.A(_05918_),
    .B(_05181_),
    .X(_05919_));
 sky130_fd_sc_hd__buf_2 _12740_ (.A(net25),
    .X(_05920_));
 sky130_fd_sc_hd__inv_2 _12741_ (.A(net26),
    .Y(_05921_));
 sky130_fd_sc_hd__and2_1 _12742_ (.A(_05920_),
    .B(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__nand2_1 _12743_ (.A(_05918_),
    .B(_05409_),
    .Y(_05923_));
 sky130_fd_sc_hd__mux4_1 _12744_ (.A0(_05493_),
    .A1(_05573_),
    .A2(_05647_),
    .A3(_05725_),
    .S0(_05918_),
    .S1(_05920_),
    .X(_05924_));
 sky130_fd_sc_hd__a32o_1 _12745_ (.A1(_05919_),
    .A2(_05922_),
    .A3(_05923_),
    .B1(_05924_),
    .B2(net26),
    .X(_05925_));
 sky130_fd_sc_hd__buf_2 _12746_ (.A(net24),
    .X(_05926_));
 sky130_fd_sc_hd__and4b_1 _12747_ (.A_N(net27),
    .B(_05925_),
    .C(net23),
    .D(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__a21oi_1 _12748_ (.A1(net23),
    .A2(_05926_),
    .B1(_05920_),
    .Y(_05928_));
 sky130_fd_sc_hd__inv_2 _12749_ (.A(net23),
    .Y(_05929_));
 sky130_fd_sc_hd__mux4_1 _12750_ (.A0(\gpout0.vpos[2] ),
    .A1(_05739_),
    .A2(_04782_),
    .A3(_04775_),
    .S0(_05918_),
    .S1(_05926_),
    .X(_05930_));
 sky130_fd_sc_hd__inv_2 _12751_ (.A(_05926_),
    .Y(_05931_));
 sky130_fd_sc_hd__mux4_1 _12752_ (.A0(_05744_),
    .A1(_05745_),
    .A2(_05177_),
    .A3(_05746_),
    .S0(_05918_),
    .S1(_05920_),
    .X(_05932_));
 sky130_fd_sc_hd__or2_1 _12753_ (.A(_05931_),
    .B(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__mux2_1 _12754_ (.A0(_05742_),
    .A1(_04787_),
    .S(_05918_),
    .X(_05934_));
 sky130_fd_sc_hd__o21a_1 _12755_ (.A1(_05926_),
    .A2(_05934_),
    .B1(net23),
    .X(_05935_));
 sky130_fd_sc_hd__a22o_1 _12756_ (.A1(_05929_),
    .A2(_05930_),
    .B1(_05933_),
    .B2(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__and4b_1 _12757_ (.A_N(_05928_),
    .B(_05936_),
    .C(net27),
    .D(net26),
    .X(_05937_));
 sky130_fd_sc_hd__mux4_1 _12758_ (.A0(net52),
    .A1(net41),
    .A2(net40),
    .A3(net42),
    .S0(net23),
    .S1(_05918_),
    .X(_05938_));
 sky130_fd_sc_hd__nor2_1 _12759_ (.A(_05920_),
    .B(_05926_),
    .Y(_05939_));
 sky130_fd_sc_hd__nor2_1 _12760_ (.A(_05929_),
    .B(net22),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_1 _12761_ (.A(net23),
    .B(_05918_),
    .Y(_05941_));
 sky130_fd_sc_hd__nor2_1 _12762_ (.A(net27),
    .B(net26),
    .Y(_05942_));
 sky130_fd_sc_hd__a21oi_1 _12763_ (.A1(_05772_),
    .A2(_05942_),
    .B1(net51),
    .Y(_05943_));
 sky130_fd_sc_hd__o2bb2a_1 _12764_ (.A1_N(net50),
    .A2_N(_05940_),
    .B1(_05941_),
    .B2(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__nor2_1 _12765_ (.A(_05920_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__a211o_1 _12766_ (.A1(_05931_),
    .A2(_05938_),
    .B1(_05939_),
    .C1(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__and4bb_1 _12767_ (.A_N(_05941_),
    .B_N(_05920_),
    .C(_05926_),
    .D(_05942_),
    .X(_05947_));
 sky130_fd_sc_hd__a22o_1 _12768_ (.A1(net27),
    .A2(_05921_),
    .B1(_05947_),
    .B2(_05772_),
    .X(_05948_));
 sky130_fd_sc_hd__nor2_1 _12769_ (.A(net23),
    .B(_05918_),
    .Y(_05949_));
 sky130_fd_sc_hd__and2_1 _12770_ (.A(_05929_),
    .B(net22),
    .X(_05950_));
 sky130_fd_sc_hd__or2_1 _12771_ (.A(net25),
    .B(net24),
    .X(_05951_));
 sky130_fd_sc_hd__a221o_1 _12772_ (.A1(net43),
    .A2(_05949_),
    .B1(_05950_),
    .B2(net46),
    .C1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__and3_1 _12773_ (.A(_05946_),
    .B(_05948_),
    .C(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__a22o_1 _12774_ (.A1(_05926_),
    .A2(_05922_),
    .B1(_05928_),
    .B2(net26),
    .X(_05954_));
 sky130_fd_sc_hd__mux4_1 _12775_ (.A0(_04588_),
    .A1(_04835_),
    .A2(_04554_),
    .A3(_04107_),
    .S0(_05918_),
    .S1(net23),
    .X(_05955_));
 sky130_fd_sc_hd__mux2_1 _12776_ (.A0(_04110_),
    .A1(_04111_),
    .S(net22),
    .X(_05956_));
 sky130_fd_sc_hd__mux4_1 _12777_ (.A0(_04103_),
    .A1(_04711_),
    .A2(_04589_),
    .A3(_04586_),
    .S0(net22),
    .S1(net23),
    .X(_05957_));
 sky130_fd_sc_hd__mux2_1 _12778_ (.A0(_05956_),
    .A1(_05957_),
    .S(_05920_),
    .X(_05958_));
 sky130_fd_sc_hd__mux2_1 _12779_ (.A0(_05955_),
    .A1(_05958_),
    .S(_05926_),
    .X(_05959_));
 sky130_fd_sc_hd__a22o_1 _12780_ (.A1(net56),
    .A2(_05940_),
    .B1(_05950_),
    .B2(net54),
    .X(_05960_));
 sky130_fd_sc_hd__a21o_1 _12781_ (.A1(net53),
    .A2(_05949_),
    .B1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__and3b_1 _12782_ (.A_N(_05920_),
    .B(_05926_),
    .C(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__or2_1 _12783_ (.A(net23),
    .B(net22),
    .X(_05963_));
 sky130_fd_sc_hd__nor2_1 _12784_ (.A(_05963_),
    .B(_05951_),
    .Y(_05964_));
 sky130_fd_sc_hd__a31o_1 _12785_ (.A1(net48),
    .A2(_05950_),
    .A3(_05939_),
    .B1(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__nor2_1 _12786_ (.A(_05941_),
    .B(_05951_),
    .Y(_05966_));
 sky130_fd_sc_hd__a32o_2 _12787_ (.A1(clknet_1_0__leaf__04767_),
    .A2(_05940_),
    .A3(_05939_),
    .B1(_05966_),
    .B2(\gpout3.clk_div[1] ),
    .X(_05967_));
 sky130_fd_sc_hd__o31a_2 _12788_ (.A1(_05962_),
    .A2(_05965_),
    .A3(_05967_),
    .B1(_05942_),
    .X(_05968_));
 sky130_fd_sc_hd__a31o_2 _12789_ (.A1(net27),
    .A2(_05954_),
    .A3(_05959_),
    .B1(_05968_),
    .X(_05969_));
 sky130_fd_sc_hd__a32o_1 _12790_ (.A1(net44),
    .A2(_05940_),
    .A3(_05939_),
    .B1(_05966_),
    .B2(_05200_),
    .X(_05970_));
 sky130_fd_sc_hd__o2bb2a_1 _12791_ (.A1_N(net72),
    .A2_N(_05950_),
    .B1(_05179_),
    .B2(_05963_),
    .X(_05971_));
 sky130_fd_sc_hd__or3_1 _12792_ (.A(_05920_),
    .B(_05931_),
    .C(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__and2b_1 _12793_ (.A_N(_05970_),
    .B(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__or3b_1 _12794_ (.A(net26),
    .B(_05973_),
    .C_N(net27),
    .X(_05974_));
 sky130_fd_sc_hd__or3b_2 _12795_ (.A(_05953_),
    .B(_05969_),
    .C_N(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__nand3_1 _12796_ (.A(_05409_),
    .B(_05942_),
    .C(_05964_),
    .Y(_05976_));
 sky130_fd_sc_hd__o31a_2 _12797_ (.A1(_05927_),
    .A2(_05937_),
    .A3(_05975_),
    .B1(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__mux2_2 _12798_ (.A0(\reg_gpout[3] ),
    .A1(clknet_1_0__leaf__05977_),
    .S(net45),
    .X(_05978_));
 sky130_fd_sc_hd__buf_1 _12799_ (.A(_05978_),
    .X(net60));
 sky130_fd_sc_hd__buf_2 _12800_ (.A(net28),
    .X(_05979_));
 sky130_fd_sc_hd__or2_1 _12801_ (.A(_05979_),
    .B(_05181_),
    .X(_05980_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(_05979_),
    .B(_05409_),
    .Y(_05981_));
 sky130_fd_sc_hd__inv_2 _12803_ (.A(net31),
    .Y(_05982_));
 sky130_fd_sc_hd__nor2_1 _12804_ (.A(_05982_),
    .B(net32),
    .Y(_05983_));
 sky130_fd_sc_hd__mux4_1 _12805_ (.A0(_05493_),
    .A1(_05573_),
    .A2(_05647_),
    .A3(_05725_),
    .S0(_05979_),
    .S1(net31),
    .X(_05984_));
 sky130_fd_sc_hd__a32o_1 _12806_ (.A1(_05980_),
    .A2(_05981_),
    .A3(_05983_),
    .B1(_05984_),
    .B2(net32),
    .X(_05985_));
 sky130_fd_sc_hd__buf_2 _12807_ (.A(net29),
    .X(_05986_));
 sky130_fd_sc_hd__buf_2 _12808_ (.A(net30),
    .X(_05987_));
 sky130_fd_sc_hd__and4b_1 _12809_ (.A_N(net33),
    .B(_05985_),
    .C(_05986_),
    .D(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__and2b_1 _12810_ (.A_N(net32),
    .B(net33),
    .X(_05989_));
 sky130_fd_sc_hd__or2_1 _12811_ (.A(_05986_),
    .B(_05979_),
    .X(_05990_));
 sky130_fd_sc_hd__inv_2 _12812_ (.A(net29),
    .Y(_05991_));
 sky130_fd_sc_hd__and2_1 _12813_ (.A(_05991_),
    .B(net28),
    .X(_05992_));
 sky130_fd_sc_hd__a2bb2o_1 _12814_ (.A1_N(_05990_),
    .A2_N(_05179_),
    .B1(net72),
    .B2(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__nor2_1 _12815_ (.A(_05991_),
    .B(net28),
    .Y(_05994_));
 sky130_fd_sc_hd__nor2_1 _12816_ (.A(net31),
    .B(net30),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2_1 _12817_ (.A(_05986_),
    .B(_05979_),
    .Y(_05996_));
 sky130_fd_sc_hd__or2_1 _12818_ (.A(net31),
    .B(net30),
    .X(_05997_));
 sky130_fd_sc_hd__nor3_1 _12819_ (.A(_05176_),
    .B(_05996_),
    .C(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__a31o_1 _12820_ (.A1(net44),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__a31o_1 _12821_ (.A1(_05982_),
    .A2(_05987_),
    .A3(_05993_),
    .B1(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__nor2_1 _12822_ (.A(net32),
    .B(net33),
    .Y(_06001_));
 sky130_fd_sc_hd__a21oi_1 _12823_ (.A1(_05772_),
    .A2(_06001_),
    .B1(net51),
    .Y(_06002_));
 sky130_fd_sc_hd__o2bb2a_1 _12824_ (.A1_N(net50),
    .A2_N(_05994_),
    .B1(_05996_),
    .B2(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__o21ai_1 _12825_ (.A1(net31),
    .A2(_06003_),
    .B1(_05987_),
    .Y(_06004_));
 sky130_fd_sc_hd__mux4_1 _12826_ (.A0(net52),
    .A1(net41),
    .A2(net40),
    .A3(net42),
    .S0(_05986_),
    .S1(_05979_),
    .X(_06005_));
 sky130_fd_sc_hd__and3b_1 _12827_ (.A_N(_05996_),
    .B(_05982_),
    .C(_05987_),
    .X(_06006_));
 sky130_fd_sc_hd__a31o_1 _12828_ (.A1(_05772_),
    .A2(_06001_),
    .A3(_06006_),
    .B1(_05989_),
    .X(_06007_));
 sky130_fd_sc_hd__nor2_1 _12829_ (.A(net29),
    .B(net28),
    .Y(_06008_));
 sky130_fd_sc_hd__a221o_1 _12830_ (.A1(net46),
    .A2(_05992_),
    .B1(_06008_),
    .B2(net43),
    .C1(_05997_),
    .X(_06009_));
 sky130_fd_sc_hd__o211a_1 _12831_ (.A1(_05982_),
    .A2(_06005_),
    .B1(_06007_),
    .C1(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__a21oi_1 _12832_ (.A1(_05986_),
    .A2(_05987_),
    .B1(net31),
    .Y(_06011_));
 sky130_fd_sc_hd__mux4_1 _12833_ (.A0(\gpout0.vpos[2] ),
    .A1(_04793_),
    .A2(_04782_),
    .A3(_04775_),
    .S0(net28),
    .S1(net30),
    .X(_06012_));
 sky130_fd_sc_hd__mux4_1 _12834_ (.A0(\gpout0.vpos[0] ),
    .A1(\gpout0.vpos[1] ),
    .A2(_05177_),
    .A3(_05746_),
    .S0(net28),
    .S1(net31),
    .X(_06013_));
 sky130_fd_sc_hd__or2b_1 _12835_ (.A(_06013_),
    .B_N(_05987_),
    .X(_06014_));
 sky130_fd_sc_hd__mux2_1 _12836_ (.A0(_04788_),
    .A1(_04787_),
    .S(net28),
    .X(_06015_));
 sky130_fd_sc_hd__o21a_1 _12837_ (.A1(_05987_),
    .A2(_06015_),
    .B1(_05986_),
    .X(_06016_));
 sky130_fd_sc_hd__a22o_1 _12838_ (.A1(_05991_),
    .A2(_06012_),
    .B1(_06014_),
    .B2(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__and4b_1 _12839_ (.A_N(_06011_),
    .B(_06017_),
    .C(net32),
    .D(net33),
    .X(_06018_));
 sky130_fd_sc_hd__and2_1 _12840_ (.A(net53),
    .B(_06008_),
    .X(_06019_));
 sky130_fd_sc_hd__a221o_1 _12841_ (.A1(net56),
    .A2(_05994_),
    .B1(_05992_),
    .B2(net54),
    .C1(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__and3_1 _12842_ (.A(_05982_),
    .B(_05987_),
    .C(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__a211oi_1 _12843_ (.A1(_04776_),
    .A2(_05979_),
    .B1(_05997_),
    .C1(_05986_),
    .Y(_06022_));
 sky130_fd_sc_hd__and4_1 _12844_ (.A(_05986_),
    .B(_05979_),
    .C(\gpout4.clk_div[1] ),
    .D(_05995_),
    .X(_06023_));
 sky130_fd_sc_hd__a31o_2 _12845_ (.A1(clknet_1_0__leaf__04767_),
    .A2(_05994_),
    .A3(_05995_),
    .B1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__o31a_2 _12846_ (.A1(_06021_),
    .A2(_06022_),
    .A3(_06024_),
    .B1(_06001_),
    .X(_06025_));
 sky130_fd_sc_hd__a211o_2 _12847_ (.A1(_06004_),
    .A2(_06010_),
    .B1(_06018_),
    .C1(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__a22o_1 _12848_ (.A1(_05987_),
    .A2(_05983_),
    .B1(_06011_),
    .B2(net32),
    .X(_06027_));
 sky130_fd_sc_hd__mux4_1 _12849_ (.A0(_04588_),
    .A1(_04835_),
    .A2(_04554_),
    .A3(_04107_),
    .S0(_05979_),
    .S1(_05986_),
    .X(_06028_));
 sky130_fd_sc_hd__mux4_1 _12850_ (.A0(_04103_),
    .A1(_04711_),
    .A2(_04589_),
    .A3(_04586_),
    .S0(net28),
    .S1(_05986_),
    .X(_06029_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(_04110_),
    .A1(_04111_),
    .S(_05979_),
    .X(_06030_));
 sky130_fd_sc_hd__mux2_1 _12852_ (.A0(_06029_),
    .A1(_06030_),
    .S(_05982_),
    .X(_06031_));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(_06028_),
    .A1(_06031_),
    .S(_05987_),
    .X(_06032_));
 sky130_fd_sc_hd__and3_1 _12854_ (.A(net33),
    .B(_06027_),
    .C(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__a211o_2 _12855_ (.A1(_05989_),
    .A2(_06000_),
    .B1(_06026_),
    .C1(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__or4_1 _12856_ (.A(net32),
    .B(net33),
    .C(_05990_),
    .D(_05997_),
    .X(_06035_));
 sky130_fd_sc_hd__o22a_2 _12857_ (.A1(_05988_),
    .A2(_06034_),
    .B1(_06035_),
    .B2(_05647_),
    .X(_06036_));
 sky130_fd_sc_hd__mux2_2 _12858_ (.A0(\reg_gpout[4] ),
    .A1(clknet_1_0__leaf__06036_),
    .S(net45),
    .X(_06037_));
 sky130_fd_sc_hd__buf_1 _12859_ (.A(_06037_),
    .X(net61));
 sky130_fd_sc_hd__inv_2 _12860_ (.A(net37),
    .Y(_06038_));
 sky130_fd_sc_hd__buf_2 _12861_ (.A(net36),
    .X(_06039_));
 sky130_fd_sc_hd__buf_2 _12862_ (.A(net35),
    .X(_06040_));
 sky130_fd_sc_hd__inv_2 _12863_ (.A(net34),
    .Y(_06041_));
 sky130_fd_sc_hd__nor2_1 _12864_ (.A(net35),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__nor2_2 _12865_ (.A(net35),
    .B(net34),
    .Y(_06043_));
 sky130_fd_sc_hd__a22o_1 _12866_ (.A1(net54),
    .A2(_06042_),
    .B1(_06043_),
    .B2(net53),
    .X(_06044_));
 sky130_fd_sc_hd__a31o_1 _12867_ (.A1(net56),
    .A2(_06040_),
    .A3(_06041_),
    .B1(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__clkbuf_4 _12868_ (.A(net34),
    .X(_06046_));
 sky130_fd_sc_hd__and2_1 _12869_ (.A(_05772_),
    .B(net36),
    .X(_06047_));
 sky130_fd_sc_hd__nor2_1 _12870_ (.A(net37),
    .B(_06039_),
    .Y(_06048_));
 sky130_fd_sc_hd__a22o_1 _12871_ (.A1(_06038_),
    .A2(_06047_),
    .B1(_06048_),
    .B2(\gpout5.clk_div[1] ),
    .X(_06049_));
 sky130_fd_sc_hd__or2_1 _12872_ (.A(net37),
    .B(net36),
    .X(_06050_));
 sky130_fd_sc_hd__a211oi_2 _12873_ (.A1(net127),
    .A2(_06040_),
    .B1(_06046_),
    .C1(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__a31o_2 _12874_ (.A1(_06040_),
    .A2(_06046_),
    .A3(_06049_),
    .B1(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__a31o_2 _12875_ (.A1(_06038_),
    .A2(_06039_),
    .A3(_06045_),
    .B1(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__nor2_1 _12876_ (.A(net38),
    .B(net39),
    .Y(_06054_));
 sky130_fd_sc_hd__nor2_1 _12877_ (.A(_06038_),
    .B(net38),
    .Y(_06055_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(net41),
    .A1(net42),
    .S(_06046_),
    .X(_06056_));
 sky130_fd_sc_hd__and4b_1 _12879_ (.A_N(_06039_),
    .B(net39),
    .C(_06055_),
    .D(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__a22o_2 _12880_ (.A1(_06053_),
    .A2(_06054_),
    .B1(_06057_),
    .B2(_06040_),
    .X(_06058_));
 sky130_fd_sc_hd__inv_2 _12881_ (.A(net39),
    .Y(_06059_));
 sky130_fd_sc_hd__or2_1 _12882_ (.A(_06046_),
    .B(_05181_),
    .X(_06060_));
 sky130_fd_sc_hd__nand2_1 _12883_ (.A(_06046_),
    .B(_05409_),
    .Y(_06061_));
 sky130_fd_sc_hd__mux4_1 _12884_ (.A0(_05493_),
    .A1(_05573_),
    .A2(_05647_),
    .A3(_05725_),
    .S0(_06046_),
    .S1(net37),
    .X(_06062_));
 sky130_fd_sc_hd__a32o_1 _12885_ (.A1(_06060_),
    .A2(_06055_),
    .A3(_06061_),
    .B1(_06062_),
    .B2(net38),
    .X(_06063_));
 sky130_fd_sc_hd__mux2_1 _12886_ (.A0(_05744_),
    .A1(_05745_),
    .S(_06046_),
    .X(_06064_));
 sky130_fd_sc_hd__mux4_1 _12887_ (.A0(_04588_),
    .A1(_04835_),
    .A2(_04554_),
    .A3(_04107_),
    .S0(net34),
    .S1(net35),
    .X(_06065_));
 sky130_fd_sc_hd__a22o_1 _12888_ (.A1(_04111_),
    .A2(_06042_),
    .B1(_06043_),
    .B2(_04110_),
    .X(_06066_));
 sky130_fd_sc_hd__mux2_1 _12889_ (.A0(_06065_),
    .A1(_06066_),
    .S(_06039_),
    .X(_06067_));
 sky130_fd_sc_hd__a31oi_1 _12890_ (.A1(_06040_),
    .A2(_06039_),
    .A3(_06064_),
    .B1(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__mux2_1 _12891_ (.A0(_05177_),
    .A1(_05746_),
    .S(net34),
    .X(_06069_));
 sky130_fd_sc_hd__nand2_1 _12892_ (.A(_06039_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__nor2_1 _12893_ (.A(_04788_),
    .B(net34),
    .Y(_06071_));
 sky130_fd_sc_hd__a211o_1 _12894_ (.A1(_04817_),
    .A2(_06046_),
    .B1(_06039_),
    .C1(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__mux4_1 _12895_ (.A0(\gpout0.vpos[2] ),
    .A1(_04793_),
    .A2(_04782_),
    .A3(_04775_),
    .S0(net34),
    .S1(net36),
    .X(_06073_));
 sky130_fd_sc_hd__o21ai_1 _12896_ (.A1(_06040_),
    .A2(_06073_),
    .B1(net37),
    .Y(_06074_));
 sky130_fd_sc_hd__a31o_1 _12897_ (.A1(_06040_),
    .A2(_06070_),
    .A3(_06072_),
    .B1(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__o211a_1 _12898_ (.A1(net37),
    .A2(_06068_),
    .B1(_06075_),
    .C1(net38),
    .X(_06076_));
 sky130_fd_sc_hd__a31o_1 _12899_ (.A1(net44),
    .A2(net35),
    .A3(_06041_),
    .B1(_06050_),
    .X(_06077_));
 sky130_fd_sc_hd__a221o_1 _12900_ (.A1(net46),
    .A2(_06042_),
    .B1(_06043_),
    .B2(net43),
    .C1(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__a31o_1 _12901_ (.A1(_06040_),
    .A2(_06046_),
    .A3(_05200_),
    .B1(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__a221o_1 _12902_ (.A1(net40),
    .A2(_06042_),
    .B1(_06043_),
    .B2(net52),
    .C1(_06038_),
    .X(_06080_));
 sky130_fd_sc_hd__nand2_1 _12903_ (.A(net72),
    .B(_06042_),
    .Y(_06081_));
 sky130_fd_sc_hd__mux2_1 _12904_ (.A0(net50),
    .A1(net51),
    .S(net34),
    .X(_06082_));
 sky130_fd_sc_hd__nand2_1 _12905_ (.A(_06040_),
    .B(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__o311a_1 _12906_ (.A1(net35),
    .A2(_06046_),
    .A3(_05179_),
    .B1(_06081_),
    .C1(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__o21ai_1 _12907_ (.A1(net37),
    .A2(_06084_),
    .B1(_06039_),
    .Y(_06085_));
 sky130_fd_sc_hd__mux4_1 _12908_ (.A0(_04103_),
    .A1(_04711_),
    .A2(_04589_),
    .A3(_04586_),
    .S0(net34),
    .S1(net35),
    .X(_06086_));
 sky130_fd_sc_hd__a31o_1 _12909_ (.A1(net37),
    .A2(_06039_),
    .A3(_06086_),
    .B1(net38),
    .X(_06087_));
 sky130_fd_sc_hd__a31o_1 _12910_ (.A1(_06079_),
    .A2(_06080_),
    .A3(_06085_),
    .B1(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__and3b_1 _12911_ (.A_N(_06076_),
    .B(net39),
    .C(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__a41o_1 _12912_ (.A1(_06040_),
    .A2(_06039_),
    .A3(_06059_),
    .A4(_06063_),
    .B1(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__nand3_1 _12913_ (.A(_06043_),
    .B(_06048_),
    .C(_06054_),
    .Y(_06091_));
 sky130_fd_sc_hd__o22a_2 _12914_ (.A1(_06058_),
    .A2(_06090_),
    .B1(_06091_),
    .B2(_05725_),
    .X(_06092_));
 sky130_fd_sc_hd__mux2_2 _12915_ (.A0(\reg_gpout[5] ),
    .A1(clknet_1_1__leaf__06092_),
    .S(net45),
    .X(_06093_));
 sky130_fd_sc_hd__buf_1 _12916_ (.A(_06093_),
    .X(net62));
 sky130_fd_sc_hd__nor3b_4 _12917_ (.A(_04563_),
    .B(_04564_),
    .C_N(\rbzero.trace_state[3] ),
    .Y(_06094_));
 sky130_fd_sc_hd__buf_8 _12918_ (.A(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__and2b_1 _12919_ (.A_N(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .X(_06096_));
 sky130_fd_sc_hd__nand2_2 _12920_ (.A(\rbzero.trace_state[1] ),
    .B(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__nor2_1 _12921_ (.A(\rbzero.trace_state[0] ),
    .B(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__buf_6 _12922_ (.A(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__buf_6 _12923_ (.A(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__buf_6 _12924_ (.A(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__inv_2 _12925_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .Y(_06102_));
 sky130_fd_sc_hd__nor2_1 _12926_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__inv_2 _12927_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .Y(_06104_));
 sky130_fd_sc_hd__inv_2 _12928_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .Y(_06105_));
 sky130_fd_sc_hd__and2_1 _12929_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__inv_2 _12930_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .Y(_06107_));
 sky130_fd_sc_hd__inv_2 _12931_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .Y(_06108_));
 sky130_fd_sc_hd__a22o_1 _12932_ (.A1(\rbzero.wall_tracer.trackDistX[3] ),
    .A2(_06107_),
    .B1(\rbzero.wall_tracer.trackDistX[2] ),
    .B2(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__inv_2 _12933_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .Y(_06110_));
 sky130_fd_sc_hd__inv_2 _12934_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .Y(_06111_));
 sky130_fd_sc_hd__o22a_1 _12935_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(_06110_),
    .B1(\rbzero.wall_tracer.trackDistX[-1] ),
    .B2(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__inv_2 _12936_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .Y(_06113_));
 sky130_fd_sc_hd__o2bb2a_1 _12937_ (.A1_N(\rbzero.wall_tracer.trackDistX[-1] ),
    .A2_N(_06111_),
    .B1(_06113_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_06114_));
 sky130_fd_sc_hd__nand2_1 _12938_ (.A(_06112_),
    .B(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__a2bb2o_1 _12939_ (.A1_N(_06104_),
    .A2_N(\rbzero.wall_tracer.trackDistX[-3] ),
    .B1(_06113_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_06116_));
 sky130_fd_sc_hd__inv_2 _12940_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .Y(_06117_));
 sky130_fd_sc_hd__a22o_1 _12941_ (.A1(_06117_),
    .A2(\rbzero.wall_tracer.trackDistX[1] ),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_06110_),
    .X(_06118_));
 sky130_fd_sc_hd__o22a_1 _12942_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_06108_),
    .B1(_06117_),
    .B2(\rbzero.wall_tracer.trackDistX[1] ),
    .X(_06119_));
 sky130_fd_sc_hd__o221a_1 _12943_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(_06105_),
    .B1(\rbzero.wall_tracer.trackDistX[3] ),
    .B2(_06107_),
    .C1(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__or4b_1 _12944_ (.A(_06115_),
    .B(_06116_),
    .C(_06118_),
    .D_N(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__a2111o_1 _12945_ (.A1(_06104_),
    .A2(\rbzero.wall_tracer.trackDistX[-3] ),
    .B1(_06106_),
    .C1(_06109_),
    .D1(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__inv_2 _12946_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .Y(_06123_));
 sky130_fd_sc_hd__inv_2 _12947_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .Y(_06124_));
 sky130_fd_sc_hd__nor2_1 _12948_ (.A(_06124_),
    .B(\rbzero.wall_tracer.trackDistY[-6] ),
    .Y(_06125_));
 sky130_fd_sc_hd__inv_2 _12949_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .Y(_06126_));
 sky130_fd_sc_hd__nor2_1 _12950_ (.A(_06126_),
    .B(\rbzero.wall_tracer.trackDistY[9] ),
    .Y(_06127_));
 sky130_fd_sc_hd__a2111o_1 _12951_ (.A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .A2(_06123_),
    .B1(_06103_),
    .C1(_06125_),
    .D1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__inv_2 _12952_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .Y(_06129_));
 sky130_fd_sc_hd__inv_2 _12953_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .Y(_06130_));
 sky130_fd_sc_hd__a22o_1 _12954_ (.A1(_06129_),
    .A2(\rbzero.wall_tracer.trackDistY[-4] ),
    .B1(_06130_),
    .B2(\rbzero.wall_tracer.trackDistY[-5] ),
    .X(_06131_));
 sky130_fd_sc_hd__a221o_1 _12955_ (.A1(\rbzero.wall_tracer.trackDistY[10] ),
    .A2(_06102_),
    .B1(_06126_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .C1(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__inv_2 _12956_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .Y(_06133_));
 sky130_fd_sc_hd__nand2_1 _12957_ (.A(_06133_),
    .B(\rbzero.wall_tracer.trackDistY[-10] ),
    .Y(_06134_));
 sky130_fd_sc_hd__inv_2 _12958_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .Y(_06135_));
 sky130_fd_sc_hd__o22a_1 _12959_ (.A1(_06133_),
    .A2(\rbzero.wall_tracer.trackDistY[-10] ),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .B2(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__nand2_1 _12960_ (.A(_06134_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__inv_2 _12961_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .Y(_06138_));
 sky130_fd_sc_hd__nor2_1 _12962_ (.A(_06138_),
    .B(\rbzero.wall_tracer.trackDistY[-9] ),
    .Y(_06139_));
 sky130_fd_sc_hd__nor2_1 _12963_ (.A(_06129_),
    .B(\rbzero.wall_tracer.trackDistY[-4] ),
    .Y(_06140_));
 sky130_fd_sc_hd__a211o_1 _12964_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(_06135_),
    .B1(_06139_),
    .C1(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__or4_1 _12965_ (.A(_06128_),
    .B(_06132_),
    .C(_06137_),
    .D(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__inv_2 _12966_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .Y(_06143_));
 sky130_fd_sc_hd__inv_2 _12967_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .Y(_06144_));
 sky130_fd_sc_hd__a2bb2o_1 _12968_ (.A1_N(_06143_),
    .A2_N(\rbzero.wall_tracer.trackDistY[7] ),
    .B1(\rbzero.wall_tracer.trackDistX[6] ),
    .B2(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__inv_2 _12969_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .Y(_06146_));
 sky130_fd_sc_hd__inv_2 _12970_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .Y(_06147_));
 sky130_fd_sc_hd__or2_1 _12971_ (.A(_06147_),
    .B(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_06148_));
 sky130_fd_sc_hd__o21ai_1 _12972_ (.A1(\rbzero.wall_tracer.trackDistY[5] ),
    .A2(_06146_),
    .B1(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__a2bb2o_1 _12973_ (.A1_N(\rbzero.wall_tracer.trackDistX[6] ),
    .A2_N(_06144_),
    .B1(\rbzero.wall_tracer.trackDistY[5] ),
    .B2(_06146_),
    .X(_06150_));
 sky130_fd_sc_hd__a22o_1 _12974_ (.A1(_06147_),
    .A2(\rbzero.wall_tracer.trackDistY[8] ),
    .B1(_06143_),
    .B2(\rbzero.wall_tracer.trackDistY[7] ),
    .X(_06151_));
 sky130_fd_sc_hd__or4_2 _12975_ (.A(_06145_),
    .B(_06149_),
    .C(_06150_),
    .D(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__inv_2 _12976_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .Y(_06153_));
 sky130_fd_sc_hd__a22o_1 _12977_ (.A1(_06153_),
    .A2(\rbzero.wall_tracer.trackDistY[-8] ),
    .B1(_06138_),
    .B2(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(_06154_));
 sky130_fd_sc_hd__inv_2 _12978_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .Y(_06155_));
 sky130_fd_sc_hd__inv_2 _12979_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .Y(_06156_));
 sky130_fd_sc_hd__inv_2 _12980_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .Y(_06157_));
 sky130_fd_sc_hd__a22o_1 _12981_ (.A1(_06124_),
    .A2(\rbzero.wall_tracer.trackDistY[-6] ),
    .B1(\rbzero.wall_tracer.trackDistY[-7] ),
    .B2(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__a221o_1 _12982_ (.A1(_06155_),
    .A2(\rbzero.wall_tracer.trackDistX[-7] ),
    .B1(\rbzero.wall_tracer.trackDistX[-8] ),
    .B2(_06156_),
    .C1(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__or4_1 _12983_ (.A(_06142_),
    .B(_06152_),
    .C(_06154_),
    .D(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__a21oi_1 _12984_ (.A1(_06134_),
    .A2(_06137_),
    .B1(_06139_),
    .Y(_06161_));
 sky130_fd_sc_hd__nand2_1 _12985_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(_06156_),
    .Y(_06162_));
 sky130_fd_sc_hd__o221a_1 _12986_ (.A1(\rbzero.wall_tracer.trackDistY[-7] ),
    .A2(_06157_),
    .B1(_06154_),
    .B2(_06161_),
    .C1(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__inv_2 _12987_ (.A(_06125_),
    .Y(_06164_));
 sky130_fd_sc_hd__o221a_1 _12988_ (.A1(_06130_),
    .A2(\rbzero.wall_tracer.trackDistY[-5] ),
    .B1(_06158_),
    .B2(_06163_),
    .C1(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__nor2_1 _12989_ (.A(_06131_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__nand2_1 _12990_ (.A(_06114_),
    .B(_06116_),
    .Y(_06167_));
 sky130_fd_sc_hd__a21o_1 _12991_ (.A1(_06112_),
    .A2(_06167_),
    .B1(_06118_),
    .X(_06168_));
 sky130_fd_sc_hd__a21o_1 _12992_ (.A1(_06119_),
    .A2(_06168_),
    .B1(_06109_),
    .X(_06169_));
 sky130_fd_sc_hd__o221a_1 _12993_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(_06105_),
    .B1(\rbzero.wall_tracer.trackDistX[3] ),
    .B2(_06107_),
    .C1(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__o32a_1 _12994_ (.A1(_06122_),
    .A2(_06140_),
    .A3(_06166_),
    .B1(_06170_),
    .B2(_06106_),
    .X(_06171_));
 sky130_fd_sc_hd__and2b_1 _12995_ (.A_N(_06145_),
    .B(_06150_),
    .X(_06172_));
 sky130_fd_sc_hd__o21ai_1 _12996_ (.A1(_06151_),
    .A2(_06172_),
    .B1(_06148_),
    .Y(_06173_));
 sky130_fd_sc_hd__o21a_1 _12997_ (.A1(_06152_),
    .A2(_06171_),
    .B1(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__nor2_1 _12998_ (.A(_06127_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__a221o_1 _12999_ (.A1(\rbzero.wall_tracer.trackDistY[10] ),
    .A2(_06102_),
    .B1(_06126_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .C1(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__o21ai_1 _13000_ (.A1(_06122_),
    .A2(_06160_),
    .B1(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__nor2_2 _13001_ (.A(_06103_),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__or3b_1 _13002_ (.A(_04563_),
    .B(_04564_),
    .C_N(\rbzero.trace_state[3] ),
    .X(_06179_));
 sky130_fd_sc_hd__clkbuf_2 _13003_ (.A(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__clkbuf_4 _13004_ (.A(\rbzero.map_rom.f3 ),
    .X(_06181_));
 sky130_fd_sc_hd__inv_2 _13005_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .Y(_06182_));
 sky130_fd_sc_hd__clkinv_2 _13006_ (.A(_06181_),
    .Y(_06183_));
 sky130_fd_sc_hd__clkbuf_4 _13007_ (.A(\rbzero.map_rom.f2 ),
    .X(_06184_));
 sky130_fd_sc_hd__inv_2 _13008_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .Y(_06185_));
 sky130_fd_sc_hd__clkinv_2 _13009_ (.A(\rbzero.map_rom.i_col[4] ),
    .Y(_06186_));
 sky130_fd_sc_hd__clkinv_2 _13010_ (.A(\rbzero.map_rom.d6 ),
    .Y(_06187_));
 sky130_fd_sc_hd__o22a_1 _13011_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_06186_),
    .B1(_06187_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .X(_06188_));
 sky130_fd_sc_hd__o221a_1 _13012_ (.A1(_04804_),
    .A2(_06184_),
    .B1(\rbzero.wall_tracer.mapY[5] ),
    .B2(_06185_),
    .C1(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__inv_2 _13013_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .Y(_06190_));
 sky130_fd_sc_hd__o22a_1 _13014_ (.A1(_04803_),
    .A2(\rbzero.map_rom.i_row[4] ),
    .B1(_06190_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .X(_06191_));
 sky130_fd_sc_hd__inv_2 _13015_ (.A(\rbzero.map_rom.c6 ),
    .Y(_06192_));
 sky130_fd_sc_hd__inv_2 _13016_ (.A(\rbzero.map_rom.b6 ),
    .Y(_06193_));
 sky130_fd_sc_hd__clkinv_2 _13017_ (.A(\rbzero.map_rom.a6 ),
    .Y(_06194_));
 sky130_fd_sc_hd__clkinv_2 _13018_ (.A(\rbzero.map_rom.i_row[4] ),
    .Y(_06195_));
 sky130_fd_sc_hd__o22a_1 _13019_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_06194_),
    .B1(_06195_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .X(_06196_));
 sky130_fd_sc_hd__o221a_1 _13020_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_06192_),
    .B1(_06193_),
    .B2(\rbzero.debug_overlay.playerY[2] ),
    .C1(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__o2111a_1 _13021_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_06183_),
    .B1(_06189_),
    .C1(_06191_),
    .D1(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__o221a_1 _13022_ (.A1(_04801_),
    .A2(_06181_),
    .B1(\rbzero.map_rom.b6 ),
    .B2(_06182_),
    .C1(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__clkinv_2 _13023_ (.A(_06184_),
    .Y(_06200_));
 sky130_fd_sc_hd__o2bb2a_1 _13024_ (.A1_N(\rbzero.debug_overlay.playerX[4] ),
    .A2_N(_06186_),
    .B1(_06200_),
    .B2(\rbzero.debug_overlay.playerX[2] ),
    .X(_06201_));
 sky130_fd_sc_hd__or4_1 _13025_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(\rbzero.wall_tracer.mapY[9] ),
    .C(\rbzero.wall_tracer.mapY[8] ),
    .D(\rbzero.wall_tracer.mapY[10] ),
    .X(_06202_));
 sky130_fd_sc_hd__xor2_1 _13026_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(\rbzero.map_rom.f1 ),
    .X(_06203_));
 sky130_fd_sc_hd__inv_2 _13027_ (.A(\rbzero.map_rom.f4 ),
    .Y(_06204_));
 sky130_fd_sc_hd__a22o_1 _13028_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_06187_),
    .B1(_06194_),
    .B2(\rbzero.debug_overlay.playerY[3] ),
    .X(_06205_));
 sky130_fd_sc_hd__a221o_1 _13029_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_06204_),
    .B1(_06192_),
    .B2(\rbzero.debug_overlay.playerY[1] ),
    .C1(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__or4_1 _13030_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(\rbzero.wall_tracer.mapX[10] ),
    .C(_06203_),
    .D(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__inv_2 _13031_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .Y(_06208_));
 sky130_fd_sc_hd__a211oi_1 _13032_ (.A1(_06208_),
    .A2(\rbzero.wall_tracer.mapX[5] ),
    .B1(\rbzero.wall_tracer.mapX[7] ),
    .C1(\rbzero.wall_tracer.mapX[6] ),
    .Y(_06209_));
 sky130_fd_sc_hd__o221a_1 _13033_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_06204_),
    .B1(\rbzero.wall_tracer.mapX[5] ),
    .B2(_06208_),
    .C1(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__nor2_1 _13034_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(\rbzero.wall_tracer.mapY[7] ),
    .Y(_06211_));
 sky130_fd_sc_hd__and4bb_1 _13035_ (.A_N(_06202_),
    .B_N(_06207_),
    .C(_06210_),
    .D(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__and3_1 _13036_ (.A(_06199_),
    .B(_06201_),
    .C(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__or4_1 _13037_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(\rbzero.wall_tracer.visualWallDist[6] ),
    .C(\rbzero.wall_tracer.visualWallDist[5] ),
    .D(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_06214_));
 sky130_fd_sc_hd__or4_1 _13038_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(\rbzero.wall_tracer.visualWallDist[2] ),
    .C(\rbzero.wall_tracer.visualWallDist[1] ),
    .D(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_06215_));
 sky130_fd_sc_hd__or4_1 _13039_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(\rbzero.wall_tracer.visualWallDist[-2] ),
    .C(\rbzero.wall_tracer.visualWallDist[-3] ),
    .D(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__or4_1 _13040_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(\rbzero.wall_tracer.visualWallDist[8] ),
    .C(_06214_),
    .D(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__or3b_4 _13041_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_06213_),
    .C_N(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__a21oi_1 _13042_ (.A1(_04831_),
    .A2(_04830_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .Y(_06219_));
 sky130_fd_sc_hd__clkbuf_4 _13043_ (.A(\rbzero.map_rom.f4 ),
    .X(_06220_));
 sky130_fd_sc_hd__nand2_1 _13044_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__or2_1 _13045_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06220_),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_4 _13046_ (.A(\rbzero.map_rom.f1 ),
    .X(_06223_));
 sky130_fd_sc_hd__xnor2_1 _13047_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__o221ai_1 _13048_ (.A1(\rbzero.map_overlay.i_mapdx[1] ),
    .A2(_06183_),
    .B1(_06200_),
    .B2(\rbzero.map_overlay.i_mapdx[2] ),
    .C1(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__a221o_1 _13049_ (.A1(\rbzero.map_overlay.i_mapdx[1] ),
    .A2(_06183_),
    .B1(_06221_),
    .B2(_06222_),
    .C1(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__a221o_1 _13050_ (.A1(\rbzero.map_overlay.i_mapdx[2] ),
    .A2(_06200_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .B2(_04831_),
    .C1(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__nor3_2 _13051_ (.A(_06218_),
    .B(_06219_),
    .C(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__clkbuf_4 _13052_ (.A(\rbzero.map_rom.d6 ),
    .X(_06229_));
 sky130_fd_sc_hd__and3_1 _13053_ (.A(\rbzero.map_rom.b6 ),
    .B(\rbzero.map_rom.a6 ),
    .C(\rbzero.map_rom.i_row[4] ),
    .X(_06230_));
 sky130_fd_sc_hd__or4_1 _13054_ (.A(\rbzero.map_rom.c6 ),
    .B(\rbzero.map_rom.b6 ),
    .C(\rbzero.map_rom.a6 ),
    .D(\rbzero.map_rom.i_row[4] ),
    .X(_06231_));
 sky130_fd_sc_hd__nor2_1 _13055_ (.A(_06229_),
    .B(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__a31o_1 _13056_ (.A1(_06229_),
    .A2(\rbzero.map_rom.c6 ),
    .A3(_06230_),
    .B1(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__nand2_1 _13057_ (.A(_06184_),
    .B(\rbzero.map_rom.b6 ),
    .Y(_06234_));
 sky130_fd_sc_hd__xnor2_1 _13058_ (.A(_06229_),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06235_));
 sky130_fd_sc_hd__nor2_1 _13059_ (.A(_06220_),
    .B(\rbzero.map_rom.d6 ),
    .Y(_06236_));
 sky130_fd_sc_hd__a21oi_1 _13060_ (.A1(_06181_),
    .A2(_06235_),
    .B1(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__and4_1 _13061_ (.A(_06220_),
    .B(_06181_),
    .C(_06184_),
    .D(\rbzero.map_rom.i_col[4] ),
    .X(_06238_));
 sky130_fd_sc_hd__a2bb2o_1 _13062_ (.A1_N(_06234_),
    .A2_N(_06237_),
    .B1(_06238_),
    .B2(_06223_),
    .X(_06239_));
 sky130_fd_sc_hd__or4_1 _13063_ (.A(_06220_),
    .B(_06181_),
    .C(_06184_),
    .D(\rbzero.map_rom.i_col[4] ),
    .X(_06240_));
 sky130_fd_sc_hd__or2_1 _13064_ (.A(\rbzero.map_rom.f2 ),
    .B(\rbzero.map_rom.b6 ),
    .X(_06241_));
 sky130_fd_sc_hd__nand2_1 _13065_ (.A(_06181_),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06242_));
 sky130_fd_sc_hd__or2_1 _13066_ (.A(_06181_),
    .B(\rbzero.map_rom.c6 ),
    .X(_06243_));
 sky130_fd_sc_hd__and4_1 _13067_ (.A(_06241_),
    .B(_06234_),
    .C(_06242_),
    .D(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__or3b_1 _13068_ (.A(\rbzero.map_rom.a6 ),
    .B(_06236_),
    .C_N(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__a221o_1 _13069_ (.A1(_06220_),
    .A2(_06229_),
    .B1(_06240_),
    .B2(_06245_),
    .C1(_06223_),
    .X(_06246_));
 sky130_fd_sc_hd__or3_1 _13070_ (.A(_06220_),
    .B(_06229_),
    .C(_06241_),
    .X(_06247_));
 sky130_fd_sc_hd__or4bb_1 _13071_ (.A(_06233_),
    .B(_06239_),
    .C_N(_06246_),
    .D_N(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__inv_2 _13072_ (.A(_06223_),
    .Y(_06249_));
 sky130_fd_sc_hd__a22o_1 _13073_ (.A1(_06223_),
    .A2(\rbzero.map_rom.c6 ),
    .B1(_06193_),
    .B2(_06204_),
    .X(_06250_));
 sky130_fd_sc_hd__a221o_1 _13074_ (.A1(_06183_),
    .A2(_06187_),
    .B1(_06192_),
    .B2(_06249_),
    .C1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__xnor2_1 _13075_ (.A(_06184_),
    .B(\rbzero.map_rom.a6 ),
    .Y(_06252_));
 sky130_fd_sc_hd__a221o_1 _13076_ (.A1(_06181_),
    .A2(_06229_),
    .B1(\rbzero.map_rom.b6 ),
    .B2(_06220_),
    .C1(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__and4_1 _13077_ (.A(_06223_),
    .B(\rbzero.map_rom.c6 ),
    .C(\rbzero.map_rom.a6 ),
    .D(_06195_),
    .X(_06254_));
 sky130_fd_sc_hd__or4b_1 _13078_ (.A(_06181_),
    .B(\rbzero.map_rom.i_col[4] ),
    .C(_06247_),
    .D_N(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__o21ai_1 _13079_ (.A1(_06251_),
    .A2(_06253_),
    .B1(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__o21ba_1 _13080_ (.A1(_06248_),
    .A2(_06256_),
    .B1_N(_06218_),
    .X(_06257_));
 sky130_fd_sc_hd__or2_2 _13081_ (.A(_06228_),
    .B(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__nor2_1 _13082_ (.A(_06180_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__xor2_1 _13083_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(_06229_),
    .X(_06260_));
 sky130_fd_sc_hd__a221o_1 _13084_ (.A1(\rbzero.map_overlay.i_mapdy[1] ),
    .A2(_06192_),
    .B1(_06194_),
    .B2(\rbzero.map_overlay.i_mapdy[3] ),
    .C1(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__o2bb2a_1 _13085_ (.A1_N(\rbzero.map_overlay.i_mapdy[2] ),
    .A2_N(_06193_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_04820_),
    .X(_06262_));
 sky130_fd_sc_hd__o221a_1 _13086_ (.A1(\rbzero.map_overlay.i_mapdy[1] ),
    .A2(_06192_),
    .B1(_06193_),
    .B2(\rbzero.map_overlay.i_mapdy[2] ),
    .C1(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__o221a_1 _13087_ (.A1(\rbzero.map_overlay.i_mapdy[3] ),
    .A2(_06194_),
    .B1(_06195_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__or3b_2 _13088_ (.A(_06261_),
    .B(_06232_),
    .C_N(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__a22o_1 _13089_ (.A1(\rbzero.map_overlay.i_otherx[3] ),
    .A2(_06249_),
    .B1(_06186_),
    .B2(\rbzero.map_overlay.i_otherx[4] ),
    .X(_06266_));
 sky130_fd_sc_hd__xor2_1 _13090_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .B(\rbzero.map_rom.i_row[4] ),
    .X(_06267_));
 sky130_fd_sc_hd__xor2_1 _13091_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(\rbzero.map_rom.c6 ),
    .X(_06268_));
 sky130_fd_sc_hd__inv_2 _13092_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .Y(_06269_));
 sky130_fd_sc_hd__o22a_1 _13093_ (.A1(_06269_),
    .A2(_06184_),
    .B1(_06186_),
    .B2(\rbzero.map_overlay.i_otherx[4] ),
    .X(_06270_));
 sky130_fd_sc_hd__or4b_1 _13094_ (.A(_06266_),
    .B(_06267_),
    .C(_06268_),
    .D_N(_06270_),
    .X(_06271_));
 sky130_fd_sc_hd__o22ai_1 _13095_ (.A1(\rbzero.map_overlay.i_othery[0] ),
    .A2(_06187_),
    .B1(_06193_),
    .B2(\rbzero.map_overlay.i_othery[2] ),
    .Y(_06272_));
 sky130_fd_sc_hd__a221o_1 _13096_ (.A1(\rbzero.map_overlay.i_othery[0] ),
    .A2(_06187_),
    .B1(_06194_),
    .B2(\rbzero.map_overlay.i_othery[3] ),
    .C1(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__a2bb2o_1 _13097_ (.A1_N(\rbzero.map_overlay.i_othery[3] ),
    .A2_N(_06194_),
    .B1(_06269_),
    .B2(_06184_),
    .X(_06274_));
 sky130_fd_sc_hd__a221o_1 _13098_ (.A1(_04842_),
    .A2(_06181_),
    .B1(_06193_),
    .B2(\rbzero.map_overlay.i_othery[2] ),
    .C1(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__a2bb2o_1 _13099_ (.A1_N(\rbzero.map_overlay.i_otherx[0] ),
    .A2_N(_06204_),
    .B1(_06223_),
    .B2(_04839_),
    .X(_06276_));
 sky130_fd_sc_hd__a221o_1 _13100_ (.A1(\rbzero.map_overlay.i_otherx[0] ),
    .A2(_06204_),
    .B1(_06183_),
    .B2(\rbzero.map_overlay.i_otherx[1] ),
    .C1(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__or3_1 _13101_ (.A(_06273_),
    .B(_06275_),
    .C(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__or2_1 _13102_ (.A(_06271_),
    .B(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__a21oi_4 _13103_ (.A1(_06265_),
    .A2(_06279_),
    .B1(_06218_),
    .Y(_06280_));
 sky130_fd_sc_hd__nor2_1 _13104_ (.A(_06258_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nor2_1 _13105_ (.A(_06180_),
    .B(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__or2_2 _13106_ (.A(_04566_),
    .B(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__a21oi_2 _13107_ (.A1(_06178_),
    .A2(_06259_),
    .B1(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__o21ai_4 _13108_ (.A1(_06095_),
    .A2(_06101_),
    .B1(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__clkbuf_4 _13109_ (.A(_06285_),
    .X(_06286_));
 sky130_fd_sc_hd__buf_4 _13110_ (.A(_06180_),
    .X(_06287_));
 sky130_fd_sc_hd__buf_6 _13111_ (.A(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__nor2_2 _13112_ (.A(_06288_),
    .B(_06286_),
    .Y(_06289_));
 sky130_fd_sc_hd__nand2_1 _13113_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_06290_));
 sky130_fd_sc_hd__or2_1 _13114_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_06291_));
 sky130_fd_sc_hd__nand3_1 _13115_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .C(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_1 _13116_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_06293_));
 sky130_fd_sc_hd__or2_1 _13117_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_06294_));
 sky130_fd_sc_hd__nand2_1 _13118_ (.A(_06293_),
    .B(_06294_),
    .Y(_06295_));
 sky130_fd_sc_hd__nand2_1 _13119_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06296_));
 sky130_fd_sc_hd__or2_1 _13120_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_06297_));
 sky130_fd_sc_hd__nand2_1 _13121_ (.A(_06296_),
    .B(_06297_),
    .Y(_06298_));
 sky130_fd_sc_hd__nor2_1 _13122_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06299_));
 sky130_fd_sc_hd__and2_1 _13123_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_06300_));
 sky130_fd_sc_hd__nor2_1 _13124_ (.A(_06299_),
    .B(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__or3b_1 _13125_ (.A(_06295_),
    .B(_06298_),
    .C_N(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__or2_1 _13126_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06303_));
 sky130_fd_sc_hd__xor2_2 _13127_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06304_));
 sky130_fd_sc_hd__and2_1 _13128_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06305_));
 sky130_fd_sc_hd__a31o_1 _13129_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_06304_),
    .B1(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__and2_1 _13130_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06307_));
 sky130_fd_sc_hd__a221o_2 _13131_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_06303_),
    .B2(_06306_),
    .C1(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__or2_2 _13132_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_06309_));
 sky130_fd_sc_hd__nand2_1 _13133_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_06310_));
 sky130_fd_sc_hd__or2_1 _13134_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_06311_));
 sky130_fd_sc_hd__and2_1 _13135_ (.A(_06310_),
    .B(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__nand4b_2 _13136_ (.A_N(_06302_),
    .B(_06308_),
    .C(_06309_),
    .D(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__nor2_1 _13137_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_06314_));
 sky130_fd_sc_hd__nand2_1 _13138_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06315_));
 sky130_fd_sc_hd__a2111o_1 _13139_ (.A1(_06310_),
    .A2(_06315_),
    .B1(_06299_),
    .C1(_06298_),
    .D1(_06295_),
    .X(_06316_));
 sky130_fd_sc_hd__o211a_1 _13140_ (.A1(_06314_),
    .A2(_06296_),
    .B1(_06316_),
    .C1(_06293_),
    .X(_06317_));
 sky130_fd_sc_hd__nand2_1 _13141_ (.A(_06291_),
    .B(_06290_),
    .Y(_06318_));
 sky130_fd_sc_hd__nand2_1 _13142_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_06319_));
 sky130_fd_sc_hd__or2_1 _13143_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_06320_));
 sky130_fd_sc_hd__nand2_1 _13144_ (.A(_06319_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__a211o_1 _13145_ (.A1(_06313_),
    .A2(_06317_),
    .B1(_06318_),
    .C1(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__nor2_1 _13146_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06323_));
 sky130_fd_sc_hd__a31oi_1 _13147_ (.A1(_06290_),
    .A2(_06292_),
    .A3(_06322_),
    .B1(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__or2_1 _13148_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_06325_));
 sky130_fd_sc_hd__nand2_1 _13149_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06326_));
 sky130_fd_sc_hd__nand2_1 _13150_ (.A(_06325_),
    .B(_06326_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand2_1 _13151_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_06328_));
 sky130_fd_sc_hd__o21a_2 _13152_ (.A1(_06324_),
    .A2(_06327_),
    .B1(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__a41o_1 _13153_ (.A1(_06290_),
    .A2(_06292_),
    .A3(_06322_),
    .A4(_06326_),
    .B1(_06323_),
    .X(_06330_));
 sky130_fd_sc_hd__nand2_1 _13154_ (.A(_06325_),
    .B(_06328_),
    .Y(_06331_));
 sky130_fd_sc_hd__xor2_2 _13155_ (.A(_06330_),
    .B(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__and2b_1 _13156_ (.A_N(_06323_),
    .B(_06326_),
    .X(_06333_));
 sky130_fd_sc_hd__a31oi_1 _13157_ (.A1(_06290_),
    .A2(_06292_),
    .A3(_06322_),
    .B1(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__and4_1 _13158_ (.A(_06290_),
    .B(_06292_),
    .C(_06322_),
    .D(_06333_),
    .X(_06335_));
 sky130_fd_sc_hd__or2_1 _13159_ (.A(_06334_),
    .B(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__nand3_1 _13160_ (.A(_06309_),
    .B(_06308_),
    .C(_06312_),
    .Y(_06337_));
 sky130_fd_sc_hd__a311o_1 _13161_ (.A1(_06310_),
    .A2(_06337_),
    .A3(_06315_),
    .B1(_06299_),
    .C1(_06298_),
    .X(_06338_));
 sky130_fd_sc_hd__or2_1 _13162_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_06339_));
 sky130_fd_sc_hd__a32o_1 _13163_ (.A1(_06309_),
    .A2(_06308_),
    .A3(_06312_),
    .B1(\rbzero.wall_tracer.rayAddendY[3] ),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .X(_06340_));
 sky130_fd_sc_hd__a221o_1 _13164_ (.A1(_06296_),
    .A2(_06297_),
    .B1(_06339_),
    .B2(_06340_),
    .C1(_06300_),
    .X(_06341_));
 sky130_fd_sc_hd__and2_1 _13165_ (.A(_06338_),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__a21o_1 _13166_ (.A1(_06313_),
    .A2(_06317_),
    .B1(_06321_),
    .X(_06343_));
 sky130_fd_sc_hd__a21o_1 _13167_ (.A1(_06319_),
    .A2(_06343_),
    .B1(_06318_),
    .X(_06344_));
 sky130_fd_sc_hd__nand3_1 _13168_ (.A(_06319_),
    .B(_06343_),
    .C(_06318_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _13169_ (.A(_06344_),
    .B(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a21oi_1 _13170_ (.A1(_06313_),
    .A2(_06317_),
    .B1(_06321_),
    .Y(_06347_));
 sky130_fd_sc_hd__and3_1 _13171_ (.A(_06321_),
    .B(_06313_),
    .C(_06317_),
    .X(_06348_));
 sky130_fd_sc_hd__nor2_1 _13172_ (.A(_06347_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__xor2_1 _13173_ (.A(_06301_),
    .B(_06340_),
    .X(_06350_));
 sky130_fd_sc_hd__a21o_1 _13174_ (.A1(_06309_),
    .A2(_06308_),
    .B1(_06312_),
    .X(_06351_));
 sky130_fd_sc_hd__and2_1 _13175_ (.A(_06337_),
    .B(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__nand2_1 _13176_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_06353_));
 sky130_fd_sc_hd__nand2_1 _13177_ (.A(_06309_),
    .B(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__a21o_1 _13178_ (.A1(_06303_),
    .A2(_06306_),
    .B1(_06307_),
    .X(_06355_));
 sky130_fd_sc_hd__xnor2_2 _13179_ (.A(_06354_),
    .B(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__nand2_1 _13180_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_06357_));
 sky130_fd_sc_hd__xnor2_2 _13181_ (.A(_06357_),
    .B(_06304_),
    .Y(_06358_));
 sky130_fd_sc_hd__and2b_1 _13182_ (.A_N(_06307_),
    .B(_06303_),
    .X(_06359_));
 sky130_fd_sc_hd__xor2_2 _13183_ (.A(_06359_),
    .B(_06306_),
    .X(_06360_));
 sky130_fd_sc_hd__xor2_2 _13184_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_06361_));
 sky130_fd_sc_hd__or4_1 _13185_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C(_06360_),
    .D(_06361_),
    .X(_06362_));
 sky130_fd_sc_hd__or4_1 _13186_ (.A(_06352_),
    .B(_06356_),
    .C(_06358_),
    .D(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__nor3_1 _13187_ (.A(_06349_),
    .B(_06350_),
    .C(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__a21o_1 _13188_ (.A1(_06296_),
    .A2(_06338_),
    .B1(_06295_),
    .X(_06365_));
 sky130_fd_sc_hd__nand3_1 _13189_ (.A(_06295_),
    .B(_06296_),
    .C(_06338_),
    .Y(_06366_));
 sky130_fd_sc_hd__nand2_1 _13190_ (.A(_06365_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__and3_1 _13191_ (.A(_06346_),
    .B(_06364_),
    .C(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__or4b_2 _13192_ (.A(_06332_),
    .B(_06336_),
    .C(_06342_),
    .D_N(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__nand2_8 _13193_ (.A(_06329_),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__buf_4 _13194_ (.A(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__buf_2 _13195_ (.A(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__o21a_1 _13196_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(\rbzero.wall_tracer.mapY[5] ),
    .B1(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__xnor2_1 _13197_ (.A(_06190_),
    .B(_06371_),
    .Y(_06374_));
 sky130_fd_sc_hd__xnor2_1 _13198_ (.A(_06195_),
    .B(_06371_),
    .Y(_06375_));
 sky130_fd_sc_hd__or2_1 _13199_ (.A(\rbzero.map_rom.a6 ),
    .B(_06371_),
    .X(_06376_));
 sky130_fd_sc_hd__inv_2 _13200_ (.A(_06371_),
    .Y(_06377_));
 sky130_fd_sc_hd__xnor2_1 _13201_ (.A(_06192_),
    .B(_06371_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_1 _13202_ (.A(_06229_),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__o21ai_1 _13203_ (.A1(_06192_),
    .A2(_06377_),
    .B1(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__xnor2_1 _13204_ (.A(_06193_),
    .B(_06371_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _13205_ (.A(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__o21ai_1 _13206_ (.A1(_06193_),
    .A2(_06377_),
    .B1(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__nand2_1 _13207_ (.A(\rbzero.map_rom.a6 ),
    .B(_06371_),
    .Y(_06384_));
 sky130_fd_sc_hd__or2b_1 _13208_ (.A(_06383_),
    .B_N(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__and3_1 _13209_ (.A(_06375_),
    .B(_06376_),
    .C(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__and2_1 _13210_ (.A(_06374_),
    .B(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__xor2_1 _13211_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_06371_),
    .X(_06388_));
 sky130_fd_sc_hd__o21a_1 _13212_ (.A1(_06373_),
    .A2(_06387_),
    .B1(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nor3_1 _13213_ (.A(_06388_),
    .B(_06373_),
    .C(_06387_),
    .Y(_06390_));
 sky130_fd_sc_hd__nor2_1 _13214_ (.A(_06389_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__a22o_1 _13215_ (.A1(\rbzero.wall_tracer.mapY[6] ),
    .A2(_06286_),
    .B1(_06289_),
    .B2(_06391_),
    .X(_00386_));
 sky130_fd_sc_hd__xor2_1 _13216_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .B(_06371_),
    .X(_06392_));
 sky130_fd_sc_hd__a21o_1 _13217_ (.A1(\rbzero.wall_tracer.mapY[6] ),
    .A2(_06372_),
    .B1(_06389_),
    .X(_06393_));
 sky130_fd_sc_hd__xor2_1 _13218_ (.A(_06392_),
    .B(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__a22o_1 _13219_ (.A1(\rbzero.wall_tracer.mapY[7] ),
    .A2(_06286_),
    .B1(_06289_),
    .B2(_06394_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _13220_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06372_),
    .X(_06395_));
 sky130_fd_sc_hd__nor2_1 _13221_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06372_),
    .Y(_06396_));
 sky130_fd_sc_hd__nor2_1 _13222_ (.A(_06395_),
    .B(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__o41a_1 _13223_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(\rbzero.wall_tracer.mapY[5] ),
    .A3(\rbzero.wall_tracer.mapY[7] ),
    .A4(\rbzero.wall_tracer.mapY[6] ),
    .B1(_06372_),
    .X(_06398_));
 sky130_fd_sc_hd__a31o_1 _13224_ (.A1(_06388_),
    .A2(_06387_),
    .A3(_06392_),
    .B1(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__xor2_1 _13225_ (.A(_06397_),
    .B(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__a22o_1 _13226_ (.A1(\rbzero.wall_tracer.mapY[8] ),
    .A2(_06286_),
    .B1(_06289_),
    .B2(_06400_),
    .X(_00388_));
 sky130_fd_sc_hd__a21o_1 _13227_ (.A1(_06397_),
    .A2(_06399_),
    .B1(_06395_),
    .X(_06401_));
 sky130_fd_sc_hd__xnor2_1 _13228_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(_06372_),
    .Y(_06402_));
 sky130_fd_sc_hd__xnor2_1 _13229_ (.A(_06401_),
    .B(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__a22o_1 _13230_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06286_),
    .B1(_06289_),
    .B2(_06403_),
    .X(_00389_));
 sky130_fd_sc_hd__o21a_1 _13231_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06372_),
    .B1(_06401_),
    .X(_06404_));
 sky130_fd_sc_hd__a21oi_1 _13232_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06372_),
    .B1(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__xor2_1 _13233_ (.A(\rbzero.wall_tracer.mapY[10] ),
    .B(_06372_),
    .X(_06406_));
 sky130_fd_sc_hd__xnor2_1 _13234_ (.A(_06405_),
    .B(_06406_),
    .Y(_06407_));
 sky130_fd_sc_hd__a22o_1 _13235_ (.A1(\rbzero.wall_tracer.mapY[10] ),
    .A2(_06286_),
    .B1(_06289_),
    .B2(_06407_),
    .X(_00390_));
 sky130_fd_sc_hd__nand2_1 _13236_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_06408_));
 sky130_fd_sc_hd__or2_1 _13237_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_06409_));
 sky130_fd_sc_hd__or2_1 _13238_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_06410_));
 sky130_fd_sc_hd__and2_1 _13239_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_06411_));
 sky130_fd_sc_hd__nor2_1 _13240_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_06412_));
 sky130_fd_sc_hd__nor2_1 _13241_ (.A(_06411_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__and2_1 _13242_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06414_));
 sky130_fd_sc_hd__nor2_1 _13243_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_06415_));
 sky130_fd_sc_hd__nor2_1 _13244_ (.A(_06414_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__xor2_2 _13245_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06417_));
 sky130_fd_sc_hd__o21a_1 _13246_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_06414_),
    .X(_06418_));
 sky130_fd_sc_hd__a21o_1 _13247_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[6] ),
    .B1(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__a21o_1 _13248_ (.A1(_06416_),
    .A2(_06417_),
    .B1(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__xor2_2 _13249_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_06421_));
 sky130_fd_sc_hd__nor2_1 _13250_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06422_));
 sky130_fd_sc_hd__nor2_1 _13251_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06423_));
 sky130_fd_sc_hd__nand2_1 _13252_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_06424_));
 sky130_fd_sc_hd__nor2_1 _13253_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _13254_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06426_));
 sky130_fd_sc_hd__nand2_1 _13255_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06427_));
 sky130_fd_sc_hd__o211a_1 _13256_ (.A1(_06424_),
    .A2(_06425_),
    .B1(_06426_),
    .C1(_06427_),
    .X(_06428_));
 sky130_fd_sc_hd__nand2_1 _13257_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06429_));
 sky130_fd_sc_hd__o31ai_4 _13258_ (.A1(_06422_),
    .A2(_06423_),
    .A3(_06428_),
    .B1(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__and2_1 _13259_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_06431_));
 sky130_fd_sc_hd__nor2_1 _13260_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_06432_));
 sky130_fd_sc_hd__nor2_2 _13261_ (.A(_06431_),
    .B(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__o21a_1 _13262_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[4] ),
    .B1(_06431_),
    .X(_06434_));
 sky130_fd_sc_hd__a21o_1 _13263_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[4] ),
    .B1(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__a311o_1 _13264_ (.A1(_06421_),
    .A2(_06430_),
    .A3(_06433_),
    .B1(_06435_),
    .C1(_06419_),
    .X(_06436_));
 sky130_fd_sc_hd__nand2_1 _13265_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_06437_));
 sky130_fd_sc_hd__or2b_1 _13266_ (.A(_06411_),
    .B_N(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__a31o_1 _13267_ (.A1(_06413_),
    .A2(_06420_),
    .A3(_06436_),
    .B1(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__and2_1 _13268_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_06440_));
 sky130_fd_sc_hd__a31o_1 _13269_ (.A1(_06409_),
    .A2(_06410_),
    .A3(_06439_),
    .B1(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__nor2_1 _13270_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_06442_));
 sky130_fd_sc_hd__a21o_1 _13271_ (.A1(_06408_),
    .A2(_06441_),
    .B1(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__o211a_2 _13272_ (.A1(_06324_),
    .A2(_06327_),
    .B1(_04561_),
    .C1(_06328_),
    .X(_06444_));
 sky130_fd_sc_hd__nor2_1 _13273_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_04562_),
    .Y(_06445_));
 sky130_fd_sc_hd__inv_2 _13274_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06446_));
 sky130_fd_sc_hd__o21a_1 _13275_ (.A1(_06444_),
    .A2(_06445_),
    .B1(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__a21oi_1 _13276_ (.A1(_04578_),
    .A2(_06443_),
    .B1(_06447_),
    .Y(_06448_));
 sky130_fd_sc_hd__or2_2 _13277_ (.A(_04578_),
    .B(_06444_),
    .X(_06449_));
 sky130_fd_sc_hd__nor2_1 _13278_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_04562_),
    .Y(_06450_));
 sky130_fd_sc_hd__a211o_2 _13279_ (.A1(_06408_),
    .A2(_06441_),
    .B1(_06446_),
    .C1(_06442_),
    .X(_06451_));
 sky130_fd_sc_hd__o21a_2 _13280_ (.A1(_06449_),
    .A2(_06450_),
    .B1(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__and2b_1 _13281_ (.A_N(_06442_),
    .B(_06408_),
    .X(_06453_));
 sky130_fd_sc_hd__xnor2_1 _13282_ (.A(_06441_),
    .B(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__nand2_1 _13283_ (.A(_04578_),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__inv_2 _13284_ (.A(_04561_),
    .Y(_06456_));
 sky130_fd_sc_hd__buf_2 _13285_ (.A(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__a21o_1 _13286_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_06457_),
    .B1(_04578_),
    .X(_06458_));
 sky130_fd_sc_hd__a21o_1 _13287_ (.A1(_04562_),
    .A2(_06332_),
    .B1(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__or3_1 _13288_ (.A(_06457_),
    .B(_06334_),
    .C(_06335_),
    .X(_06460_));
 sky130_fd_sc_hd__clkinv_4 _13289_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .Y(_06461_));
 sky130_fd_sc_hd__a21oi_1 _13290_ (.A1(_06461_),
    .A2(_06457_),
    .B1(_04577_),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_1 _13291_ (.A(_06410_),
    .B(_06439_),
    .Y(_06463_));
 sky130_fd_sc_hd__nand2_1 _13292_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_06464_));
 sky130_fd_sc_hd__nand2_1 _13293_ (.A(_06409_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__xnor2_2 _13294_ (.A(_06463_),
    .B(_06465_),
    .Y(_06466_));
 sky130_fd_sc_hd__o2bb2a_1 _13295_ (.A1_N(_06460_),
    .A2_N(_06462_),
    .B1(_06446_),
    .B2(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__a21boi_2 _13296_ (.A1(_06455_),
    .A2(_06459_),
    .B1_N(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__nor2_1 _13297_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_04562_),
    .Y(_06469_));
 sky130_fd_sc_hd__o21a_2 _13298_ (.A1(_06449_),
    .A2(_06469_),
    .B1(_06451_),
    .X(_06470_));
 sky130_fd_sc_hd__a31o_1 _13299_ (.A1(_06421_),
    .A2(_06430_),
    .A3(_06433_),
    .B1(_06435_),
    .X(_06471_));
 sky130_fd_sc_hd__a21oi_1 _13300_ (.A1(_06416_),
    .A2(_06471_),
    .B1(_06414_),
    .Y(_06472_));
 sky130_fd_sc_hd__xnor2_2 _13301_ (.A(_06417_),
    .B(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__or2_1 _13302_ (.A(_06446_),
    .B(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__a21o_1 _13303_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_06457_),
    .B1(_04577_),
    .X(_06475_));
 sky130_fd_sc_hd__a31o_1 _13304_ (.A1(_04561_),
    .A2(_06365_),
    .A3(_06366_),
    .B1(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__xnor2_2 _13305_ (.A(_06416_),
    .B(_06471_),
    .Y(_06477_));
 sky130_fd_sc_hd__and3_1 _13306_ (.A(_04561_),
    .B(_06338_),
    .C(_06341_),
    .X(_06478_));
 sky130_fd_sc_hd__a21o_1 _13307_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_06457_),
    .B1(_04577_),
    .X(_06479_));
 sky130_fd_sc_hd__o2bb2a_2 _13308_ (.A1_N(_04577_),
    .A2_N(_06477_),
    .B1(_06478_),
    .B2(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__a21o_1 _13309_ (.A1(_06430_),
    .A2(_06433_),
    .B1(_06431_),
    .X(_06481_));
 sky130_fd_sc_hd__xnor2_2 _13310_ (.A(_06421_),
    .B(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__nand2_1 _13311_ (.A(_04577_),
    .B(_06482_),
    .Y(_06483_));
 sky130_fd_sc_hd__a21o_1 _13312_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_06457_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06484_));
 sky130_fd_sc_hd__a21o_1 _13313_ (.A1(_04561_),
    .A2(_06350_),
    .B1(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__xnor2_2 _13314_ (.A(_06430_),
    .B(_06433_),
    .Y(_06486_));
 sky130_fd_sc_hd__a21o_1 _13315_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_06457_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06487_));
 sky130_fd_sc_hd__and3_1 _13316_ (.A(_04561_),
    .B(_06337_),
    .C(_06351_),
    .X(_06488_));
 sky130_fd_sc_hd__o2bb2a_2 _13317_ (.A1_N(_04577_),
    .A2_N(_06486_),
    .B1(_06487_),
    .B2(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__or2b_1 _13318_ (.A(_06425_),
    .B_N(_06426_),
    .X(_06490_));
 sky130_fd_sc_hd__xor2_1 _13319_ (.A(_06424_),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__mux2_1 _13320_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_06358_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06492_));
 sky130_fd_sc_hd__mux2_4 _13321_ (.A0(_06491_),
    .A1(_06492_),
    .S(_06446_),
    .X(_06493_));
 sky130_fd_sc_hd__mux2_1 _13322_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06494_));
 sky130_fd_sc_hd__mux2_2 _13323_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_06494_),
    .S(_06446_),
    .X(_06495_));
 sky130_fd_sc_hd__mux2_1 _13324_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06496_));
 sky130_fd_sc_hd__mux2_2 _13325_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_06496_),
    .S(_06446_),
    .X(_06497_));
 sky130_fd_sc_hd__or2_1 _13326_ (.A(_06495_),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__mux2_1 _13327_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_06361_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06499_));
 sky130_fd_sc_hd__or2_1 _13328_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_06500_));
 sky130_fd_sc_hd__and3_1 _13329_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .B(_06424_),
    .C(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__a21o_2 _13330_ (.A1(_06446_),
    .A2(_06499_),
    .B1(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__nor2_1 _13331_ (.A(_06498_),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__and2b_1 _13332_ (.A_N(_06493_),
    .B(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__o21ai_1 _13333_ (.A1(_06424_),
    .A2(_06425_),
    .B1(_06426_),
    .Y(_06505_));
 sky130_fd_sc_hd__and2b_1 _13334_ (.A_N(_06423_),
    .B(_06427_),
    .X(_06506_));
 sky130_fd_sc_hd__xnor2_1 _13335_ (.A(_06505_),
    .B(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__nand2_1 _13336_ (.A(_04561_),
    .B(_06360_),
    .Y(_06508_));
 sky130_fd_sc_hd__a21oi_1 _13337_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_06456_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06509_));
 sky130_fd_sc_hd__a22o_2 _13338_ (.A1(\rbzero.wall_tracer.rcp_sel[0] ),
    .A2(_06507_),
    .B1(_06508_),
    .B2(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__nand2_1 _13339_ (.A(_06504_),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__nor2_1 _13340_ (.A(_06423_),
    .B(_06428_),
    .Y(_06512_));
 sky130_fd_sc_hd__or2b_1 _13341_ (.A(_06422_),
    .B_N(_06429_),
    .X(_06513_));
 sky130_fd_sc_hd__xnor2_1 _13342_ (.A(_06512_),
    .B(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__mux2_1 _13343_ (.A0(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A1(_06356_),
    .S(_04561_),
    .X(_06515_));
 sky130_fd_sc_hd__mux2_2 _13344_ (.A0(_06514_),
    .A1(_06515_),
    .S(_06446_),
    .X(_06516_));
 sky130_fd_sc_hd__a2111o_1 _13345_ (.A1(_06483_),
    .A2(_06485_),
    .B1(_06489_),
    .C1(_06511_),
    .D1(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__a211oi_2 _13346_ (.A1(_06474_),
    .A2(_06476_),
    .B1(_06480_),
    .C1(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_1 _13347_ (.A(_06410_),
    .B(_06437_),
    .Y(_06519_));
 sky130_fd_sc_hd__a31o_1 _13348_ (.A1(_06413_),
    .A2(_06420_),
    .A3(_06436_),
    .B1(_06411_),
    .X(_06520_));
 sky130_fd_sc_hd__xnor2_1 _13349_ (.A(_06519_),
    .B(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__or2_1 _13350_ (.A(_06446_),
    .B(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__a21o_1 _13351_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_06457_),
    .B1(_04577_),
    .X(_06523_));
 sky130_fd_sc_hd__a31o_1 _13352_ (.A1(_04561_),
    .A2(_06344_),
    .A3(_06345_),
    .B1(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__or3_1 _13353_ (.A(_06457_),
    .B(_06347_),
    .C(_06348_),
    .X(_06525_));
 sky130_fd_sc_hd__a21oi_1 _13354_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_06457_),
    .B1(_04577_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand2_1 _13355_ (.A(_06420_),
    .B(_06436_),
    .Y(_06527_));
 sky130_fd_sc_hd__xor2_2 _13356_ (.A(_06413_),
    .B(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__a22o_2 _13357_ (.A1(_06525_),
    .A2(_06526_),
    .B1(_06528_),
    .B2(_04577_),
    .X(_06529_));
 sky130_fd_sc_hd__a21boi_1 _13358_ (.A1(_06522_),
    .A2(_06524_),
    .B1_N(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__and2_1 _13359_ (.A(_06518_),
    .B(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__nand4_4 _13360_ (.A(_06452_),
    .B(_06468_),
    .C(_06470_),
    .D(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__nor2_1 _13361_ (.A(_04578_),
    .B(_06444_),
    .Y(_06533_));
 sky130_fd_sc_hd__o21a_1 _13362_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_04562_),
    .B1(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__nor2_1 _13363_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_04562_),
    .Y(_06535_));
 sky130_fd_sc_hd__nor2_1 _13364_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_04562_),
    .Y(_06536_));
 sky130_fd_sc_hd__o31a_2 _13365_ (.A1(_04578_),
    .A2(_06444_),
    .A3(_06536_),
    .B1(_06451_),
    .X(_06537_));
 sky130_fd_sc_hd__nor2_1 _13366_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_04562_),
    .Y(_06538_));
 sky130_fd_sc_hd__o31a_1 _13367_ (.A1(_04578_),
    .A2(_06444_),
    .A3(_06538_),
    .B1(_06451_),
    .X(_06539_));
 sky130_fd_sc_hd__o211ai_2 _13368_ (.A1(_06449_),
    .A2(_06535_),
    .B1(_06537_),
    .C1(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__nor2_1 _13369_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_04562_),
    .Y(_06541_));
 sky130_fd_sc_hd__o21ai_1 _13370_ (.A1(_06449_),
    .A2(_06541_),
    .B1(_06451_),
    .Y(_06542_));
 sky130_fd_sc_hd__buf_2 _13371_ (.A(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__o31a_1 _13372_ (.A1(_06532_),
    .A2(_06534_),
    .A3(_06540_),
    .B1(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__mux2_1 _13373_ (.A0(_06448_),
    .A1(_06447_),
    .S(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__or3_1 _13374_ (.A(_06532_),
    .B(_06534_),
    .C(_06540_),
    .X(_06546_));
 sky130_fd_sc_hd__and4bb_1 _13375_ (.A_N(_06541_),
    .B_N(_06546_),
    .C(_06445_),
    .D(_06533_),
    .X(_06547_));
 sky130_fd_sc_hd__o21ai_1 _13376_ (.A1(_06449_),
    .A2(_06535_),
    .B1(_06537_),
    .Y(_06548_));
 sky130_fd_sc_hd__o211ai_1 _13377_ (.A1(_06532_),
    .A2(_06548_),
    .B1(_06539_),
    .C1(_06543_),
    .Y(_06549_));
 sky130_fd_sc_hd__and2_1 _13378_ (.A(_06542_),
    .B(_06548_),
    .X(_06550_));
 sky130_fd_sc_hd__a211o_1 _13379_ (.A1(_06543_),
    .A2(_06532_),
    .B1(_06539_),
    .C1(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__a21oi_1 _13380_ (.A1(_06408_),
    .A2(_06441_),
    .B1(_06442_),
    .Y(_06552_));
 sky130_fd_sc_hd__a21oi_1 _13381_ (.A1(_04578_),
    .A2(_06552_),
    .B1(_06534_),
    .Y(_06553_));
 sky130_fd_sc_hd__o211ai_1 _13382_ (.A1(_06532_),
    .A2(_06540_),
    .B1(_06553_),
    .C1(_06543_),
    .Y(_06554_));
 sky130_fd_sc_hd__and2_1 _13383_ (.A(_06542_),
    .B(_06540_),
    .X(_06555_));
 sky130_fd_sc_hd__a211o_1 _13384_ (.A1(_06543_),
    .A2(_06532_),
    .B1(_06553_),
    .C1(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__and4_1 _13385_ (.A(_06549_),
    .B(_06551_),
    .C(_06554_),
    .D(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__or3b_1 _13386_ (.A(_06545_),
    .B(_06547_),
    .C_N(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__o21a_1 _13387_ (.A1(_06449_),
    .A2(_06535_),
    .B1(_06451_),
    .X(_06559_));
 sky130_fd_sc_hd__inv_2 _13388_ (.A(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__o21a_1 _13389_ (.A1(_06532_),
    .A2(_06560_),
    .B1(_06543_),
    .X(_06561_));
 sky130_fd_sc_hd__xnor2_2 _13390_ (.A(_06537_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__nand2_1 _13391_ (.A(_06543_),
    .B(_06532_),
    .Y(_06563_));
 sky130_fd_sc_hd__xnor2_2 _13392_ (.A(_06560_),
    .B(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__o31a_1 _13393_ (.A1(_04578_),
    .A2(_06444_),
    .A3(_06541_),
    .B1(_06451_),
    .X(_06565_));
 sky130_fd_sc_hd__clkbuf_4 _13394_ (.A(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__a31o_1 _13395_ (.A1(_06468_),
    .A2(_06470_),
    .A3(_06531_),
    .B1(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__xor2_4 _13396_ (.A(_06452_),
    .B(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__or3_1 _13397_ (.A(_06562_),
    .B(_06564_),
    .C(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__nor2_1 _13398_ (.A(_06558_),
    .B(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__nor2_1 _13399_ (.A(_06566_),
    .B(_06518_),
    .Y(_06571_));
 sky130_fd_sc_hd__xor2_1 _13400_ (.A(_06529_),
    .B(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__nand2_1 _13401_ (.A(_06455_),
    .B(_06459_),
    .Y(_06573_));
 sky130_fd_sc_hd__a31o_1 _13402_ (.A1(_06467_),
    .A2(_06518_),
    .A3(_06530_),
    .B1(_06565_),
    .X(_06574_));
 sky130_fd_sc_hd__xor2_2 _13403_ (.A(_06573_),
    .B(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__a21oi_1 _13404_ (.A1(_06518_),
    .A2(_06530_),
    .B1(_06566_),
    .Y(_06576_));
 sky130_fd_sc_hd__xnor2_2 _13405_ (.A(_06467_),
    .B(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__nand2_1 _13406_ (.A(_06522_),
    .B(_06524_),
    .Y(_06578_));
 sky130_fd_sc_hd__a21o_1 _13407_ (.A1(_06529_),
    .A2(_06518_),
    .B1(_06565_),
    .X(_06579_));
 sky130_fd_sc_hd__xnor2_1 _13408_ (.A(_06578_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__or3b_1 _13409_ (.A(_06575_),
    .B(_06577_),
    .C_N(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__a21oi_2 _13410_ (.A1(_06468_),
    .A2(_06531_),
    .B1(_06566_),
    .Y(_06582_));
 sky130_fd_sc_hd__xnor2_4 _13411_ (.A(_06470_),
    .B(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__nor2_2 _13412_ (.A(_06581_),
    .B(_06583_),
    .Y(_06584_));
 sky130_fd_sc_hd__and2_1 _13413_ (.A(_06572_),
    .B(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__nand2_1 _13414_ (.A(_06570_),
    .B(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__buf_4 _13415_ (.A(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__nand2_1 _13416_ (.A(_06474_),
    .B(_06476_),
    .Y(_06588_));
 sky130_fd_sc_hd__o21ba_1 _13417_ (.A1(_06480_),
    .A2(_06517_),
    .B1_N(_06566_),
    .X(_06589_));
 sky130_fd_sc_hd__xnor2_1 _13418_ (.A(_06588_),
    .B(_06589_),
    .Y(_06590_));
 sky130_fd_sc_hd__clkbuf_2 _13419_ (.A(_06590_),
    .X(_06591_));
 sky130_fd_sc_hd__nor2_1 _13420_ (.A(_06511_),
    .B(_06516_),
    .Y(_06592_));
 sky130_fd_sc_hd__or2_2 _13421_ (.A(_06566_),
    .B(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__xnor2_4 _13422_ (.A(_06489_),
    .B(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__nand2_2 _13423_ (.A(_06483_),
    .B(_06485_),
    .Y(_06595_));
 sky130_fd_sc_hd__inv_2 _13424_ (.A(_06489_),
    .Y(_06596_));
 sky130_fd_sc_hd__a21oi_2 _13425_ (.A1(_06596_),
    .A2(_06592_),
    .B1(_06566_),
    .Y(_06597_));
 sky130_fd_sc_hd__xnor2_4 _13426_ (.A(_06595_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__nor2b_1 _13427_ (.A(_06566_),
    .B_N(_06511_),
    .Y(_06599_));
 sky130_fd_sc_hd__xor2_2 _13428_ (.A(_06516_),
    .B(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__or3_1 _13429_ (.A(_06594_),
    .B(_06598_),
    .C(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__nand2_2 _13430_ (.A(_06543_),
    .B(_06517_),
    .Y(_06602_));
 sky130_fd_sc_hd__xor2_2 _13431_ (.A(_06480_),
    .B(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__or2_2 _13432_ (.A(_06504_),
    .B(_06566_),
    .X(_06604_));
 sky130_fd_sc_hd__xnor2_4 _13433_ (.A(_06510_),
    .B(_06604_),
    .Y(_06605_));
 sky130_fd_sc_hd__and3b_1 _13434_ (.A_N(_06601_),
    .B(_06603_),
    .C(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__nor2_1 _13435_ (.A(_06564_),
    .B(_06568_),
    .Y(_06607_));
 sky130_fd_sc_hd__nor4b_2 _13436_ (.A(_06545_),
    .B(_06562_),
    .C(_06547_),
    .D_N(_06557_),
    .Y(_06608_));
 sky130_fd_sc_hd__and3_1 _13437_ (.A(_06607_),
    .B(_06608_),
    .C(_06585_),
    .X(_06609_));
 sky130_fd_sc_hd__and3b_1 _13438_ (.A_N(_06591_),
    .B(_06606_),
    .C(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__nor2_2 _13439_ (.A(_06503_),
    .B(_06566_),
    .Y(_06611_));
 sky130_fd_sc_hd__xnor2_4 _13440_ (.A(_06493_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__and2_2 _13441_ (.A(_06498_),
    .B(_06543_),
    .X(_06613_));
 sky130_fd_sc_hd__xor2_4 _13442_ (.A(_06502_),
    .B(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__xnor2_1 _13443_ (.A(_06596_),
    .B(_06593_),
    .Y(_06615_));
 sky130_fd_sc_hd__nor2_1 _13444_ (.A(_06615_),
    .B(_06598_),
    .Y(_06616_));
 sky130_fd_sc_hd__and4b_1 _13445_ (.A_N(_06591_),
    .B(_06603_),
    .C(_06616_),
    .D(_06609_),
    .X(_06617_));
 sky130_fd_sc_hd__a31oi_4 _13446_ (.A1(_06610_),
    .A2(_06612_),
    .A3(_06614_),
    .B1(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__and3b_1 _13447_ (.A_N(_06591_),
    .B(_06603_),
    .C(_06609_),
    .X(_06619_));
 sky130_fd_sc_hd__nor2_1 _13448_ (.A(_06601_),
    .B(_06605_),
    .Y(_06620_));
 sky130_fd_sc_hd__nor2_1 _13449_ (.A(_06591_),
    .B(_06603_),
    .Y(_06621_));
 sky130_fd_sc_hd__and4_1 _13450_ (.A(_06607_),
    .B(_06608_),
    .C(_06585_),
    .D(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__and3_1 _13451_ (.A(_06607_),
    .B(_06608_),
    .C(_06583_),
    .X(_06623_));
 sky130_fd_sc_hd__inv_2 _13452_ (.A(_06575_),
    .Y(_06624_));
 sky130_fd_sc_hd__inv_2 _13453_ (.A(_06583_),
    .Y(_06625_));
 sky130_fd_sc_hd__xnor2_2 _13454_ (.A(_06529_),
    .B(_06571_),
    .Y(_06626_));
 sky130_fd_sc_hd__a32o_1 _13455_ (.A1(_06624_),
    .A2(_06577_),
    .A3(_06625_),
    .B1(_06584_),
    .B2(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__and3_1 _13456_ (.A(_06607_),
    .B(_06608_),
    .C(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__nand2_1 _13457_ (.A(_06549_),
    .B(_06551_),
    .Y(_06629_));
 sky130_fd_sc_hd__and2_1 _13458_ (.A(_06554_),
    .B(_06556_),
    .X(_06630_));
 sky130_fd_sc_hd__a221o_1 _13459_ (.A1(_06629_),
    .A2(_06630_),
    .B1(_06564_),
    .B2(_06608_),
    .C1(_06545_),
    .X(_06631_));
 sky130_fd_sc_hd__or4_2 _13460_ (.A(_06622_),
    .B(_06623_),
    .C(_06628_),
    .D(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__xnor2_1 _13461_ (.A(_06502_),
    .B(_06613_),
    .Y(_06633_));
 sky130_fd_sc_hd__nand2_1 _13462_ (.A(_06612_),
    .B(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__inv_2 _13463_ (.A(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(_06495_),
    .B(_06543_),
    .Y(_06636_));
 sky130_fd_sc_hd__xor2_2 _13465_ (.A(_06497_),
    .B(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__and3_1 _13466_ (.A(_06495_),
    .B(_06635_),
    .C(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__and4b_1 _13467_ (.A_N(_06591_),
    .B(_06606_),
    .C(_06638_),
    .D(_06609_),
    .X(_06639_));
 sky130_fd_sc_hd__clkbuf_4 _13468_ (.A(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__a211oi_4 _13469_ (.A1(_06619_),
    .A2(_06620_),
    .B1(_06632_),
    .C1(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_1 _13470_ (.A(_06618_),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__clkbuf_4 _13471_ (.A(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__clkbuf_4 _13472_ (.A(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__clkbuf_4 _13473_ (.A(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__buf_2 _13474_ (.A(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__and4b_1 _13475_ (.A_N(_06591_),
    .B(_06606_),
    .C(_06504_),
    .D(_06609_),
    .X(_06647_));
 sky130_fd_sc_hd__clkbuf_4 _13476_ (.A(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__xnor2_2 _13477_ (.A(_06480_),
    .B(_06602_),
    .Y(_06649_));
 sky130_fd_sc_hd__buf_4 _13478_ (.A(_06609_),
    .X(_06650_));
 sky130_fd_sc_hd__o31a_2 _13479_ (.A1(_06591_),
    .A2(_06649_),
    .A3(_06616_),
    .B1(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__xnor2_1 _13480_ (.A(_06497_),
    .B(_06636_),
    .Y(_06652_));
 sky130_fd_sc_hd__nor2_1 _13481_ (.A(_06626_),
    .B(_06590_),
    .Y(_06653_));
 sky130_fd_sc_hd__and4b_1 _13482_ (.A_N(_06601_),
    .B(_06603_),
    .C(_06605_),
    .D(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__and4_1 _13483_ (.A(_06584_),
    .B(_06635_),
    .C(_06652_),
    .D(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__and4_1 _13484_ (.A(_06584_),
    .B(_06598_),
    .C(_06603_),
    .D(_06653_),
    .X(_06656_));
 sky130_fd_sc_hd__inv_2 _13485_ (.A(_06558_),
    .Y(_06657_));
 sky130_fd_sc_hd__o41a_1 _13486_ (.A1(_06569_),
    .A2(_06583_),
    .A3(_06655_),
    .A4(_06656_),
    .B1(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__or4_1 _13487_ (.A(_06648_),
    .B(_06640_),
    .C(_06651_),
    .D(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__buf_2 _13488_ (.A(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__clkbuf_4 _13489_ (.A(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__a31o_4 _13490_ (.A1(_06610_),
    .A2(_06612_),
    .A3(_06614_),
    .B1(_06617_),
    .X(_06662_));
 sky130_fd_sc_hd__and3_1 _13491_ (.A(_06607_),
    .B(_06608_),
    .C(_06656_),
    .X(_06663_));
 sky130_fd_sc_hd__inv_2 _13492_ (.A(_06564_),
    .Y(_06664_));
 sky130_fd_sc_hd__xor2_2 _13493_ (.A(_06493_),
    .B(_06611_),
    .X(_06665_));
 sky130_fd_sc_hd__nor2_1 _13494_ (.A(_06577_),
    .B(_06580_),
    .Y(_06666_));
 sky130_fd_sc_hd__nor3b_1 _13495_ (.A(_06575_),
    .B(_06583_),
    .C_N(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__a311o_1 _13496_ (.A1(_06584_),
    .A2(_06665_),
    .A3(_06654_),
    .B1(_06667_),
    .C1(_06568_),
    .X(_06668_));
 sky130_fd_sc_hd__and3_1 _13497_ (.A(_06664_),
    .B(_06608_),
    .C(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__or3_1 _13498_ (.A(_06545_),
    .B(_06547_),
    .C(_06557_),
    .X(_06670_));
 sky130_fd_sc_hd__or3b_1 _13499_ (.A(_06663_),
    .B(_06669_),
    .C_N(_06670_),
    .X(_06671_));
 sky130_fd_sc_hd__nand3_2 _13500_ (.A(_06570_),
    .B(_06626_),
    .C(_06584_),
    .Y(_06672_));
 sky130_fd_sc_hd__or4b_4 _13501_ (.A(_06648_),
    .B(_06623_),
    .C(_06671_),
    .D_N(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__or2_1 _13502_ (.A(_06662_),
    .B(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__buf_2 _13503_ (.A(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__and3_1 _13504_ (.A(_06598_),
    .B(_06618_),
    .C(_06641_),
    .X(_06676_));
 sky130_fd_sc_hd__a21o_1 _13505_ (.A1(_06594_),
    .A2(_06644_),
    .B1(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__nor2_4 _13506_ (.A(_06662_),
    .B(_06673_),
    .Y(_06678_));
 sky130_fd_sc_hd__a21o_1 _13507_ (.A1(_06618_),
    .A2(_06641_),
    .B1(_06649_),
    .X(_06679_));
 sky130_fd_sc_hd__a211o_2 _13508_ (.A1(_06619_),
    .A2(_06620_),
    .B1(_06632_),
    .C1(_06640_),
    .X(_06680_));
 sky130_fd_sc_hd__or3_1 _13509_ (.A(_06591_),
    .B(_06662_),
    .C(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__and3_1 _13510_ (.A(_06678_),
    .B(_06679_),
    .C(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__a21o_1 _13511_ (.A1(_06675_),
    .A2(_06677_),
    .B1(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__nor4_4 _13512_ (.A(_06648_),
    .B(_06640_),
    .C(_06651_),
    .D(_06658_),
    .Y(_06684_));
 sky130_fd_sc_hd__nand2_2 _13513_ (.A(_06684_),
    .B(_06678_),
    .Y(_06685_));
 sky130_fd_sc_hd__inv_2 _13514_ (.A(_06605_),
    .Y(_06686_));
 sky130_fd_sc_hd__and3_1 _13515_ (.A(_06600_),
    .B(_06618_),
    .C(_06641_),
    .X(_06687_));
 sky130_fd_sc_hd__a21oi_1 _13516_ (.A1(_06686_),
    .A2(_06644_),
    .B1(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__mux2_1 _13517_ (.A0(_06665_),
    .A1(_06614_),
    .S(_06643_),
    .X(_06689_));
 sky130_fd_sc_hd__nor2_4 _13518_ (.A(_06660_),
    .B(_06678_),
    .Y(_06690_));
 sky130_fd_sc_hd__a2bb2o_1 _13519_ (.A1_N(_06685_),
    .A2_N(_06688_),
    .B1(_06689_),
    .B2(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__o21a_1 _13520_ (.A1(_06575_),
    .A2(_06666_),
    .B1(_06625_),
    .X(_06692_));
 sky130_fd_sc_hd__a211o_1 _13521_ (.A1(_06570_),
    .A2(_06692_),
    .B1(_06663_),
    .C1(_06628_),
    .X(_06693_));
 sky130_fd_sc_hd__or2_1 _13522_ (.A(_06651_),
    .B(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__nor2_1 _13523_ (.A(_06660_),
    .B(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__or3_4 _13524_ (.A(_06651_),
    .B(_06663_),
    .C(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__a211o_1 _13525_ (.A1(_06661_),
    .A2(_06683_),
    .B1(_06691_),
    .C1(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__and3_1 _13526_ (.A(_06580_),
    .B(_06618_),
    .C(_06641_),
    .X(_06698_));
 sky130_fd_sc_hd__a21oi_1 _13527_ (.A1(_06572_),
    .A2(_06644_),
    .B1(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(_06575_),
    .A1(_06577_),
    .S(_06643_),
    .X(_06700_));
 sky130_fd_sc_hd__clkbuf_4 _13529_ (.A(_06678_),
    .X(_06701_));
 sky130_fd_sc_hd__mux2_1 _13530_ (.A0(_06699_),
    .A1(_06700_),
    .S(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__o21a_1 _13531_ (.A1(_06661_),
    .A2(_06702_),
    .B1(_06587_),
    .X(_06703_));
 sky130_fd_sc_hd__a21o_4 _13532_ (.A1(_06673_),
    .A2(_06680_),
    .B1(_06662_),
    .X(_06704_));
 sky130_fd_sc_hd__xnor2_4 _13533_ (.A(_06684_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__xnor2_2 _13534_ (.A(_06684_),
    .B(_06694_),
    .Y(_06706_));
 sky130_fd_sc_hd__a21o_1 _13535_ (.A1(_06684_),
    .A2(_06704_),
    .B1(_06706_),
    .X(_06707_));
 sky130_fd_sc_hd__a21oi_2 _13536_ (.A1(_06672_),
    .A2(_06707_),
    .B1(_06587_),
    .Y(_06708_));
 sky130_fd_sc_hd__nand2_1 _13537_ (.A(_06705_),
    .B(_06708_),
    .Y(_06709_));
 sky130_fd_sc_hd__nand2_1 _13538_ (.A(_06495_),
    .B(_06644_),
    .Y(_06710_));
 sky130_fd_sc_hd__nor2_4 _13539_ (.A(_06662_),
    .B(_06680_),
    .Y(_06711_));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(_06633_),
    .A1(_06637_),
    .S(_06711_),
    .X(_06712_));
 sky130_fd_sc_hd__o21ba_1 _13541_ (.A1(_06673_),
    .A2(_06643_),
    .B1_N(_06704_),
    .X(_06713_));
 sky130_fd_sc_hd__o22a_1 _13542_ (.A1(_06675_),
    .A2(_06710_),
    .B1(_06712_),
    .B2(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__o2bb2a_4 _13543_ (.A1_N(_06697_),
    .A2_N(_06703_),
    .B1(_06709_),
    .B2(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__clkbuf_4 _13544_ (.A(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__mux4_1 _13545_ (.A0(_06605_),
    .A1(_06633_),
    .A2(_06637_),
    .A3(_06612_),
    .S0(_06701_),
    .S1(_06711_),
    .X(_06717_));
 sky130_fd_sc_hd__nor2_2 _13546_ (.A(_06587_),
    .B(_06705_),
    .Y(_06718_));
 sky130_fd_sc_hd__nand2_2 _13547_ (.A(_06672_),
    .B(_06707_),
    .Y(_06719_));
 sky130_fd_sc_hd__nor2_4 _13548_ (.A(_06587_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__nand2_2 _13549_ (.A(_06684_),
    .B(_06674_),
    .Y(_06721_));
 sky130_fd_sc_hd__or2_1 _13550_ (.A(_06721_),
    .B(_06710_),
    .X(_06722_));
 sky130_fd_sc_hd__a22o_1 _13551_ (.A1(_06717_),
    .A2(_06718_),
    .B1(_06720_),
    .B2(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__clkbuf_4 _13552_ (.A(_06713_),
    .X(_06724_));
 sky130_fd_sc_hd__a21o_1 _13553_ (.A1(_06594_),
    .A2(_06644_),
    .B1(_06687_),
    .X(_06725_));
 sky130_fd_sc_hd__o21bai_4 _13554_ (.A1(_06673_),
    .A2(_06644_),
    .B1_N(_06704_),
    .Y(_06726_));
 sky130_fd_sc_hd__o211a_1 _13555_ (.A1(_06598_),
    .A2(_06645_),
    .B1(_06726_),
    .C1(_06679_),
    .X(_06727_));
 sky130_fd_sc_hd__a211o_1 _13556_ (.A1(_06724_),
    .A2(_06725_),
    .B1(_06727_),
    .C1(_06709_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_4 _13557_ (.A(_06706_),
    .X(_06729_));
 sky130_fd_sc_hd__clkbuf_4 _13558_ (.A(_06684_),
    .X(_06730_));
 sky130_fd_sc_hd__clkbuf_4 _13559_ (.A(_06701_),
    .X(_06731_));
 sky130_fd_sc_hd__and3_1 _13560_ (.A(_06674_),
    .B(_06679_),
    .C(_06681_),
    .X(_06732_));
 sky130_fd_sc_hd__a21o_1 _13561_ (.A1(_06731_),
    .A2(_06699_),
    .B1(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__and3_1 _13562_ (.A(_06568_),
    .B(_06618_),
    .C(_06641_),
    .X(_06734_));
 sky130_fd_sc_hd__a211o_1 _13563_ (.A1(_06583_),
    .A2(_06644_),
    .B1(_06734_),
    .C1(_06675_),
    .X(_06735_));
 sky130_fd_sc_hd__o211a_1 _13564_ (.A1(_06701_),
    .A2(_06700_),
    .B1(_06735_),
    .C1(_06661_),
    .X(_06736_));
 sky130_fd_sc_hd__a21o_1 _13565_ (.A1(_06730_),
    .A2(_06733_),
    .B1(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__and2_1 _13566_ (.A(_06629_),
    .B(_06645_),
    .X(_06738_));
 sky130_fd_sc_hd__mux2_1 _13567_ (.A0(_06562_),
    .A1(_06564_),
    .S(_06645_),
    .X(_06739_));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(_06738_),
    .A1(_06739_),
    .S(_06675_),
    .X(_06740_));
 sky130_fd_sc_hd__a211o_1 _13569_ (.A1(_06729_),
    .A2(_06737_),
    .B1(_06740_),
    .C1(_06650_),
    .X(_06741_));
 sky130_fd_sc_hd__and3b_2 _13570_ (.A_N(_06723_),
    .B(_06728_),
    .C(_06741_),
    .X(_06742_));
 sky130_fd_sc_hd__inv_2 _13571_ (.A(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__a21o_2 _13572_ (.A1(_06672_),
    .A2(_06707_),
    .B1(_06586_),
    .X(_06744_));
 sky130_fd_sc_hd__xnor2_2 _13573_ (.A(_06660_),
    .B(_06704_),
    .Y(_06745_));
 sky130_fd_sc_hd__mux2_1 _13574_ (.A0(_06495_),
    .A1(_06652_),
    .S(_06642_),
    .X(_06746_));
 sky130_fd_sc_hd__or3b_1 _13575_ (.A(_06745_),
    .B(_06713_),
    .C_N(_06746_),
    .X(_06747_));
 sky130_fd_sc_hd__or2_1 _13576_ (.A(_06744_),
    .B(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__mux2_1 _13577_ (.A0(_06598_),
    .A1(_06649_),
    .S(_06711_),
    .X(_06749_));
 sky130_fd_sc_hd__a21o_1 _13578_ (.A1(_06618_),
    .A2(_06641_),
    .B1(_06600_),
    .X(_06750_));
 sky130_fd_sc_hd__or3_1 _13579_ (.A(_06594_),
    .B(_06662_),
    .C(_06680_),
    .X(_06751_));
 sky130_fd_sc_hd__a21o_1 _13580_ (.A1(_06750_),
    .A2(_06751_),
    .B1(_06701_),
    .X(_06752_));
 sky130_fd_sc_hd__o211ai_1 _13581_ (.A1(_06675_),
    .A2(_06749_),
    .B1(_06752_),
    .C1(_06661_),
    .Y(_06753_));
 sky130_fd_sc_hd__mux2_1 _13582_ (.A0(_06633_),
    .A1(_06637_),
    .S(_06643_),
    .X(_06754_));
 sky130_fd_sc_hd__mux2_1 _13583_ (.A0(_06605_),
    .A1(_06612_),
    .S(_06643_),
    .X(_06755_));
 sky130_fd_sc_hd__o221a_1 _13584_ (.A1(_06721_),
    .A2(_06754_),
    .B1(_06685_),
    .B2(_06755_),
    .C1(_06706_),
    .X(_06756_));
 sky130_fd_sc_hd__or3_1 _13585_ (.A(_06626_),
    .B(_06662_),
    .C(_06680_),
    .X(_06757_));
 sky130_fd_sc_hd__a21o_1 _13586_ (.A1(_06618_),
    .A2(_06641_),
    .B1(_06591_),
    .X(_06758_));
 sky130_fd_sc_hd__a21o_1 _13587_ (.A1(_06757_),
    .A2(_06758_),
    .B1(_06701_),
    .X(_06759_));
 sky130_fd_sc_hd__and3_1 _13588_ (.A(_06577_),
    .B(_06618_),
    .C(_06641_),
    .X(_06760_));
 sky130_fd_sc_hd__a21oi_1 _13589_ (.A1(_06618_),
    .A2(_06641_),
    .B1(_06580_),
    .Y(_06761_));
 sky130_fd_sc_hd__or3_1 _13590_ (.A(_06674_),
    .B(_06760_),
    .C(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__or2_1 _13591_ (.A(_06660_),
    .B(_06694_),
    .X(_06763_));
 sky130_fd_sc_hd__a21oi_1 _13592_ (.A1(_06759_),
    .A2(_06762_),
    .B1(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__a211o_1 _13593_ (.A1(_06753_),
    .A2(_06756_),
    .B1(_06764_),
    .C1(_06650_),
    .X(_06765_));
 sky130_fd_sc_hd__a211o_1 _13594_ (.A1(_06594_),
    .A2(_06644_),
    .B1(_06676_),
    .C1(_06675_),
    .X(_06766_));
 sky130_fd_sc_hd__a211o_1 _13595_ (.A1(_06686_),
    .A2(_06643_),
    .B1(_06687_),
    .C1(_06701_),
    .X(_06767_));
 sky130_fd_sc_hd__a21oi_1 _13596_ (.A1(_06766_),
    .A2(_06767_),
    .B1(_06684_),
    .Y(_06768_));
 sky130_fd_sc_hd__o211a_1 _13597_ (.A1(_06637_),
    .A2(_06644_),
    .B1(_06690_),
    .C1(_06710_),
    .X(_06769_));
 sky130_fd_sc_hd__nor2_1 _13598_ (.A(_06685_),
    .B(_06689_),
    .Y(_06770_));
 sky130_fd_sc_hd__o31a_1 _13599_ (.A1(_06768_),
    .A2(_06769_),
    .A3(_06770_),
    .B1(_06706_),
    .X(_06771_));
 sky130_fd_sc_hd__a211oi_2 _13600_ (.A1(_06730_),
    .A2(_06733_),
    .B1(_06736_),
    .C1(_06729_),
    .Y(_06772_));
 sky130_fd_sc_hd__a211o_1 _13601_ (.A1(_06748_),
    .A2(_06765_),
    .B1(_06771_),
    .C1(_06772_),
    .X(_06773_));
 sky130_fd_sc_hd__o32a_1 _13602_ (.A1(_06684_),
    .A2(_06731_),
    .A3(_06710_),
    .B1(_06717_),
    .B2(_06745_),
    .X(_06774_));
 sky130_fd_sc_hd__a31o_1 _13603_ (.A1(_06684_),
    .A2(_06766_),
    .A3(_06767_),
    .B1(_06696_),
    .X(_06775_));
 sky130_fd_sc_hd__a21oi_1 _13604_ (.A1(_06661_),
    .A2(_06733_),
    .B1(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__o21a_1 _13605_ (.A1(_06731_),
    .A2(_06700_),
    .B1(_06735_),
    .X(_06777_));
 sky130_fd_sc_hd__o21ai_1 _13606_ (.A1(_06763_),
    .A2(_06777_),
    .B1(_06587_),
    .Y(_06778_));
 sky130_fd_sc_hd__o22a_4 _13607_ (.A1(_06744_),
    .A2(_06774_),
    .B1(_06776_),
    .B2(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__clkbuf_4 _13608_ (.A(_06745_),
    .X(_06780_));
 sky130_fd_sc_hd__mux4_1 _13609_ (.A0(_06495_),
    .A1(_06665_),
    .A2(_06614_),
    .A3(_06652_),
    .S0(_06643_),
    .S1(_06678_),
    .X(_06781_));
 sky130_fd_sc_hd__nand2_1 _13610_ (.A(_06708_),
    .B(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__and3_1 _13611_ (.A(_06678_),
    .B(_06757_),
    .C(_06758_),
    .X(_06783_));
 sky130_fd_sc_hd__a21oi_1 _13612_ (.A1(_06675_),
    .A2(_06749_),
    .B1(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__nand2_1 _13613_ (.A(_06750_),
    .B(_06751_),
    .Y(_06785_));
 sky130_fd_sc_hd__o221a_1 _13614_ (.A1(_06785_),
    .A2(_06685_),
    .B1(_06755_),
    .B2(_06721_),
    .C1(_06706_),
    .X(_06786_));
 sky130_fd_sc_hd__o21a_1 _13615_ (.A1(_06684_),
    .A2(_06784_),
    .B1(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__mux2_1 _13616_ (.A0(_06624_),
    .A1(_06625_),
    .S(_06711_),
    .X(_06788_));
 sky130_fd_sc_hd__or3_1 _13617_ (.A(_06678_),
    .B(_06760_),
    .C(_06761_),
    .X(_06789_));
 sky130_fd_sc_hd__a21bo_1 _13618_ (.A1(_06701_),
    .A2(_06788_),
    .B1_N(_06789_),
    .X(_06790_));
 sky130_fd_sc_hd__a21o_1 _13619_ (.A1(_06695_),
    .A2(_06790_),
    .B1(_06650_),
    .X(_06791_));
 sky130_fd_sc_hd__o22a_4 _13620_ (.A1(_06780_),
    .A2(_06782_),
    .B1(_06787_),
    .B2(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__o21a_1 _13621_ (.A1(_06675_),
    .A2(_06749_),
    .B1(_06752_),
    .X(_06793_));
 sky130_fd_sc_hd__a31o_1 _13622_ (.A1(_06661_),
    .A2(_06759_),
    .A3(_06762_),
    .B1(_06696_),
    .X(_06794_));
 sky130_fd_sc_hd__a21oi_1 _13623_ (.A1(_06730_),
    .A2(_06793_),
    .B1(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__clkinv_2 _13624_ (.A(_06568_),
    .Y(_06796_));
 sky130_fd_sc_hd__mux2_1 _13625_ (.A0(_06664_),
    .A1(_06796_),
    .S(_06643_),
    .X(_06797_));
 sky130_fd_sc_hd__mux2_1 _13626_ (.A0(_06788_),
    .A1(_06797_),
    .S(_06701_),
    .X(_06798_));
 sky130_fd_sc_hd__a21o_1 _13627_ (.A1(_06695_),
    .A2(_06798_),
    .B1(_06650_),
    .X(_06799_));
 sky130_fd_sc_hd__nand2_1 _13628_ (.A(_06726_),
    .B(_06746_),
    .Y(_06800_));
 sky130_fd_sc_hd__xnor2_1 _13629_ (.A(_06516_),
    .B(_06599_),
    .Y(_06801_));
 sky130_fd_sc_hd__mux4_1 _13630_ (.A0(_06801_),
    .A1(_06612_),
    .A2(_06633_),
    .A3(_06605_),
    .S0(_06701_),
    .S1(_06711_),
    .X(_06802_));
 sky130_fd_sc_hd__mux2_1 _13631_ (.A0(_06800_),
    .A1(_06802_),
    .S(_06705_),
    .X(_06803_));
 sky130_fd_sc_hd__o22a_2 _13632_ (.A1(_06795_),
    .A2(_06799_),
    .B1(_06803_),
    .B2(_06744_),
    .X(_06804_));
 sky130_fd_sc_hd__a2111o_4 _13633_ (.A1(_06773_),
    .A2(_06715_),
    .B1(_06779_),
    .C1(_06792_),
    .D1(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__a211o_1 _13634_ (.A1(_06675_),
    .A2(_06677_),
    .B1(_06682_),
    .C1(_06661_),
    .X(_06806_));
 sky130_fd_sc_hd__o211a_1 _13635_ (.A1(_06730_),
    .A2(_06702_),
    .B1(_06806_),
    .C1(_06729_),
    .X(_06807_));
 sky130_fd_sc_hd__a21o_1 _13636_ (.A1(_06583_),
    .A2(_06645_),
    .B1(_06734_),
    .X(_06808_));
 sky130_fd_sc_hd__nand2_1 _13637_ (.A(_06690_),
    .B(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__or2b_1 _13638_ (.A(_06685_),
    .B_N(_06739_),
    .X(_06810_));
 sky130_fd_sc_hd__nand2_1 _13639_ (.A(_06726_),
    .B(_06725_),
    .Y(_06811_));
 sky130_fd_sc_hd__mux2_1 _13640_ (.A0(_06686_),
    .A1(_06665_),
    .S(_06711_),
    .X(_06812_));
 sky130_fd_sc_hd__a21oi_1 _13641_ (.A1(_06713_),
    .A2(_06812_),
    .B1(_06745_),
    .Y(_06813_));
 sky130_fd_sc_hd__a221o_1 _13642_ (.A1(_06745_),
    .A2(_06714_),
    .B1(_06811_),
    .B2(_06813_),
    .C1(_06744_),
    .X(_06814_));
 sky130_fd_sc_hd__and4b_1 _13643_ (.A_N(_06807_),
    .B(_06809_),
    .C(_06810_),
    .D(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__clkbuf_4 _13644_ (.A(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__nor2_1 _13645_ (.A(_06731_),
    .B(_06797_),
    .Y(_06817_));
 sky130_fd_sc_hd__mux2_1 _13646_ (.A0(_06629_),
    .A1(_06562_),
    .S(_06645_),
    .X(_06818_));
 sky130_fd_sc_hd__nand2_1 _13647_ (.A(_06731_),
    .B(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__mux4_1 _13648_ (.A0(_06594_),
    .A1(_06600_),
    .A2(_06686_),
    .A3(_06598_),
    .S0(_06643_),
    .S1(_06674_),
    .X(_06820_));
 sky130_fd_sc_hd__mux2_1 _13649_ (.A0(_06781_),
    .A1(_06820_),
    .S(_06705_),
    .X(_06821_));
 sky130_fd_sc_hd__mux2_1 _13650_ (.A0(_06784_),
    .A1(_06790_),
    .S(_06660_),
    .X(_06822_));
 sky130_fd_sc_hd__o2bb2a_1 _13651_ (.A1_N(_06708_),
    .A2_N(_06821_),
    .B1(_06822_),
    .B2(_06696_),
    .X(_06823_));
 sky130_fd_sc_hd__and3b_1 _13652_ (.A_N(_06817_),
    .B(_06819_),
    .C(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__buf_2 _13653_ (.A(_06824_),
    .X(_06825_));
 sky130_fd_sc_hd__a21o_1 _13654_ (.A1(_06805_),
    .A2(_06816_),
    .B1(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__or2_1 _13655_ (.A(_06743_),
    .B(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__clkbuf_4 _13656_ (.A(_06827_),
    .X(_06828_));
 sky130_fd_sc_hd__clkbuf_4 _13657_ (.A(_06711_),
    .X(_06829_));
 sky130_fd_sc_hd__mux4_1 _13658_ (.A0(_06591_),
    .A1(_06594_),
    .A2(_06598_),
    .A3(_06649_),
    .S0(_06829_),
    .S1(_06731_),
    .X(_06830_));
 sky130_fd_sc_hd__nand2_1 _13659_ (.A(_06705_),
    .B(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__clkbuf_4 _13660_ (.A(_06708_),
    .X(_06832_));
 sky130_fd_sc_hd__o211a_1 _13661_ (.A1(_06705_),
    .A2(_06802_),
    .B1(_06831_),
    .C1(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__nand4_1 _13662_ (.A(_06730_),
    .B(_06693_),
    .C(_06759_),
    .D(_06762_),
    .Y(_06834_));
 sky130_fd_sc_hd__buf_2 _13663_ (.A(_06675_),
    .X(_06835_));
 sky130_fd_sc_hd__nor2_1 _13664_ (.A(_06630_),
    .B(_06829_),
    .Y(_06836_));
 sky130_fd_sc_hd__a211oi_1 _13665_ (.A1(_06835_),
    .A2(_06818_),
    .B1(_06836_),
    .C1(_06650_),
    .Y(_06837_));
 sky130_fd_sc_hd__o211a_1 _13666_ (.A1(_06730_),
    .A2(_06798_),
    .B1(_06834_),
    .C1(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__a211oi_2 _13667_ (.A1(_06747_),
    .A2(_06720_),
    .B1(_06833_),
    .C1(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__clkbuf_4 _13668_ (.A(_06839_),
    .X(_06840_));
 sky130_fd_sc_hd__xnor2_4 _13669_ (.A(_06828_),
    .B(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__nor2_1 _13670_ (.A(_06716_),
    .B(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__nand2_2 _13671_ (.A(_06748_),
    .B(_06765_),
    .Y(_06843_));
 sky130_fd_sc_hd__clkbuf_4 _13672_ (.A(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__clkinv_4 _13673_ (.A(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__buf_6 _13674_ (.A(_06826_),
    .X(_06846_));
 sky130_fd_sc_hd__buf_4 _13675_ (.A(_06742_),
    .X(_06847_));
 sky130_fd_sc_hd__nand2_1 _13676_ (.A(_06847_),
    .B(_06840_),
    .Y(_06848_));
 sky130_fd_sc_hd__inv_2 _13677_ (.A(_06648_),
    .Y(_06849_));
 sky130_fd_sc_hd__o21ai_4 _13678_ (.A1(_06846_),
    .A2(_06848_),
    .B1(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__nor2_1 _13679_ (.A(_06845_),
    .B(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__nand2_1 _13680_ (.A(_06842_),
    .B(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__buf_2 _13681_ (.A(_06792_),
    .X(_06853_));
 sky130_fd_sc_hd__nor2_1 _13682_ (.A(_06853_),
    .B(_06850_),
    .Y(_06854_));
 sky130_fd_sc_hd__nand2_1 _13683_ (.A(_06842_),
    .B(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__nor2_1 _13684_ (.A(_06853_),
    .B(_06841_),
    .Y(_06856_));
 sky130_fd_sc_hd__o21bai_1 _13685_ (.A1(_06716_),
    .A2(_06850_),
    .B1_N(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__nand2_1 _13686_ (.A(_06855_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__xnor2_1 _13687_ (.A(_06852_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__xnor2_4 _13688_ (.A(_06847_),
    .B(_06846_),
    .Y(_06860_));
 sky130_fd_sc_hd__or2_1 _13689_ (.A(_06853_),
    .B(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__clkbuf_4 _13690_ (.A(_06804_),
    .X(_06862_));
 sky130_fd_sc_hd__xnor2_4 _13691_ (.A(_06805_),
    .B(_06816_),
    .Y(_06863_));
 sky130_fd_sc_hd__nor2_1 _13692_ (.A(_06862_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__nand3_4 _13693_ (.A(_06805_),
    .B(_06825_),
    .C(_06816_),
    .Y(_06865_));
 sky130_fd_sc_hd__a21oi_1 _13694_ (.A1(_06846_),
    .A2(_06865_),
    .B1(_06779_),
    .Y(_06866_));
 sky130_fd_sc_hd__xnor2_1 _13695_ (.A(_06864_),
    .B(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__xnor2_1 _13696_ (.A(_06861_),
    .B(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__buf_4 _13697_ (.A(_06773_),
    .X(_06869_));
 sky130_fd_sc_hd__a21oi_2 _13698_ (.A1(_06869_),
    .A2(_06715_),
    .B1(_06792_),
    .Y(_06870_));
 sky130_fd_sc_hd__xnor2_2 _13699_ (.A(_06779_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__and3_1 _13700_ (.A(_06869_),
    .B(_06715_),
    .C(_06792_),
    .X(_06872_));
 sky130_fd_sc_hd__nor2_2 _13701_ (.A(_06870_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__or4_1 _13702_ (.A(_06825_),
    .B(_06816_),
    .C(_06871_),
    .D(_06873_),
    .X(_06874_));
 sky130_fd_sc_hd__a211o_1 _13703_ (.A1(_06869_),
    .A2(_06715_),
    .B1(_06779_),
    .C1(_06792_),
    .X(_06875_));
 sky130_fd_sc_hd__nor2_2 _13704_ (.A(_06875_),
    .B(_06862_),
    .Y(_06876_));
 sky130_fd_sc_hd__clkbuf_4 _13705_ (.A(_06816_),
    .X(_06877_));
 sky130_fd_sc_hd__clkbuf_4 _13706_ (.A(_06825_),
    .X(_06878_));
 sky130_fd_sc_hd__o22ai_2 _13707_ (.A1(_06877_),
    .A2(_06871_),
    .B1(_06873_),
    .B2(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand3_1 _13708_ (.A(_06876_),
    .B(_06874_),
    .C(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__nand2_1 _13709_ (.A(_06874_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__and2b_1 _13710_ (.A_N(_06868_),
    .B(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__nor2_1 _13711_ (.A(_06792_),
    .B(_06863_),
    .Y(_06883_));
 sky130_fd_sc_hd__or2_1 _13712_ (.A(_06716_),
    .B(_06860_),
    .X(_06884_));
 sky130_fd_sc_hd__nor2_1 _13713_ (.A(_06779_),
    .B(_06863_),
    .Y(_06885_));
 sky130_fd_sc_hd__a21oi_2 _13714_ (.A1(_06846_),
    .A2(_06865_),
    .B1(_06792_),
    .Y(_06886_));
 sky130_fd_sc_hd__xnor2_1 _13715_ (.A(_06885_),
    .B(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__o2bb2a_1 _13716_ (.A1_N(_06866_),
    .A2_N(_06883_),
    .B1(_06884_),
    .B2(_06887_),
    .X(_06888_));
 sky130_fd_sc_hd__xnor2_1 _13717_ (.A(_06881_),
    .B(_06868_),
    .Y(_06889_));
 sky130_fd_sc_hd__and2b_1 _13718_ (.A_N(_06888_),
    .B(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__nor2_1 _13719_ (.A(_06882_),
    .B(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__or2_1 _13720_ (.A(_06771_),
    .B(_06772_),
    .X(_06892_));
 sky130_fd_sc_hd__clkbuf_4 _13721_ (.A(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__buf_2 _13722_ (.A(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__or2_1 _13723_ (.A(_06894_),
    .B(_06841_),
    .X(_06895_));
 sky130_fd_sc_hd__or3_2 _13724_ (.A(_06845_),
    .B(_06850_),
    .C(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__xnor2_1 _13725_ (.A(_06842_),
    .B(_06851_),
    .Y(_06897_));
 sky130_fd_sc_hd__or2_1 _13726_ (.A(_06896_),
    .B(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__xnor2_1 _13727_ (.A(_06859_),
    .B(_06891_),
    .Y(_06899_));
 sky130_fd_sc_hd__or2_1 _13728_ (.A(_06898_),
    .B(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__o21ai_2 _13729_ (.A1(_06859_),
    .A2(_06891_),
    .B1(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__xnor2_4 _13730_ (.A(_06843_),
    .B(_06893_),
    .Y(_06902_));
 sky130_fd_sc_hd__nor2_1 _13731_ (.A(_06648_),
    .B(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__xor2_2 _13732_ (.A(_06869_),
    .B(_06715_),
    .X(_06904_));
 sky130_fd_sc_hd__and2_1 _13733_ (.A(_06840_),
    .B(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__xnor2_1 _13734_ (.A(_06903_),
    .B(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__and2_1 _13735_ (.A(_06742_),
    .B(_06904_),
    .X(_06907_));
 sky130_fd_sc_hd__nor2_2 _13736_ (.A(_06771_),
    .B(_06772_),
    .Y(_06908_));
 sky130_fd_sc_hd__mux2_1 _13737_ (.A0(_06908_),
    .A1(_06845_),
    .S(_06840_),
    .X(_06909_));
 sky130_fd_sc_hd__nand2_1 _13738_ (.A(_06908_),
    .B(_06839_),
    .Y(_06910_));
 sky130_fd_sc_hd__nor2_1 _13739_ (.A(_06845_),
    .B(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__a21oi_1 _13740_ (.A1(_06907_),
    .A2(_06909_),
    .B1(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__xnor2_1 _13741_ (.A(_06906_),
    .B(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__nand2_1 _13742_ (.A(_06875_),
    .B(_06804_),
    .Y(_06914_));
 sky130_fd_sc_hd__and2_1 _13743_ (.A(_06805_),
    .B(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__clkbuf_4 _13744_ (.A(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__nor2_1 _13745_ (.A(_06916_),
    .B(_06877_),
    .Y(_06917_));
 sky130_fd_sc_hd__nor2_1 _13746_ (.A(_06878_),
    .B(_06871_),
    .Y(_06918_));
 sky130_fd_sc_hd__or2_4 _13747_ (.A(_06870_),
    .B(_06872_),
    .X(_06919_));
 sky130_fd_sc_hd__nand2_1 _13748_ (.A(_06847_),
    .B(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__xnor2_1 _13749_ (.A(_06918_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__xnor2_1 _13750_ (.A(_06917_),
    .B(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__xor2_1 _13751_ (.A(_06913_),
    .B(_06922_),
    .X(_06923_));
 sky130_fd_sc_hd__xnor2_1 _13752_ (.A(_06907_),
    .B(_06909_),
    .Y(_06924_));
 sky130_fd_sc_hd__xnor2_4 _13753_ (.A(_06869_),
    .B(_06715_),
    .Y(_06925_));
 sky130_fd_sc_hd__or2_1 _13754_ (.A(_06825_),
    .B(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__xnor2_1 _13755_ (.A(_06844_),
    .B(_06908_),
    .Y(_06927_));
 sky130_fd_sc_hd__a21boi_1 _13756_ (.A1(_06847_),
    .A2(_06927_),
    .B1_N(_06910_),
    .Y(_06928_));
 sky130_fd_sc_hd__o2bb2a_1 _13757_ (.A1_N(_06847_),
    .A2_N(_06911_),
    .B1(_06926_),
    .B2(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__xnor2_1 _13758_ (.A(_06924_),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__inv_2 _13759_ (.A(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__a21o_1 _13760_ (.A1(_06874_),
    .A2(_06879_),
    .B1(_06876_),
    .X(_06932_));
 sky130_fd_sc_hd__and2_1 _13761_ (.A(_06880_),
    .B(_06932_),
    .X(_06933_));
 sky130_fd_sc_hd__nor2_1 _13762_ (.A(_06924_),
    .B(_06929_),
    .Y(_06934_));
 sky130_fd_sc_hd__a21oi_1 _13763_ (.A1(_06931_),
    .A2(_06933_),
    .B1(_06934_),
    .Y(_06935_));
 sky130_fd_sc_hd__xnor2_1 _13764_ (.A(_06923_),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__xnor2_1 _13765_ (.A(_06888_),
    .B(_06889_),
    .Y(_06937_));
 sky130_fd_sc_hd__or2b_1 _13766_ (.A(_06935_),
    .B_N(_06923_),
    .X(_06938_));
 sky130_fd_sc_hd__a21bo_1 _13767_ (.A1(_06936_),
    .A2(_06937_),
    .B1_N(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__nand2_1 _13768_ (.A(_06903_),
    .B(_06905_),
    .Y(_06940_));
 sky130_fd_sc_hd__nand2_1 _13769_ (.A(_06904_),
    .B(_06940_),
    .Y(_06941_));
 sky130_fd_sc_hd__nor2_1 _13770_ (.A(_06916_),
    .B(_06878_),
    .Y(_06942_));
 sky130_fd_sc_hd__clkbuf_4 _13771_ (.A(_06871_),
    .X(_06943_));
 sky130_fd_sc_hd__nor2_1 _13772_ (.A(_06743_),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2_1 _13773_ (.A(_06840_),
    .B(_06919_),
    .Y(_06945_));
 sky130_fd_sc_hd__xnor2_1 _13774_ (.A(_06944_),
    .B(_06945_),
    .Y(_06946_));
 sky130_fd_sc_hd__xnor2_1 _13775_ (.A(_06942_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__xor2_1 _13776_ (.A(_06941_),
    .B(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__or2_1 _13777_ (.A(_06906_),
    .B(_06912_),
    .X(_06949_));
 sky130_fd_sc_hd__o21ai_1 _13778_ (.A1(_06913_),
    .A2(_06922_),
    .B1(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__and2_1 _13779_ (.A(_06948_),
    .B(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__nor2_1 _13780_ (.A(_06948_),
    .B(_06950_),
    .Y(_06952_));
 sky130_fd_sc_hd__or2_1 _13781_ (.A(_06951_),
    .B(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__and2_2 _13782_ (.A(_06846_),
    .B(_06865_),
    .X(_06954_));
 sky130_fd_sc_hd__nor2_1 _13783_ (.A(_06862_),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__o2bb2ai_1 _13784_ (.A1_N(_06955_),
    .A2_N(_06885_),
    .B1(_06867_),
    .B2(_06861_),
    .Y(_06956_));
 sky130_fd_sc_hd__nor2_1 _13785_ (.A(_06743_),
    .B(_06873_),
    .Y(_06957_));
 sky130_fd_sc_hd__a22oi_2 _13786_ (.A1(_06918_),
    .A2(_06957_),
    .B1(_06921_),
    .B2(_06917_),
    .Y(_06958_));
 sky130_fd_sc_hd__buf_2 _13787_ (.A(_06779_),
    .X(_06959_));
 sky130_fd_sc_hd__nor2_1 _13788_ (.A(_06959_),
    .B(_06860_),
    .Y(_06960_));
 sky130_fd_sc_hd__nor2_1 _13789_ (.A(_06876_),
    .B(_06877_),
    .Y(_06961_));
 sky130_fd_sc_hd__xnor2_1 _13790_ (.A(_06955_),
    .B(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__xnor2_1 _13791_ (.A(_06960_),
    .B(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__xnor2_1 _13792_ (.A(_06958_),
    .B(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__xnor2_1 _13793_ (.A(_06956_),
    .B(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__xnor2_1 _13794_ (.A(_06953_),
    .B(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__xor2_1 _13795_ (.A(_06939_),
    .B(_06966_),
    .X(_06967_));
 sky130_fd_sc_hd__xnor2_1 _13796_ (.A(_06898_),
    .B(_06899_),
    .Y(_06968_));
 sky130_fd_sc_hd__and2b_1 _13797_ (.A_N(_06966_),
    .B(_06939_),
    .X(_06969_));
 sky130_fd_sc_hd__o21ba_1 _13798_ (.A1(_06967_),
    .A2(_06968_),
    .B1_N(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__nor2_1 _13799_ (.A(_06953_),
    .B(_06965_),
    .Y(_06971_));
 sky130_fd_sc_hd__nand2b_1 _13800_ (.A_N(_06943_),
    .B(_06840_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand2_1 _13801_ (.A(_06849_),
    .B(_06919_),
    .Y(_06973_));
 sky130_fd_sc_hd__xnor2_1 _13802_ (.A(_06972_),
    .B(_06973_),
    .Y(_06974_));
 sky130_fd_sc_hd__nand2_2 _13803_ (.A(_06805_),
    .B(_06914_),
    .Y(_06975_));
 sky130_fd_sc_hd__nand2_1 _13804_ (.A(_06975_),
    .B(_06847_),
    .Y(_06976_));
 sky130_fd_sc_hd__xnor2_1 _13805_ (.A(_06974_),
    .B(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__o21ai_1 _13806_ (.A1(_06925_),
    .A2(_06947_),
    .B1(_06940_),
    .Y(_06978_));
 sky130_fd_sc_hd__or2b_1 _13807_ (.A(_06977_),
    .B_N(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__or2b_1 _13808_ (.A(_06978_),
    .B_N(_06977_),
    .X(_06980_));
 sky130_fd_sc_hd__nand2_1 _13809_ (.A(_06979_),
    .B(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__or3_1 _13810_ (.A(_06959_),
    .B(_06860_),
    .C(_06962_),
    .X(_06982_));
 sky130_fd_sc_hd__a21bo_1 _13811_ (.A1(_06955_),
    .A2(_06961_),
    .B1_N(_06982_),
    .X(_06983_));
 sky130_fd_sc_hd__or2_1 _13812_ (.A(_06920_),
    .B(_06972_),
    .X(_06984_));
 sky130_fd_sc_hd__nand2_1 _13813_ (.A(_06942_),
    .B(_06946_),
    .Y(_06985_));
 sky130_fd_sc_hd__nor2_1 _13814_ (.A(_06805_),
    .B(_06878_),
    .Y(_06986_));
 sky130_fd_sc_hd__or2_1 _13815_ (.A(_06862_),
    .B(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__o2bb2a_1 _13816_ (.A1_N(_06743_),
    .A2_N(_06986_),
    .B1(_06987_),
    .B2(_06860_),
    .X(_06988_));
 sky130_fd_sc_hd__a21oi_1 _13817_ (.A1(_06984_),
    .A2(_06985_),
    .B1(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__and3_1 _13818_ (.A(_06984_),
    .B(_06985_),
    .C(_06988_),
    .X(_06990_));
 sky130_fd_sc_hd__or2_1 _13819_ (.A(_06989_),
    .B(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__xnor2_1 _13820_ (.A(_06983_),
    .B(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__xnor2_1 _13821_ (.A(_06981_),
    .B(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__o21ai_1 _13822_ (.A1(_06951_),
    .A2(_06971_),
    .B1(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__or3_1 _13823_ (.A(_06951_),
    .B(_06971_),
    .C(_06993_),
    .X(_06995_));
 sky130_fd_sc_hd__nand2_1 _13824_ (.A(_06994_),
    .B(_06995_),
    .Y(_06996_));
 sky130_fd_sc_hd__or2_1 _13825_ (.A(_06852_),
    .B(_06858_),
    .X(_06997_));
 sky130_fd_sc_hd__and2b_1 _13826_ (.A_N(_06958_),
    .B(_06963_),
    .X(_06998_));
 sky130_fd_sc_hd__a21o_1 _13827_ (.A1(_06956_),
    .A2(_06964_),
    .B1(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__nor2_1 _13828_ (.A(_06959_),
    .B(_06841_),
    .Y(_07000_));
 sky130_fd_sc_hd__xor2_1 _13829_ (.A(_06854_),
    .B(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__xnor2_1 _13830_ (.A(_06855_),
    .B(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__xnor2_1 _13831_ (.A(_06999_),
    .B(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__nor2_1 _13832_ (.A(_06997_),
    .B(_07003_),
    .Y(_07004_));
 sky130_fd_sc_hd__and2_1 _13833_ (.A(_06997_),
    .B(_07003_),
    .X(_07005_));
 sky130_fd_sc_hd__nor2_1 _13834_ (.A(_07004_),
    .B(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__xnor2_1 _13835_ (.A(_06996_),
    .B(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__xnor2_2 _13836_ (.A(_06970_),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__xnor2_2 _13837_ (.A(_06901_),
    .B(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__xnor2_1 _13838_ (.A(_06884_),
    .B(_06887_),
    .Y(_07010_));
 sky130_fd_sc_hd__nor2_1 _13839_ (.A(_06959_),
    .B(_06916_),
    .Y(_07011_));
 sky130_fd_sc_hd__nor4_1 _13840_ (.A(_06862_),
    .B(_06877_),
    .C(_06943_),
    .D(_06873_),
    .Y(_07012_));
 sky130_fd_sc_hd__o22a_1 _13841_ (.A1(_06862_),
    .A2(_06871_),
    .B1(_06873_),
    .B2(_06877_),
    .X(_07013_));
 sky130_fd_sc_hd__nor2_1 _13842_ (.A(_07012_),
    .B(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__a21o_1 _13843_ (.A1(_07011_),
    .A2(_07014_),
    .B1(_07012_),
    .X(_07015_));
 sky130_fd_sc_hd__or2b_1 _13844_ (.A(_07010_),
    .B_N(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__nor2_2 _13845_ (.A(_06716_),
    .B(_06863_),
    .Y(_07017_));
 sky130_fd_sc_hd__nor2_1 _13846_ (.A(_06845_),
    .B(_06860_),
    .Y(_07018_));
 sky130_fd_sc_hd__a21o_1 _13847_ (.A1(_06846_),
    .A2(_06865_),
    .B1(_06715_),
    .X(_07019_));
 sky130_fd_sc_hd__xnor2_1 _13848_ (.A(_06883_),
    .B(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__a22oi_2 _13849_ (.A1(_06886_),
    .A2(_07017_),
    .B1(_07018_),
    .B2(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__xnor2_1 _13850_ (.A(_07015_),
    .B(_07010_),
    .Y(_07022_));
 sky130_fd_sc_hd__or2b_1 _13851_ (.A(_07021_),
    .B_N(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__xnor2_1 _13852_ (.A(_06896_),
    .B(_06897_),
    .Y(_07024_));
 sky130_fd_sc_hd__a21oi_1 _13853_ (.A1(_07016_),
    .A2(_07023_),
    .B1(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__xnor2_1 _13854_ (.A(_06931_),
    .B(_06933_),
    .Y(_07026_));
 sky130_fd_sc_hd__a21oi_1 _13855_ (.A1(_06847_),
    .A2(_06911_),
    .B1(_06928_),
    .Y(_07027_));
 sky130_fd_sc_hd__xor2_2 _13856_ (.A(_06926_),
    .B(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__or4b_1 _13857_ (.A(_06893_),
    .B(_06825_),
    .C(_06902_),
    .D_N(_06742_),
    .X(_07029_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(_06816_),
    .B(_06925_),
    .Y(_07030_));
 sky130_fd_sc_hd__a2bb2o_1 _13859_ (.A1_N(_06825_),
    .A2_N(_06902_),
    .B1(_06908_),
    .B2(_06742_),
    .X(_07031_));
 sky130_fd_sc_hd__nand3_1 _13860_ (.A(_07029_),
    .B(_07030_),
    .C(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__and2_1 _13861_ (.A(_07029_),
    .B(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__xnor2_2 _13862_ (.A(_07028_),
    .B(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__xnor2_2 _13863_ (.A(_07011_),
    .B(_07014_),
    .Y(_07035_));
 sky130_fd_sc_hd__or2_1 _13864_ (.A(_07028_),
    .B(_07033_),
    .X(_07036_));
 sky130_fd_sc_hd__o21ai_1 _13865_ (.A1(_07034_),
    .A2(_07035_),
    .B1(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__xnor2_1 _13866_ (.A(_07026_),
    .B(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__xnor2_1 _13867_ (.A(_07021_),
    .B(_07022_),
    .Y(_07039_));
 sky130_fd_sc_hd__and2b_1 _13868_ (.A_N(_07026_),
    .B(_07037_),
    .X(_07040_));
 sky130_fd_sc_hd__a21oi_1 _13869_ (.A1(_07038_),
    .A2(_07039_),
    .B1(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__xnor2_1 _13870_ (.A(_06936_),
    .B(_06937_),
    .Y(_07042_));
 sky130_fd_sc_hd__xnor2_1 _13871_ (.A(_07041_),
    .B(_07042_),
    .Y(_07043_));
 sky130_fd_sc_hd__nand2_1 _13872_ (.A(_07016_),
    .B(_07023_),
    .Y(_07044_));
 sky130_fd_sc_hd__xor2_1 _13873_ (.A(_07044_),
    .B(_07024_),
    .X(_07045_));
 sky130_fd_sc_hd__or2_1 _13874_ (.A(_07041_),
    .B(_07042_),
    .X(_07046_));
 sky130_fd_sc_hd__o21a_1 _13875_ (.A1(_07043_),
    .A2(_07045_),
    .B1(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__xor2_1 _13876_ (.A(_06967_),
    .B(_06968_),
    .X(_07048_));
 sky130_fd_sc_hd__xnor2_1 _13877_ (.A(_07047_),
    .B(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__or2b_1 _13878_ (.A(_07047_),
    .B_N(_07048_),
    .X(_07050_));
 sky130_fd_sc_hd__a21boi_2 _13879_ (.A1(_07025_),
    .A2(_07049_),
    .B1_N(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__xnor2_2 _13880_ (.A(_07009_),
    .B(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__xnor2_1 _13881_ (.A(_07018_),
    .B(_07020_),
    .Y(_07053_));
 sky130_fd_sc_hd__or2_1 _13882_ (.A(_06805_),
    .B(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__clkbuf_4 _13883_ (.A(_06908_),
    .X(_07055_));
 sky130_fd_sc_hd__xnor2_4 _13884_ (.A(_06743_),
    .B(_06846_),
    .Y(_07056_));
 sky130_fd_sc_hd__a21oi_4 _13885_ (.A1(_06846_),
    .A2(_06865_),
    .B1(_06845_),
    .Y(_07057_));
 sky130_fd_sc_hd__xor2_2 _13886_ (.A(_07017_),
    .B(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__a32oi_4 _13887_ (.A1(_07055_),
    .A2(_07056_),
    .A3(_07058_),
    .B1(_07057_),
    .B2(_07017_),
    .Y(_07059_));
 sky130_fd_sc_hd__xnor2_1 _13888_ (.A(_06876_),
    .B(_07053_),
    .Y(_07060_));
 sky130_fd_sc_hd__or2b_1 _13889_ (.A(_07059_),
    .B_N(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__inv_2 _13890_ (.A(_06850_),
    .Y(_07062_));
 sky130_fd_sc_hd__clkinv_2 _13891_ (.A(_06841_),
    .Y(_07063_));
 sky130_fd_sc_hd__a22o_1 _13892_ (.A1(_07055_),
    .A2(_07062_),
    .B1(_07063_),
    .B2(_06844_),
    .X(_07064_));
 sky130_fd_sc_hd__nand2_1 _13893_ (.A(_06896_),
    .B(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__a21oi_1 _13894_ (.A1(_07054_),
    .A2(_07061_),
    .B1(_07065_),
    .Y(_07066_));
 sky130_fd_sc_hd__or2_1 _13895_ (.A(_07034_),
    .B(_07035_),
    .X(_07067_));
 sky130_fd_sc_hd__nand2_1 _13896_ (.A(_07034_),
    .B(_07035_),
    .Y(_07068_));
 sky130_fd_sc_hd__a21o_1 _13897_ (.A1(_07029_),
    .A2(_07031_),
    .B1(_07030_),
    .X(_07069_));
 sky130_fd_sc_hd__nand2_2 _13898_ (.A(_07032_),
    .B(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__or2_1 _13899_ (.A(_06862_),
    .B(_06925_),
    .X(_07071_));
 sky130_fd_sc_hd__nor2_1 _13900_ (.A(_06893_),
    .B(_06816_),
    .Y(_07072_));
 sky130_fd_sc_hd__or3b_1 _13901_ (.A(_06825_),
    .B(_06902_),
    .C_N(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__o22ai_1 _13902_ (.A1(_06893_),
    .A2(_06878_),
    .B1(_06877_),
    .B2(_06902_),
    .Y(_07074_));
 sky130_fd_sc_hd__nand2_1 _13903_ (.A(_07073_),
    .B(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__o21a_1 _13904_ (.A1(_07071_),
    .A2(_07075_),
    .B1(_07073_),
    .X(_07076_));
 sky130_fd_sc_hd__xnor2_2 _13905_ (.A(_07070_),
    .B(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__mux2_1 _13906_ (.A0(_06873_),
    .A1(_06853_),
    .S(_06862_),
    .X(_07078_));
 sky130_fd_sc_hd__o22ai_4 _13907_ (.A1(_07070_),
    .A2(_07076_),
    .B1(_07077_),
    .B2(_07078_),
    .Y(_07079_));
 sky130_fd_sc_hd__xnor2_1 _13908_ (.A(_07034_),
    .B(_07035_),
    .Y(_07080_));
 sky130_fd_sc_hd__xnor2_2 _13909_ (.A(_07080_),
    .B(_07079_),
    .Y(_07081_));
 sky130_fd_sc_hd__xnor2_2 _13910_ (.A(_07059_),
    .B(_07060_),
    .Y(_07082_));
 sky130_fd_sc_hd__a32oi_4 _13911_ (.A1(_07067_),
    .A2(_07068_),
    .A3(_07079_),
    .B1(_07081_),
    .B2(_07082_),
    .Y(_07083_));
 sky130_fd_sc_hd__xnor2_1 _13912_ (.A(_07038_),
    .B(_07039_),
    .Y(_07084_));
 sky130_fd_sc_hd__xor2_1 _13913_ (.A(_07083_),
    .B(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__and3_1 _13914_ (.A(_07054_),
    .B(_07061_),
    .C(_07065_),
    .X(_07086_));
 sky130_fd_sc_hd__nor2_1 _13915_ (.A(_07066_),
    .B(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__nor2_1 _13916_ (.A(_07083_),
    .B(_07084_),
    .Y(_07088_));
 sky130_fd_sc_hd__a21oi_1 _13917_ (.A1(_07085_),
    .A2(_07087_),
    .B1(_07088_),
    .Y(_07089_));
 sky130_fd_sc_hd__xnor2_1 _13918_ (.A(_07043_),
    .B(_07045_),
    .Y(_07090_));
 sky130_fd_sc_hd__xor2_1 _13919_ (.A(_07089_),
    .B(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__xnor2_1 _13920_ (.A(_07066_),
    .B(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__nand2_1 _13921_ (.A(_06869_),
    .B(_06716_),
    .Y(_07093_));
 sky130_fd_sc_hd__nor2_1 _13922_ (.A(_06959_),
    .B(_06853_),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2_1 _13923_ (.A(_06908_),
    .B(_07056_),
    .Y(_07095_));
 sky130_fd_sc_hd__xnor2_1 _13924_ (.A(_07095_),
    .B(_07058_),
    .Y(_07096_));
 sky130_fd_sc_hd__xnor2_1 _13925_ (.A(_06875_),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__inv_2 _13926_ (.A(_06863_),
    .Y(_07098_));
 sky130_fd_sc_hd__and3_1 _13927_ (.A(_07055_),
    .B(_07098_),
    .C(_07057_),
    .X(_07099_));
 sky130_fd_sc_hd__and2_1 _13928_ (.A(_07097_),
    .B(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__a31o_1 _13929_ (.A1(_07093_),
    .A2(_07094_),
    .A3(_07096_),
    .B1(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__and3_1 _13930_ (.A(_07055_),
    .B(_07063_),
    .C(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__xor2_1 _13931_ (.A(_07077_),
    .B(_07078_),
    .X(_07103_));
 sky130_fd_sc_hd__xnor2_1 _13932_ (.A(_07071_),
    .B(_07075_),
    .Y(_07104_));
 sky130_fd_sc_hd__nor2_1 _13933_ (.A(_06804_),
    .B(_06902_),
    .Y(_07105_));
 sky130_fd_sc_hd__or2_1 _13934_ (.A(_06779_),
    .B(_06925_),
    .X(_07106_));
 sky130_fd_sc_hd__xnor2_1 _13935_ (.A(_07072_),
    .B(_07105_),
    .Y(_07107_));
 sky130_fd_sc_hd__o2bb2a_1 _13936_ (.A1_N(_07072_),
    .A2_N(_07105_),
    .B1(_07106_),
    .B2(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__xnor2_1 _13937_ (.A(_07104_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__and2_1 _13938_ (.A(_06959_),
    .B(_06853_),
    .X(_07110_));
 sky130_fd_sc_hd__o32a_1 _13939_ (.A1(_07093_),
    .A2(_07094_),
    .A3(_07110_),
    .B1(_06916_),
    .B2(_06716_),
    .X(_07111_));
 sky130_fd_sc_hd__or2_1 _13940_ (.A(_07104_),
    .B(_07108_),
    .X(_07112_));
 sky130_fd_sc_hd__o21a_1 _13941_ (.A1(_07109_),
    .A2(_07111_),
    .B1(_07112_),
    .X(_07113_));
 sky130_fd_sc_hd__xnor2_1 _13942_ (.A(_07103_),
    .B(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__xor2_1 _13943_ (.A(_07097_),
    .B(_07099_),
    .X(_07115_));
 sky130_fd_sc_hd__and2b_1 _13944_ (.A_N(_07113_),
    .B(_07103_),
    .X(_07116_));
 sky130_fd_sc_hd__a21oi_1 _13945_ (.A1(_07114_),
    .A2(_07115_),
    .B1(_07116_),
    .Y(_07117_));
 sky130_fd_sc_hd__xnor2_1 _13946_ (.A(_07081_),
    .B(_07082_),
    .Y(_07118_));
 sky130_fd_sc_hd__xnor2_1 _13947_ (.A(_07117_),
    .B(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__xor2_1 _13948_ (.A(_06895_),
    .B(_07101_),
    .X(_07120_));
 sky130_fd_sc_hd__or2_1 _13949_ (.A(_07117_),
    .B(_07118_),
    .X(_07121_));
 sky130_fd_sc_hd__o21a_1 _13950_ (.A1(_07119_),
    .A2(_07120_),
    .B1(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__xor2_1 _13951_ (.A(_07085_),
    .B(_07087_),
    .X(_07123_));
 sky130_fd_sc_hd__xnor2_1 _13952_ (.A(_07122_),
    .B(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__and2b_1 _13953_ (.A_N(_07122_),
    .B(_07123_),
    .X(_07125_));
 sky130_fd_sc_hd__a21oi_1 _13954_ (.A1(_07102_),
    .A2(_07124_),
    .B1(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__nor2_1 _13955_ (.A(_07092_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__xnor2_1 _13956_ (.A(_07025_),
    .B(_07049_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand2_1 _13957_ (.A(_07066_),
    .B(_07091_),
    .Y(_07129_));
 sky130_fd_sc_hd__o21a_1 _13958_ (.A1(_07089_),
    .A2(_07090_),
    .B1(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__nor2_1 _13959_ (.A(_07128_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__and2_1 _13960_ (.A(_07128_),
    .B(_07130_),
    .X(_07132_));
 sky130_fd_sc_hd__nor2_1 _13961_ (.A(_07131_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_1 _13962_ (.A(_07127_),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__xor2_1 _13963_ (.A(_07102_),
    .B(_07124_),
    .X(_07135_));
 sky130_fd_sc_hd__xnor2_1 _13964_ (.A(_07106_),
    .B(_07107_),
    .Y(_07136_));
 sky130_fd_sc_hd__nor2_1 _13965_ (.A(_06893_),
    .B(_06779_),
    .Y(_07137_));
 sky130_fd_sc_hd__or2_1 _13966_ (.A(_06853_),
    .B(_06925_),
    .X(_07138_));
 sky130_fd_sc_hd__buf_2 _13967_ (.A(_06902_),
    .X(_07139_));
 sky130_fd_sc_hd__o22a_1 _13968_ (.A1(_06893_),
    .A2(_06804_),
    .B1(_07139_),
    .B2(_06779_),
    .X(_07140_));
 sky130_fd_sc_hd__a21o_1 _13969_ (.A1(_07105_),
    .A2(_07137_),
    .B1(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__o2bb2a_1 _13970_ (.A1_N(_07105_),
    .A2_N(_07137_),
    .B1(_07138_),
    .B2(_07141_),
    .X(_07142_));
 sky130_fd_sc_hd__or2_1 _13971_ (.A(_07136_),
    .B(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__nor2_1 _13972_ (.A(_06845_),
    .B(_06916_),
    .Y(_07144_));
 sky130_fd_sc_hd__nor2_1 _13973_ (.A(_06869_),
    .B(_06853_),
    .Y(_07145_));
 sky130_fd_sc_hd__mux2_1 _13974_ (.A0(_06959_),
    .A1(_07145_),
    .S(_06716_),
    .X(_07146_));
 sky130_fd_sc_hd__xnor2_1 _13975_ (.A(_07144_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__xnor2_1 _13976_ (.A(_07136_),
    .B(_07142_),
    .Y(_07148_));
 sky130_fd_sc_hd__or2_1 _13977_ (.A(_07147_),
    .B(_07148_),
    .X(_07149_));
 sky130_fd_sc_hd__xnor2_1 _13978_ (.A(_07109_),
    .B(_07111_),
    .Y(_07150_));
 sky130_fd_sc_hd__a21o_1 _13979_ (.A1(_07143_),
    .A2(_07149_),
    .B1(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__clkbuf_4 _13980_ (.A(_06863_),
    .X(_07152_));
 sky130_fd_sc_hd__o22a_1 _13981_ (.A1(_06893_),
    .A2(_06954_),
    .B1(_07152_),
    .B2(_06845_),
    .X(_07153_));
 sky130_fd_sc_hd__nor2_1 _13982_ (.A(_07099_),
    .B(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__or2_1 _13983_ (.A(_06779_),
    .B(_06792_),
    .X(_07155_));
 sky130_fd_sc_hd__a2bb2o_1 _13984_ (.A1_N(_06716_),
    .A2_N(_07155_),
    .B1(_07144_),
    .B2(_07146_),
    .X(_07156_));
 sky130_fd_sc_hd__nand2_1 _13985_ (.A(_07154_),
    .B(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__or2_1 _13986_ (.A(_07154_),
    .B(_07156_),
    .X(_07158_));
 sky130_fd_sc_hd__and2_1 _13987_ (.A(_07157_),
    .B(_07158_),
    .X(_07159_));
 sky130_fd_sc_hd__nand3_1 _13988_ (.A(_07150_),
    .B(_07143_),
    .C(_07149_),
    .Y(_07160_));
 sky130_fd_sc_hd__nand3_1 _13989_ (.A(_07151_),
    .B(_07159_),
    .C(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__xnor2_1 _13990_ (.A(_07114_),
    .B(_07115_),
    .Y(_07162_));
 sky130_fd_sc_hd__a21oi_1 _13991_ (.A1(_07151_),
    .A2(_07161_),
    .B1(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__and3_1 _13992_ (.A(_07151_),
    .B(_07161_),
    .C(_07162_),
    .X(_07164_));
 sky130_fd_sc_hd__or2_1 _13993_ (.A(_07163_),
    .B(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__nor2_1 _13994_ (.A(_07157_),
    .B(_07165_),
    .Y(_07166_));
 sky130_fd_sc_hd__xor2_1 _13995_ (.A(_07119_),
    .B(_07120_),
    .X(_07167_));
 sky130_fd_sc_hd__o21a_1 _13996_ (.A1(_07163_),
    .A2(_07166_),
    .B1(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__xor2_1 _13997_ (.A(_07092_),
    .B(_07126_),
    .X(_07169_));
 sky130_fd_sc_hd__and3_1 _13998_ (.A(_07135_),
    .B(_07168_),
    .C(_07169_),
    .X(_07170_));
 sky130_fd_sc_hd__nand2_1 _13999_ (.A(_07135_),
    .B(_07168_),
    .Y(_07171_));
 sky130_fd_sc_hd__xnor2_1 _14000_ (.A(_07171_),
    .B(_07169_),
    .Y(_07172_));
 sky130_fd_sc_hd__or3_1 _14001_ (.A(_07167_),
    .B(_07163_),
    .C(_07166_),
    .X(_07173_));
 sky130_fd_sc_hd__and3b_1 _14002_ (.A_N(_07168_),
    .B(_07173_),
    .C(_07135_),
    .X(_07174_));
 sky130_fd_sc_hd__and2_1 _14003_ (.A(_07157_),
    .B(_07165_),
    .X(_07175_));
 sky130_fd_sc_hd__nor2_1 _14004_ (.A(_07166_),
    .B(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__nor2_1 _14005_ (.A(_06716_),
    .B(_06853_),
    .Y(_07177_));
 sky130_fd_sc_hd__nor2_1 _14006_ (.A(_06845_),
    .B(_06943_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_1 _14007_ (.A(_07177_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__xnor2_1 _14008_ (.A(_07177_),
    .B(_07178_),
    .Y(_07180_));
 sky130_fd_sc_hd__nand2_1 _14009_ (.A(_07055_),
    .B(_06975_),
    .Y(_07181_));
 sky130_fd_sc_hd__or2_1 _14010_ (.A(_07180_),
    .B(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__or2_1 _14011_ (.A(_06894_),
    .B(_07152_),
    .X(_07183_));
 sky130_fd_sc_hd__a21o_1 _14012_ (.A1(_07179_),
    .A2(_07182_),
    .B1(_07183_),
    .X(_07184_));
 sky130_fd_sc_hd__a21o_1 _14013_ (.A1(_07151_),
    .A2(_07160_),
    .B1(_07159_),
    .X(_07185_));
 sky130_fd_sc_hd__and2_1 _14014_ (.A(_07161_),
    .B(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__nand2_1 _14015_ (.A(_07147_),
    .B(_07148_),
    .Y(_07187_));
 sky130_fd_sc_hd__xnor2_1 _14016_ (.A(_07138_),
    .B(_07141_),
    .Y(_07188_));
 sky130_fd_sc_hd__a21o_1 _14017_ (.A1(_06844_),
    .A2(_07055_),
    .B1(_06716_),
    .X(_07189_));
 sky130_fd_sc_hd__o21ba_1 _14018_ (.A1(_06853_),
    .A2(_07139_),
    .B1_N(_07137_),
    .X(_07190_));
 sky130_fd_sc_hd__or2_1 _14019_ (.A(_06869_),
    .B(_07155_),
    .X(_07191_));
 sky130_fd_sc_hd__o21a_1 _14020_ (.A1(_07189_),
    .A2(_07190_),
    .B1(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__or2_1 _14021_ (.A(_07188_),
    .B(_07192_),
    .X(_07193_));
 sky130_fd_sc_hd__nand2_1 _14022_ (.A(_07180_),
    .B(_07181_),
    .Y(_07194_));
 sky130_fd_sc_hd__nand2_1 _14023_ (.A(_07182_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__nand2_1 _14024_ (.A(_07188_),
    .B(_07192_),
    .Y(_07196_));
 sky130_fd_sc_hd__nand2_1 _14025_ (.A(_07193_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__or2_1 _14026_ (.A(_07195_),
    .B(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__nand2_1 _14027_ (.A(_07193_),
    .B(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__nand3_1 _14028_ (.A(_07183_),
    .B(_07179_),
    .C(_07182_),
    .Y(_07200_));
 sky130_fd_sc_hd__nand2_1 _14029_ (.A(_07184_),
    .B(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__nand2_1 _14030_ (.A(_07149_),
    .B(_07187_),
    .Y(_07202_));
 sky130_fd_sc_hd__xnor2_1 _14031_ (.A(_07202_),
    .B(_07199_),
    .Y(_07203_));
 sky130_fd_sc_hd__and2b_1 _14032_ (.A_N(_07201_),
    .B(_07203_),
    .X(_07204_));
 sky130_fd_sc_hd__a31o_1 _14033_ (.A1(_07149_),
    .A2(_07187_),
    .A3(_07199_),
    .B1(_07204_),
    .X(_07205_));
 sky130_fd_sc_hd__xnor2_1 _14034_ (.A(_07186_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand2_1 _14035_ (.A(_07186_),
    .B(_07205_),
    .Y(_07207_));
 sky130_fd_sc_hd__o21ai_1 _14036_ (.A1(_07184_),
    .A2(_07206_),
    .B1(_07207_),
    .Y(_07208_));
 sky130_fd_sc_hd__and3_1 _14037_ (.A(_07174_),
    .B(_07176_),
    .C(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__xor2_1 _14038_ (.A(_07172_),
    .B(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__a2bb2o_1 _14039_ (.A1_N(_06894_),
    .A2_N(_06943_),
    .B1(_06919_),
    .B2(_06844_),
    .X(_07211_));
 sky130_fd_sc_hd__a21boi_1 _14040_ (.A1(_07189_),
    .A2(_07190_),
    .B1_N(_07192_),
    .Y(_07212_));
 sky130_fd_sc_hd__nand2_1 _14041_ (.A(_07195_),
    .B(_07197_),
    .Y(_07213_));
 sky130_fd_sc_hd__and2_1 _14042_ (.A(_07198_),
    .B(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__a21oi_1 _14043_ (.A1(_07211_),
    .A2(_07212_),
    .B1(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__o21ai_1 _14044_ (.A1(_06844_),
    .A2(_07177_),
    .B1(_07055_),
    .Y(_07216_));
 sky130_fd_sc_hd__xor2_1 _14045_ (.A(_07201_),
    .B(_07203_),
    .X(_07217_));
 sky130_fd_sc_hd__o211ai_1 _14046_ (.A1(_07215_),
    .A2(_07216_),
    .B1(_07191_),
    .C1(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__a32o_1 _14047_ (.A1(_07214_),
    .A2(_07211_),
    .A3(_07212_),
    .B1(_07145_),
    .B2(_06959_),
    .X(_07219_));
 sky130_fd_sc_hd__a21boi_1 _14048_ (.A1(_07184_),
    .A2(_07206_),
    .B1_N(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__o2111a_1 _14049_ (.A1(_07176_),
    .A2(_07208_),
    .B1(_07218_),
    .C1(_07220_),
    .D1(_07174_),
    .X(_07221_));
 sky130_fd_sc_hd__nand2_1 _14050_ (.A(_07172_),
    .B(_07209_),
    .Y(_07222_));
 sky130_fd_sc_hd__a21bo_1 _14051_ (.A1(_07210_),
    .A2(_07221_),
    .B1_N(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__nor2_1 _14052_ (.A(_07127_),
    .B(_07170_),
    .Y(_07224_));
 sky130_fd_sc_hd__xnor2_1 _14053_ (.A(_07133_),
    .B(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__a22o_1 _14054_ (.A1(_07133_),
    .A2(_07170_),
    .B1(_07223_),
    .B2(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__a21o_1 _14055_ (.A1(_07127_),
    .A2(_07133_),
    .B1(_07131_),
    .X(_07227_));
 sky130_fd_sc_hd__xnor2_1 _14056_ (.A(_07052_),
    .B(_07227_),
    .Y(_07228_));
 sky130_fd_sc_hd__a2bb2o_2 _14057_ (.A1_N(_07052_),
    .A2_N(_07134_),
    .B1(_07226_),
    .B2(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__a21o_1 _14058_ (.A1(_06999_),
    .A2(_07002_),
    .B1(_07004_),
    .X(_07230_));
 sky130_fd_sc_hd__or2b_1 _14059_ (.A(_06996_),
    .B_N(_07006_),
    .X(_07231_));
 sky130_fd_sc_hd__or2b_1 _14060_ (.A(_06981_),
    .B_N(_06992_),
    .X(_07232_));
 sky130_fd_sc_hd__nor2_1 _14061_ (.A(_06648_),
    .B(_06943_),
    .Y(_07233_));
 sky130_fd_sc_hd__and2_1 _14062_ (.A(_06975_),
    .B(_06840_),
    .X(_07234_));
 sky130_fd_sc_hd__xnor2_1 _14063_ (.A(_07233_),
    .B(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__clkbuf_4 _14064_ (.A(_06873_),
    .X(_07236_));
 sky130_fd_sc_hd__o22ai_2 _14065_ (.A1(_07236_),
    .A2(_06972_),
    .B1(_06974_),
    .B2(_06976_),
    .Y(_07237_));
 sky130_fd_sc_hd__o2bb2a_1 _14066_ (.A1_N(_06877_),
    .A2_N(_07056_),
    .B1(_07098_),
    .B2(_06743_),
    .X(_07238_));
 sky130_fd_sc_hd__xnor2_1 _14067_ (.A(_07237_),
    .B(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__a21oi_1 _14068_ (.A1(_06876_),
    .A2(_06743_),
    .B1(_06846_),
    .Y(_07240_));
 sky130_fd_sc_hd__xor2_1 _14069_ (.A(_07239_),
    .B(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__or2_1 _14070_ (.A(_07235_),
    .B(_07241_),
    .X(_07242_));
 sky130_fd_sc_hd__nand2_1 _14071_ (.A(_07235_),
    .B(_07241_),
    .Y(_07243_));
 sky130_fd_sc_hd__nand2_1 _14072_ (.A(_07242_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__a21o_1 _14073_ (.A1(_06979_),
    .A2(_07232_),
    .B1(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__nand3_1 _14074_ (.A(_06979_),
    .B(_07232_),
    .C(_07244_),
    .Y(_07246_));
 sky130_fd_sc_hd__and2_1 _14075_ (.A(_07245_),
    .B(_07246_),
    .X(_07247_));
 sky130_fd_sc_hd__or2b_1 _14076_ (.A(_06855_),
    .B_N(_07001_),
    .X(_07248_));
 sky130_fd_sc_hd__and2b_1 _14077_ (.A_N(_06991_),
    .B(_06983_),
    .X(_07249_));
 sky130_fd_sc_hd__nor2_1 _14078_ (.A(_06862_),
    .B(_06841_),
    .Y(_07250_));
 sky130_fd_sc_hd__or2_1 _14079_ (.A(_06959_),
    .B(_06850_),
    .X(_07251_));
 sky130_fd_sc_hd__or3b_1 _14080_ (.A(_07250_),
    .B(_07251_),
    .C_N(_06856_),
    .X(_07252_));
 sky130_fd_sc_hd__xnor2_1 _14081_ (.A(_07251_),
    .B(_07250_),
    .Y(_07253_));
 sky130_fd_sc_hd__a21o_1 _14082_ (.A1(_06854_),
    .A2(_07000_),
    .B1(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__and2_1 _14083_ (.A(_07252_),
    .B(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__o21ai_1 _14084_ (.A1(_06989_),
    .A2(_07249_),
    .B1(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__or3_1 _14085_ (.A(_06989_),
    .B(_07249_),
    .C(_07255_),
    .X(_07257_));
 sky130_fd_sc_hd__nand2_1 _14086_ (.A(_07256_),
    .B(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__xor2_1 _14087_ (.A(_07248_),
    .B(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__xnor2_1 _14088_ (.A(_07247_),
    .B(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__a21o_1 _14089_ (.A1(_06994_),
    .A2(_07231_),
    .B1(_07260_),
    .X(_07261_));
 sky130_fd_sc_hd__nand3_1 _14090_ (.A(_06994_),
    .B(_07231_),
    .C(_07260_),
    .Y(_07262_));
 sky130_fd_sc_hd__and2_1 _14091_ (.A(_07261_),
    .B(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__xnor2_2 _14092_ (.A(_07230_),
    .B(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__or2b_1 _14093_ (.A(_06970_),
    .B_N(_07007_),
    .X(_07265_));
 sky130_fd_sc_hd__a21boi_2 _14094_ (.A1(_06901_),
    .A2(_07008_),
    .B1_N(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__xor2_2 _14095_ (.A(_07264_),
    .B(_07266_),
    .X(_07267_));
 sky130_fd_sc_hd__and2b_1 _14096_ (.A_N(_07052_),
    .B(_07131_),
    .X(_07268_));
 sky130_fd_sc_hd__nor2_1 _14097_ (.A(_07009_),
    .B(_07051_),
    .Y(_07269_));
 sky130_fd_sc_hd__nor3_1 _14098_ (.A(_07269_),
    .B(_07267_),
    .C(_07268_),
    .Y(_07270_));
 sky130_fd_sc_hd__and2_1 _14099_ (.A(_07269_),
    .B(_07267_),
    .X(_07271_));
 sky130_fd_sc_hd__a211oi_2 _14100_ (.A1(_07267_),
    .A2(_07268_),
    .B1(_07270_),
    .C1(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__xnor2_2 _14101_ (.A(_07229_),
    .B(_07272_),
    .Y(_07273_));
 sky130_fd_sc_hd__xor2_1 _14102_ (.A(_07226_),
    .B(_07228_),
    .X(_07274_));
 sky130_fd_sc_hd__xnor2_1 _14103_ (.A(_07223_),
    .B(_07225_),
    .Y(_07275_));
 sky130_fd_sc_hd__xnor2_1 _14104_ (.A(_07210_),
    .B(_07221_),
    .Y(_07276_));
 sky130_fd_sc_hd__nor2_1 _14105_ (.A(_07275_),
    .B(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__nor2_1 _14106_ (.A(_07274_),
    .B(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__nand2_1 _14107_ (.A(_07273_),
    .B(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__a22o_1 _14108_ (.A1(_07267_),
    .A2(_07268_),
    .B1(_07272_),
    .B2(_07229_),
    .X(_07280_));
 sky130_fd_sc_hd__nand2_1 _14109_ (.A(_07230_),
    .B(_07263_),
    .Y(_07281_));
 sky130_fd_sc_hd__o21a_1 _14110_ (.A1(_07248_),
    .A2(_07258_),
    .B1(_07256_),
    .X(_07282_));
 sky130_fd_sc_hd__nand2_1 _14111_ (.A(_07247_),
    .B(_07259_),
    .Y(_07283_));
 sky130_fd_sc_hd__nor2_1 _14112_ (.A(_06648_),
    .B(_06916_),
    .Y(_07284_));
 sky130_fd_sc_hd__nand2_1 _14113_ (.A(_07233_),
    .B(_07234_),
    .Y(_07285_));
 sky130_fd_sc_hd__nor2_1 _14114_ (.A(_06878_),
    .B(_06860_),
    .Y(_07286_));
 sky130_fd_sc_hd__nand2_1 _14115_ (.A(_06840_),
    .B(_07098_),
    .Y(_07287_));
 sky130_fd_sc_hd__nand2_2 _14116_ (.A(_06846_),
    .B(_06865_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand2_1 _14117_ (.A(_06847_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__xnor2_1 _14118_ (.A(_07287_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__xnor2_1 _14119_ (.A(_07286_),
    .B(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__xor2_1 _14120_ (.A(_07285_),
    .B(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__xor2_1 _14121_ (.A(_06828_),
    .B(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__xnor2_1 _14122_ (.A(_07284_),
    .B(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__or2_1 _14123_ (.A(_07242_),
    .B(_07294_),
    .X(_07295_));
 sky130_fd_sc_hd__nand2_1 _14124_ (.A(_07242_),
    .B(_07294_),
    .Y(_07296_));
 sky130_fd_sc_hd__nand2_1 _14125_ (.A(_07295_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__or2b_1 _14126_ (.A(_07239_),
    .B_N(_07240_),
    .X(_07298_));
 sky130_fd_sc_hd__a21bo_1 _14127_ (.A1(_07237_),
    .A2(_07238_),
    .B1_N(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__or2_1 _14128_ (.A(_06862_),
    .B(_06850_),
    .X(_07300_));
 sky130_fd_sc_hd__or3_1 _14129_ (.A(_06959_),
    .B(_06841_),
    .C(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__nor2_1 _14130_ (.A(_06877_),
    .B(_06841_),
    .Y(_07302_));
 sky130_fd_sc_hd__xnor2_1 _14131_ (.A(_07300_),
    .B(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__xnor2_1 _14132_ (.A(_07301_),
    .B(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__xnor2_1 _14133_ (.A(_07299_),
    .B(_07304_),
    .Y(_07305_));
 sky130_fd_sc_hd__nor2_1 _14134_ (.A(_07252_),
    .B(_07305_),
    .Y(_07306_));
 sky130_fd_sc_hd__and2_1 _14135_ (.A(_07252_),
    .B(_07305_),
    .X(_07307_));
 sky130_fd_sc_hd__nor2_1 _14136_ (.A(_07306_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__xor2_1 _14137_ (.A(_07297_),
    .B(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__a21o_1 _14138_ (.A1(_07245_),
    .A2(_07283_),
    .B1(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__nand3_1 _14139_ (.A(_07245_),
    .B(_07283_),
    .C(_07309_),
    .Y(_07311_));
 sky130_fd_sc_hd__and2_1 _14140_ (.A(_07310_),
    .B(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__or2b_1 _14141_ (.A(_07282_),
    .B_N(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__or2b_1 _14142_ (.A(_07312_),
    .B_N(_07282_),
    .X(_07314_));
 sky130_fd_sc_hd__nand2_1 _14143_ (.A(_07313_),
    .B(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__a21oi_2 _14144_ (.A1(_07261_),
    .A2(_07281_),
    .B1(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__and3_1 _14145_ (.A(_07261_),
    .B(_07281_),
    .C(_07315_),
    .X(_07317_));
 sky130_fd_sc_hd__nor2_1 _14146_ (.A(_07316_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__nor2_1 _14147_ (.A(_07264_),
    .B(_07266_),
    .Y(_07319_));
 sky130_fd_sc_hd__nor2_1 _14148_ (.A(_07319_),
    .B(_07271_),
    .Y(_07320_));
 sky130_fd_sc_hd__xnor2_1 _14149_ (.A(_07318_),
    .B(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__xor2_2 _14150_ (.A(_07280_),
    .B(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__or2_1 _14151_ (.A(_07279_),
    .B(_07322_),
    .X(_07323_));
 sky130_fd_sc_hd__a22o_1 _14152_ (.A1(_07271_),
    .A2(_07318_),
    .B1(_07321_),
    .B2(_07280_),
    .X(_07324_));
 sky130_fd_sc_hd__or2b_1 _14153_ (.A(_07297_),
    .B_N(_07308_),
    .X(_07325_));
 sky130_fd_sc_hd__nand2_1 _14154_ (.A(_07284_),
    .B(_07293_),
    .Y(_07326_));
 sky130_fd_sc_hd__and2_1 _14155_ (.A(_06840_),
    .B(_07288_),
    .X(_07327_));
 sky130_fd_sc_hd__xnor2_1 _14156_ (.A(_07098_),
    .B(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__nor2_1 _14157_ (.A(_07326_),
    .B(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__and2_1 _14158_ (.A(_07326_),
    .B(_07328_),
    .X(_07330_));
 sky130_fd_sc_hd__or2_1 _14159_ (.A(_07329_),
    .B(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__or3b_1 _14160_ (.A(_07302_),
    .B(_07300_),
    .C_N(_07000_),
    .X(_07332_));
 sky130_fd_sc_hd__nor2_1 _14161_ (.A(_06828_),
    .B(_07292_),
    .Y(_07333_));
 sky130_fd_sc_hd__a31o_1 _14162_ (.A1(_07233_),
    .A2(_07234_),
    .A3(_07291_),
    .B1(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__buf_2 _14163_ (.A(_06841_),
    .X(_07335_));
 sky130_fd_sc_hd__or3_1 _14164_ (.A(_06877_),
    .B(_07335_),
    .C(_07300_),
    .X(_07336_));
 sky130_fd_sc_hd__and3b_1 _14165_ (.A_N(_06878_),
    .B(_07062_),
    .C(_07302_),
    .X(_07337_));
 sky130_fd_sc_hd__clkbuf_4 _14166_ (.A(_06850_),
    .X(_07338_));
 sky130_fd_sc_hd__o22a_1 _14167_ (.A1(_06877_),
    .A2(_07338_),
    .B1(_06841_),
    .B2(_06878_),
    .X(_07339_));
 sky130_fd_sc_hd__nor2_1 _14168_ (.A(_07337_),
    .B(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__xnor2_1 _14169_ (.A(_07336_),
    .B(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__xnor2_1 _14170_ (.A(_07334_),
    .B(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__xnor2_1 _14171_ (.A(_07332_),
    .B(_07342_),
    .Y(_07343_));
 sky130_fd_sc_hd__xnor2_1 _14172_ (.A(_07331_),
    .B(_07343_),
    .Y(_07344_));
 sky130_fd_sc_hd__a21oi_1 _14173_ (.A1(_07295_),
    .A2(_07325_),
    .B1(_07344_),
    .Y(_07345_));
 sky130_fd_sc_hd__and3_1 _14174_ (.A(_07295_),
    .B(_07325_),
    .C(_07344_),
    .X(_07346_));
 sky130_fd_sc_hd__nor2_1 _14175_ (.A(_07345_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__a21oi_1 _14176_ (.A1(_07299_),
    .A2(_07304_),
    .B1(_07306_),
    .Y(_07348_));
 sky130_fd_sc_hd__xor2_1 _14177_ (.A(_07347_),
    .B(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__a21oi_2 _14178_ (.A1(_07310_),
    .A2(_07313_),
    .B1(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__and3_1 _14179_ (.A(_07310_),
    .B(_07313_),
    .C(_07349_),
    .X(_07351_));
 sky130_fd_sc_hd__nor2_1 _14180_ (.A(_07350_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__xor2_1 _14181_ (.A(_07316_),
    .B(_07352_),
    .X(_07353_));
 sky130_fd_sc_hd__and3_1 _14182_ (.A(_07319_),
    .B(_07318_),
    .C(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__a21oi_1 _14183_ (.A1(_07319_),
    .A2(_07318_),
    .B1(_07353_),
    .Y(_07355_));
 sky130_fd_sc_hd__nor2_1 _14184_ (.A(_07354_),
    .B(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__xor2_2 _14185_ (.A(_07324_),
    .B(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__nor2_1 _14186_ (.A(_07323_),
    .B(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__a21o_1 _14187_ (.A1(_07324_),
    .A2(_07356_),
    .B1(_07354_),
    .X(_07359_));
 sky130_fd_sc_hd__nand2_1 _14188_ (.A(_07316_),
    .B(_07352_),
    .Y(_07360_));
 sky130_fd_sc_hd__and2b_1 _14189_ (.A_N(_07348_),
    .B(_07347_),
    .X(_07361_));
 sky130_fd_sc_hd__nor2_1 _14190_ (.A(_07331_),
    .B(_07343_),
    .Y(_07362_));
 sky130_fd_sc_hd__nor2_1 _14191_ (.A(_06828_),
    .B(_07328_),
    .Y(_07363_));
 sky130_fd_sc_hd__a21o_1 _14192_ (.A1(_07098_),
    .A2(_07327_),
    .B1(_07363_),
    .X(_07364_));
 sky130_fd_sc_hd__o2bb2a_1 _14193_ (.A1_N(_06840_),
    .A2_N(_07056_),
    .B1(_06954_),
    .B2(_06648_),
    .X(_07365_));
 sky130_fd_sc_hd__a31oi_1 _14194_ (.A1(_06849_),
    .A2(_07056_),
    .A3(_07327_),
    .B1(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__and2_1 _14195_ (.A(_07364_),
    .B(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__nor2_1 _14196_ (.A(_07364_),
    .B(_07366_),
    .Y(_07368_));
 sky130_fd_sc_hd__nor2_1 _14197_ (.A(_07367_),
    .B(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__or3_1 _14198_ (.A(_07336_),
    .B(_07337_),
    .C(_07339_),
    .X(_07370_));
 sky130_fd_sc_hd__nor2_1 _14199_ (.A(_06828_),
    .B(_07363_),
    .Y(_07371_));
 sky130_fd_sc_hd__o22a_1 _14200_ (.A1(_06878_),
    .A2(_07338_),
    .B1(_07335_),
    .B2(_06743_),
    .X(_07372_));
 sky130_fd_sc_hd__or4_1 _14201_ (.A(_06743_),
    .B(_06878_),
    .C(_07338_),
    .D(_07335_),
    .X(_07373_));
 sky130_fd_sc_hd__or3b_1 _14202_ (.A(_07337_),
    .B(_07372_),
    .C_N(_07373_),
    .X(_07374_));
 sky130_fd_sc_hd__or2_1 _14203_ (.A(_07371_),
    .B(_07374_),
    .X(_07375_));
 sky130_fd_sc_hd__xor2_1 _14204_ (.A(_07370_),
    .B(_07375_),
    .X(_07376_));
 sky130_fd_sc_hd__nand2_1 _14205_ (.A(_07369_),
    .B(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__or2_1 _14206_ (.A(_07369_),
    .B(_07376_),
    .X(_07378_));
 sky130_fd_sc_hd__and2_1 _14207_ (.A(_07377_),
    .B(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__o21a_1 _14208_ (.A1(_07329_),
    .A2(_07362_),
    .B1(_07379_),
    .X(_07380_));
 sky130_fd_sc_hd__nor3_1 _14209_ (.A(_07329_),
    .B(_07362_),
    .C(_07379_),
    .Y(_07381_));
 sky130_fd_sc_hd__nor2_1 _14210_ (.A(_07380_),
    .B(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__nor2_1 _14211_ (.A(_07332_),
    .B(_07342_),
    .Y(_07383_));
 sky130_fd_sc_hd__a21oi_1 _14212_ (.A1(_07334_),
    .A2(_07341_),
    .B1(_07383_),
    .Y(_07384_));
 sky130_fd_sc_hd__xnor2_1 _14213_ (.A(_07382_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__o21ai_1 _14214_ (.A1(_07345_),
    .A2(_07361_),
    .B1(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__or3_1 _14215_ (.A(_07345_),
    .B(_07361_),
    .C(_07385_),
    .X(_07387_));
 sky130_fd_sc_hd__and2_1 _14216_ (.A(_07386_),
    .B(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__xor2_1 _14217_ (.A(_07350_),
    .B(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__xnor2_1 _14218_ (.A(_07360_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__xnor2_2 _14219_ (.A(_07359_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__and2_1 _14220_ (.A(_07324_),
    .B(_07356_),
    .X(_07392_));
 sky130_fd_sc_hd__and2b_1 _14221_ (.A_N(_07384_),
    .B(_07382_),
    .X(_07393_));
 sky130_fd_sc_hd__and3_1 _14222_ (.A(_06847_),
    .B(_07367_),
    .C(_07373_),
    .X(_07394_));
 sky130_fd_sc_hd__a21oi_1 _14223_ (.A1(_06847_),
    .A2(_07373_),
    .B1(_07367_),
    .Y(_07395_));
 sky130_fd_sc_hd__nor2_1 _14224_ (.A(_07394_),
    .B(_07395_),
    .Y(_07396_));
 sky130_fd_sc_hd__o21ba_1 _14225_ (.A1(_07370_),
    .A2(_07375_),
    .B1_N(_07371_),
    .X(_07397_));
 sky130_fd_sc_hd__o21a_1 _14226_ (.A1(_07337_),
    .A2(_07396_),
    .B1(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__or3_1 _14227_ (.A(_06648_),
    .B(_06860_),
    .C(_07327_),
    .X(_07399_));
 sky130_fd_sc_hd__xor2_1 _14228_ (.A(_07377_),
    .B(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__xnor2_1 _14229_ (.A(_07398_),
    .B(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__or3_1 _14230_ (.A(_07380_),
    .B(_07393_),
    .C(_07401_),
    .X(_07402_));
 sky130_fd_sc_hd__o21a_1 _14231_ (.A1(_07287_),
    .A2(_07289_),
    .B1(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__nor2_1 _14232_ (.A(_07386_),
    .B(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__a221o_1 _14233_ (.A1(_07350_),
    .A2(_07388_),
    .B1(_07403_),
    .B2(_07386_),
    .C1(_07404_),
    .X(_07405_));
 sky130_fd_sc_hd__inv_2 _14234_ (.A(_07354_),
    .Y(_07406_));
 sky130_fd_sc_hd__a21boi_1 _14235_ (.A1(_07360_),
    .A2(_07406_),
    .B1_N(_07389_),
    .Y(_07407_));
 sky130_fd_sc_hd__a211o_1 _14236_ (.A1(_07392_),
    .A2(_07390_),
    .B1(_07405_),
    .C1(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__a21bo_2 _14237_ (.A1(_07358_),
    .A2(_07391_),
    .B1_N(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__buf_2 _14238_ (.A(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__buf_2 _14239_ (.A(_07410_),
    .X(_07411_));
 sky130_fd_sc_hd__xnor2_1 _14240_ (.A(_07279_),
    .B(_07322_),
    .Y(_07412_));
 sky130_fd_sc_hd__buf_2 _14241_ (.A(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__or2_1 _14242_ (.A(_07335_),
    .B(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__xnor2_2 _14243_ (.A(_07323_),
    .B(_07357_),
    .Y(_07415_));
 sky130_fd_sc_hd__clkbuf_4 _14244_ (.A(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__nor2_1 _14245_ (.A(_07338_),
    .B(_07416_),
    .Y(_07417_));
 sky130_fd_sc_hd__xor2_2 _14246_ (.A(_07358_),
    .B(_07391_),
    .X(_07418_));
 sky130_fd_sc_hd__buf_2 _14247_ (.A(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__nand2_1 _14248_ (.A(_07063_),
    .B(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__and3b_1 _14249_ (.A_N(_07414_),
    .B(_07417_),
    .C(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__buf_2 _14250_ (.A(_06954_),
    .X(_07422_));
 sky130_fd_sc_hd__or2_2 _14251_ (.A(_07152_),
    .B(_07410_),
    .X(_07423_));
 sky130_fd_sc_hd__or2_1 _14252_ (.A(_07422_),
    .B(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__nor2_1 _14253_ (.A(_07422_),
    .B(_07411_),
    .Y(_07425_));
 sky130_fd_sc_hd__xnor2_2 _14254_ (.A(_07423_),
    .B(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__buf_2 _14255_ (.A(_06860_),
    .X(_07427_));
 sky130_fd_sc_hd__nor2_1 _14256_ (.A(_07427_),
    .B(_07411_),
    .Y(_07428_));
 sky130_fd_sc_hd__nand2_1 _14257_ (.A(_07426_),
    .B(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__and3b_1 _14258_ (.A_N(_07411_),
    .B(_07288_),
    .C(_07056_),
    .X(_07430_));
 sky130_fd_sc_hd__a21o_1 _14259_ (.A1(_07424_),
    .A2(_07429_),
    .B1(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__or3b_1 _14260_ (.A(_07411_),
    .B(_07421_),
    .C_N(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__and2_2 _14261_ (.A(_06849_),
    .B(_07409_),
    .X(_07433_));
 sky130_fd_sc_hd__a21oi_1 _14262_ (.A1(_07288_),
    .A2(_07433_),
    .B1(_07428_),
    .Y(_07434_));
 sky130_fd_sc_hd__or2_1 _14263_ (.A(_07430_),
    .B(_07434_),
    .X(_07435_));
 sky130_fd_sc_hd__a211o_1 _14264_ (.A1(_07098_),
    .A2(_07433_),
    .B1(_07425_),
    .C1(_07428_),
    .X(_07436_));
 sky130_fd_sc_hd__buf_4 _14265_ (.A(_06648_),
    .X(_07437_));
 sky130_fd_sc_hd__a21o_1 _14266_ (.A1(_07431_),
    .A2(_07436_),
    .B1(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__nor2_1 _14267_ (.A(_07335_),
    .B(_07411_),
    .Y(_07439_));
 sky130_fd_sc_hd__nand2_1 _14268_ (.A(_07416_),
    .B(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__a31o_1 _14269_ (.A1(_07062_),
    .A2(_07419_),
    .A3(_07440_),
    .B1(_07394_),
    .X(_07441_));
 sky130_fd_sc_hd__o211ai_1 _14270_ (.A1(_07432_),
    .A2(_07435_),
    .B1(_07438_),
    .C1(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__nand2_1 _14271_ (.A(_07432_),
    .B(_07435_),
    .Y(_07443_));
 sky130_fd_sc_hd__a21oi_1 _14272_ (.A1(_07442_),
    .A2(_07443_),
    .B1(_07421_),
    .Y(_07444_));
 sky130_fd_sc_hd__or2_1 _14273_ (.A(_07273_),
    .B(_07278_),
    .X(_07445_));
 sky130_fd_sc_hd__nand2_1 _14274_ (.A(_07279_),
    .B(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__clkbuf_4 _14275_ (.A(_07446_),
    .X(_07447_));
 sky130_fd_sc_hd__or2_1 _14276_ (.A(_07338_),
    .B(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__nor2_1 _14277_ (.A(_07414_),
    .B(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__o22ai_1 _14278_ (.A1(_07335_),
    .A2(_07416_),
    .B1(_07413_),
    .B2(_07338_),
    .Y(_07450_));
 sky130_fd_sc_hd__o31a_1 _14279_ (.A1(_07338_),
    .A2(_07416_),
    .A3(_07414_),
    .B1(_07450_),
    .X(_07451_));
 sky130_fd_sc_hd__nand2_1 _14280_ (.A(_07449_),
    .B(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__clkbuf_4 _14281_ (.A(_06916_),
    .X(_07453_));
 sky130_fd_sc_hd__nor2_2 _14282_ (.A(_07453_),
    .B(_07411_),
    .Y(_07454_));
 sky130_fd_sc_hd__clkbuf_4 _14283_ (.A(_06943_),
    .X(_07455_));
 sky130_fd_sc_hd__a2bb2o_1 _14284_ (.A1_N(_07455_),
    .A2_N(_07411_),
    .B1(_07433_),
    .B2(_06919_),
    .X(_07456_));
 sky130_fd_sc_hd__and2_1 _14285_ (.A(_07056_),
    .B(_07419_),
    .X(_07457_));
 sky130_fd_sc_hd__xor2_2 _14286_ (.A(_07426_),
    .B(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__nand2_1 _14287_ (.A(_07454_),
    .B(_07456_),
    .Y(_07459_));
 sky130_fd_sc_hd__xor2_1 _14288_ (.A(_07459_),
    .B(_07458_),
    .X(_07460_));
 sky130_fd_sc_hd__nor2_1 _14289_ (.A(_07427_),
    .B(_07416_),
    .Y(_07461_));
 sky130_fd_sc_hd__and2_1 _14290_ (.A(_07288_),
    .B(_07419_),
    .X(_07462_));
 sky130_fd_sc_hd__xnor2_1 _14291_ (.A(_07423_),
    .B(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__and3_1 _14292_ (.A(_07098_),
    .B(_07425_),
    .C(_07419_),
    .X(_07464_));
 sky130_fd_sc_hd__a21oi_1 _14293_ (.A1(_07461_),
    .A2(_07463_),
    .B1(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__nor2_1 _14294_ (.A(_07460_),
    .B(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__a31o_1 _14295_ (.A1(_07454_),
    .A2(_07456_),
    .A3(_07458_),
    .B1(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__nand2_1 _14296_ (.A(_07414_),
    .B(_07417_),
    .Y(_07468_));
 sky130_fd_sc_hd__xnor2_1 _14297_ (.A(_07420_),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__inv_2 _14298_ (.A(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__xnor2_1 _14299_ (.A(_07467_),
    .B(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nand2_1 _14300_ (.A(_07467_),
    .B(_07470_),
    .Y(_07472_));
 sky130_fd_sc_hd__o21ai_1 _14301_ (.A1(_07452_),
    .A2(_07471_),
    .B1(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__xnor2_1 _14302_ (.A(_07438_),
    .B(_07441_),
    .Y(_07474_));
 sky130_fd_sc_hd__xor2_1 _14303_ (.A(_07452_),
    .B(_07471_),
    .X(_07475_));
 sky130_fd_sc_hd__inv_2 _14304_ (.A(_07433_),
    .Y(_07476_));
 sky130_fd_sc_hd__nor2_1 _14305_ (.A(_07455_),
    .B(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__or3_1 _14306_ (.A(_07437_),
    .B(_07454_),
    .C(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__xor2_1 _14307_ (.A(_07460_),
    .B(_07465_),
    .X(_07479_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(_07478_),
    .B(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__nor2_1 _14309_ (.A(_07426_),
    .B(_07428_),
    .Y(_07481_));
 sky130_fd_sc_hd__nor2_1 _14310_ (.A(_07457_),
    .B(_07429_),
    .Y(_07482_));
 sky130_fd_sc_hd__o21a_1 _14311_ (.A1(_07481_),
    .A2(_07482_),
    .B1(_07424_),
    .X(_07483_));
 sky130_fd_sc_hd__o2bb2a_1 _14312_ (.A1_N(_06975_),
    .A2_N(_07411_),
    .B1(_07483_),
    .B2(_07394_),
    .X(_07484_));
 sky130_fd_sc_hd__nor2_1 _14313_ (.A(_07480_),
    .B(_07484_),
    .Y(_07485_));
 sky130_fd_sc_hd__and2_1 _14314_ (.A(_07480_),
    .B(_07484_),
    .X(_07486_));
 sky130_fd_sc_hd__nor2_1 _14315_ (.A(_07485_),
    .B(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__a21oi_1 _14316_ (.A1(_07475_),
    .A2(_07487_),
    .B1(_07485_),
    .Y(_07488_));
 sky130_fd_sc_hd__nor2_1 _14317_ (.A(_07474_),
    .B(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__and2_1 _14318_ (.A(_07474_),
    .B(_07488_),
    .X(_07490_));
 sky130_fd_sc_hd__nor2_1 _14319_ (.A(_07489_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__a21oi_1 _14320_ (.A1(_07473_),
    .A2(_07491_),
    .B1(_07489_),
    .Y(_07492_));
 sky130_fd_sc_hd__or2_1 _14321_ (.A(_07444_),
    .B(_07492_),
    .X(_07493_));
 sky130_fd_sc_hd__mux2_1 _14322_ (.A0(_07430_),
    .A1(_07427_),
    .S(_07411_),
    .X(_07494_));
 sky130_fd_sc_hd__o21a_1 _14323_ (.A1(_07432_),
    .A2(_07435_),
    .B1(_07431_),
    .X(_07495_));
 sky130_fd_sc_hd__and2b_1 _14324_ (.A_N(_07494_),
    .B(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__inv_2 _14325_ (.A(_07442_),
    .Y(_07497_));
 sky130_fd_sc_hd__nor2_1 _14326_ (.A(_07497_),
    .B(_07496_),
    .Y(_07498_));
 sky130_fd_sc_hd__a31o_1 _14327_ (.A1(_07438_),
    .A2(_07441_),
    .A3(_07496_),
    .B1(_07498_),
    .X(_07499_));
 sky130_fd_sc_hd__nor2_1 _14328_ (.A(_07493_),
    .B(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__mux2_1 _14329_ (.A0(_07063_),
    .A1(_07427_),
    .S(_07411_),
    .X(_07501_));
 sky130_fd_sc_hd__or2_1 _14330_ (.A(_07430_),
    .B(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__a2bb2o_1 _14331_ (.A1_N(_07495_),
    .A2_N(_07502_),
    .B1(_07496_),
    .B2(_07497_),
    .X(_07503_));
 sky130_fd_sc_hd__a21oi_2 _14332_ (.A1(_07495_),
    .A2(_07502_),
    .B1(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__xor2_2 _14333_ (.A(_07500_),
    .B(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__xnor2_1 _14334_ (.A(_07473_),
    .B(_07491_),
    .Y(_07506_));
 sky130_fd_sc_hd__and2_1 _14335_ (.A(_07274_),
    .B(_07277_),
    .X(_07507_));
 sky130_fd_sc_hd__or2_1 _14336_ (.A(_07278_),
    .B(_07507_),
    .X(_07508_));
 sky130_fd_sc_hd__buf_2 _14337_ (.A(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__or2_1 _14338_ (.A(_07335_),
    .B(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__nor2_1 _14339_ (.A(_07448_),
    .B(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__and2_1 _14340_ (.A(_07414_),
    .B(_07448_),
    .X(_07512_));
 sky130_fd_sc_hd__nor2_1 _14341_ (.A(_07449_),
    .B(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__xnor2_1 _14342_ (.A(_07449_),
    .B(_07451_),
    .Y(_07514_));
 sky130_fd_sc_hd__o2bb2a_1 _14343_ (.A1_N(_07098_),
    .A2_N(_07419_),
    .B1(_07416_),
    .B2(_07422_),
    .X(_07515_));
 sky130_fd_sc_hd__nor2_1 _14344_ (.A(_07427_),
    .B(_07413_),
    .Y(_07516_));
 sky130_fd_sc_hd__nor2b_1 _14345_ (.A(_07515_),
    .B_N(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__or3_1 _14346_ (.A(_06943_),
    .B(_07236_),
    .C(_07409_),
    .X(_07518_));
 sky130_fd_sc_hd__a21oi_1 _14347_ (.A1(_07455_),
    .A2(_07236_),
    .B1(_07409_),
    .Y(_07519_));
 sky130_fd_sc_hd__and2_1 _14348_ (.A(_07518_),
    .B(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__nand2_1 _14349_ (.A(_07454_),
    .B(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__xnor2_1 _14350_ (.A(_07461_),
    .B(_07463_),
    .Y(_07522_));
 sky130_fd_sc_hd__nand3_1 _14351_ (.A(_07518_),
    .B(_07521_),
    .C(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__a21oi_1 _14352_ (.A1(_07518_),
    .A2(_07521_),
    .B1(_07522_),
    .Y(_07524_));
 sky130_fd_sc_hd__a21oi_1 _14353_ (.A1(_07517_),
    .A2(_07523_),
    .B1(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__xor2_1 _14354_ (.A(_07514_),
    .B(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__nor2_1 _14355_ (.A(_07514_),
    .B(_07525_),
    .Y(_07527_));
 sky130_fd_sc_hd__a31o_1 _14356_ (.A1(_07511_),
    .A2(_07513_),
    .A3(_07526_),
    .B1(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__xnor2_1 _14357_ (.A(_07475_),
    .B(_07487_),
    .Y(_07529_));
 sky130_fd_sc_hd__nand2_1 _14358_ (.A(_07511_),
    .B(_07513_),
    .Y(_07530_));
 sky130_fd_sc_hd__xnor2_1 _14359_ (.A(_07530_),
    .B(_07526_),
    .Y(_07531_));
 sky130_fd_sc_hd__xor2_1 _14360_ (.A(_07454_),
    .B(_07456_),
    .X(_07532_));
 sky130_fd_sc_hd__and2b_1 _14361_ (.A_N(_07524_),
    .B(_07523_),
    .X(_07533_));
 sky130_fd_sc_hd__xor2_2 _14362_ (.A(_07517_),
    .B(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__xor2_1 _14363_ (.A(_07478_),
    .B(_07479_),
    .X(_07535_));
 sky130_fd_sc_hd__and3_1 _14364_ (.A(_07532_),
    .B(_07534_),
    .C(_07535_),
    .X(_07536_));
 sky130_fd_sc_hd__a21oi_1 _14365_ (.A1(_07532_),
    .A2(_07534_),
    .B1(_07535_),
    .Y(_07537_));
 sky130_fd_sc_hd__nor2_1 _14366_ (.A(_07536_),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__a21oi_1 _14367_ (.A1(_07531_),
    .A2(_07538_),
    .B1(_07536_),
    .Y(_07539_));
 sky130_fd_sc_hd__nor2_1 _14368_ (.A(_07529_),
    .B(_07539_),
    .Y(_07540_));
 sky130_fd_sc_hd__and2_1 _14369_ (.A(_07529_),
    .B(_07539_),
    .X(_07541_));
 sky130_fd_sc_hd__nor2_1 _14370_ (.A(_07540_),
    .B(_07541_),
    .Y(_07542_));
 sky130_fd_sc_hd__a21oi_1 _14371_ (.A1(_07528_),
    .A2(_07542_),
    .B1(_07540_),
    .Y(_07543_));
 sky130_fd_sc_hd__nor2_1 _14372_ (.A(_07506_),
    .B(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__nand2_1 _14373_ (.A(_07444_),
    .B(_07492_),
    .Y(_07545_));
 sky130_fd_sc_hd__and2_1 _14374_ (.A(_07493_),
    .B(_07545_),
    .X(_07546_));
 sky130_fd_sc_hd__and2_1 _14375_ (.A(_07544_),
    .B(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__and2_1 _14376_ (.A(_07493_),
    .B(_07499_),
    .X(_07548_));
 sky130_fd_sc_hd__nor2_1 _14377_ (.A(_07500_),
    .B(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__and2_1 _14378_ (.A(_07547_),
    .B(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__nor2_1 _14379_ (.A(_07547_),
    .B(_07549_),
    .Y(_07551_));
 sky130_fd_sc_hd__nor2_1 _14380_ (.A(_07550_),
    .B(_07551_),
    .Y(_07552_));
 sky130_fd_sc_hd__inv_2 _14381_ (.A(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__nor2_1 _14382_ (.A(_07544_),
    .B(_07546_),
    .Y(_07554_));
 sky130_fd_sc_hd__nor2_1 _14383_ (.A(_07547_),
    .B(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__xnor2_2 _14384_ (.A(_07528_),
    .B(_07542_),
    .Y(_07556_));
 sky130_fd_sc_hd__xnor2_1 _14385_ (.A(_07531_),
    .B(_07538_),
    .Y(_07557_));
 sky130_fd_sc_hd__o22a_1 _14386_ (.A1(_07335_),
    .A2(_07447_),
    .B1(_07509_),
    .B2(_07338_),
    .X(_07558_));
 sky130_fd_sc_hd__nor2_1 _14387_ (.A(_07511_),
    .B(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__and2_1 _14388_ (.A(_07275_),
    .B(_07276_),
    .X(_07560_));
 sky130_fd_sc_hd__nor2_2 _14389_ (.A(_07277_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__nor2_1 _14390_ (.A(_07338_),
    .B(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__and2b_1 _14391_ (.A_N(_07510_),
    .B(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__o21ai_1 _14392_ (.A1(_07437_),
    .A2(_07559_),
    .B1(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__xnor2_1 _14393_ (.A(_07511_),
    .B(_07513_),
    .Y(_07565_));
 sky130_fd_sc_hd__and2_1 _14394_ (.A(_06975_),
    .B(_07419_),
    .X(_07566_));
 sky130_fd_sc_hd__a21bo_1 _14395_ (.A1(_07519_),
    .A2(_07566_),
    .B1_N(_07518_),
    .X(_07567_));
 sky130_fd_sc_hd__and2b_1 _14396_ (.A_N(_07516_),
    .B(_07515_),
    .X(_07568_));
 sky130_fd_sc_hd__nor2_1 _14397_ (.A(_07517_),
    .B(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__xnor2_1 _14398_ (.A(_07567_),
    .B(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__or2_1 _14399_ (.A(_07422_),
    .B(_07412_),
    .X(_07571_));
 sky130_fd_sc_hd__nor2_1 _14400_ (.A(_07152_),
    .B(_07415_),
    .Y(_07572_));
 sky130_fd_sc_hd__xnor2_1 _14401_ (.A(_07571_),
    .B(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__or3b_1 _14402_ (.A(_07427_),
    .B(_07447_),
    .C_N(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__o31a_1 _14403_ (.A1(_07152_),
    .A2(_07416_),
    .A3(_07571_),
    .B1(_07574_),
    .X(_07575_));
 sky130_fd_sc_hd__nor2_1 _14404_ (.A(_07570_),
    .B(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__a21oi_1 _14405_ (.A1(_07567_),
    .A2(_07569_),
    .B1(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__xor2_1 _14406_ (.A(_07565_),
    .B(_07577_),
    .X(_07578_));
 sky130_fd_sc_hd__xnor2_1 _14407_ (.A(_07564_),
    .B(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__xnor2_1 _14408_ (.A(_07532_),
    .B(_07534_),
    .Y(_07580_));
 sky130_fd_sc_hd__and2_1 _14409_ (.A(_07570_),
    .B(_07575_),
    .X(_07581_));
 sky130_fd_sc_hd__nor2_1 _14410_ (.A(_07576_),
    .B(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__or2_1 _14411_ (.A(_07454_),
    .B(_07520_),
    .X(_07583_));
 sky130_fd_sc_hd__clkbuf_4 _14412_ (.A(_06925_),
    .X(_07584_));
 sky130_fd_sc_hd__nor2_1 _14413_ (.A(_07584_),
    .B(_07476_),
    .Y(_07585_));
 sky130_fd_sc_hd__a211o_1 _14414_ (.A1(_07521_),
    .A2(_07583_),
    .B1(_07585_),
    .C1(_07437_),
    .X(_07586_));
 sky130_fd_sc_hd__xor2_1 _14415_ (.A(_07520_),
    .B(_07566_),
    .X(_07587_));
 sky130_fd_sc_hd__nor2_1 _14416_ (.A(_07584_),
    .B(_07410_),
    .Y(_07588_));
 sky130_fd_sc_hd__a21o_1 _14417_ (.A1(_06927_),
    .A2(_07433_),
    .B1(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__and3b_1 _14418_ (.A_N(_07410_),
    .B(_06904_),
    .C(_06927_),
    .X(_07590_));
 sky130_fd_sc_hd__a21o_1 _14419_ (.A1(_07587_),
    .A2(_07589_),
    .B1(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__xor2_1 _14420_ (.A(_07586_),
    .B(_07591_),
    .X(_07592_));
 sky130_fd_sc_hd__and2_1 _14421_ (.A(_07586_),
    .B(_07591_),
    .X(_07593_));
 sky130_fd_sc_hd__a21oi_1 _14422_ (.A1(_07582_),
    .A2(_07592_),
    .B1(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__nand2_1 _14423_ (.A(_07580_),
    .B(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__nor2_1 _14424_ (.A(_07580_),
    .B(_07594_),
    .Y(_07596_));
 sky130_fd_sc_hd__a21oi_1 _14425_ (.A1(_07579_),
    .A2(_07595_),
    .B1(_07596_),
    .Y(_07597_));
 sky130_fd_sc_hd__xnor2_1 _14426_ (.A(_07557_),
    .B(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__or2b_1 _14427_ (.A(_07564_),
    .B_N(_07578_),
    .X(_07599_));
 sky130_fd_sc_hd__o21ai_1 _14428_ (.A1(_07565_),
    .A2(_07577_),
    .B1(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__or2b_1 _14429_ (.A(_07598_),
    .B_N(_07600_),
    .X(_07601_));
 sky130_fd_sc_hd__o21a_1 _14430_ (.A1(_07557_),
    .A2(_07597_),
    .B1(_07601_),
    .X(_07602_));
 sky130_fd_sc_hd__nor2_1 _14431_ (.A(_07556_),
    .B(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__and2_1 _14432_ (.A(_07506_),
    .B(_07543_),
    .X(_07604_));
 sky130_fd_sc_hd__nor2_1 _14433_ (.A(_07544_),
    .B(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__and2_1 _14434_ (.A(_07603_),
    .B(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__xor2_1 _14435_ (.A(_07555_),
    .B(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__inv_2 _14436_ (.A(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__xor2_1 _14437_ (.A(_07603_),
    .B(_07605_),
    .X(_07609_));
 sky130_fd_sc_hd__xor2_1 _14438_ (.A(_07600_),
    .B(_07598_),
    .X(_07610_));
 sky130_fd_sc_hd__buf_2 _14439_ (.A(_07276_),
    .X(_07611_));
 sky130_fd_sc_hd__or2_1 _14440_ (.A(_07335_),
    .B(_07611_),
    .X(_07612_));
 sky130_fd_sc_hd__inv_2 _14441_ (.A(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__nand2_1 _14442_ (.A(_07562_),
    .B(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__or2_1 _14443_ (.A(_07563_),
    .B(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__or3_1 _14444_ (.A(_07437_),
    .B(_07563_),
    .C(_07559_),
    .X(_07616_));
 sky130_fd_sc_hd__nand2_1 _14445_ (.A(_07564_),
    .B(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__nor2_1 _14446_ (.A(_07236_),
    .B(_07409_),
    .Y(_07618_));
 sky130_fd_sc_hd__and2b_1 _14447_ (.A_N(_06943_),
    .B(_07418_),
    .X(_07619_));
 sky130_fd_sc_hd__xnor2_2 _14448_ (.A(_07618_),
    .B(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__nand2_1 _14449_ (.A(_07618_),
    .B(_07619_),
    .Y(_07621_));
 sky130_fd_sc_hd__o31ai_4 _14450_ (.A1(_07453_),
    .A2(_07416_),
    .A3(_07620_),
    .B1(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__o21bai_1 _14451_ (.A1(_07427_),
    .A2(_07447_),
    .B1_N(_07573_),
    .Y(_07623_));
 sky130_fd_sc_hd__and2_1 _14452_ (.A(_07574_),
    .B(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__xnor2_2 _14453_ (.A(_07622_),
    .B(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__or2_1 _14454_ (.A(_06860_),
    .B(_07508_),
    .X(_07626_));
 sky130_fd_sc_hd__nor2_1 _14455_ (.A(_07152_),
    .B(_07412_),
    .Y(_07627_));
 sky130_fd_sc_hd__nor2_1 _14456_ (.A(_07422_),
    .B(_07446_),
    .Y(_07628_));
 sky130_fd_sc_hd__nand2_1 _14457_ (.A(_07627_),
    .B(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__or2_1 _14458_ (.A(_07627_),
    .B(_07628_),
    .X(_07630_));
 sky130_fd_sc_hd__nand2_1 _14459_ (.A(_07629_),
    .B(_07630_),
    .Y(_07631_));
 sky130_fd_sc_hd__o21a_1 _14460_ (.A1(_07626_),
    .A2(_07631_),
    .B1(_07629_),
    .X(_07632_));
 sky130_fd_sc_hd__nand2_1 _14461_ (.A(_07622_),
    .B(_07624_),
    .Y(_07633_));
 sky130_fd_sc_hd__o21a_1 _14462_ (.A1(_07625_),
    .A2(_07632_),
    .B1(_07633_),
    .X(_07634_));
 sky130_fd_sc_hd__or2_1 _14463_ (.A(_07617_),
    .B(_07634_),
    .X(_07635_));
 sky130_fd_sc_hd__nand2_1 _14464_ (.A(_07617_),
    .B(_07634_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand2_1 _14465_ (.A(_07635_),
    .B(_07636_),
    .Y(_07637_));
 sky130_fd_sc_hd__o21ai_1 _14466_ (.A1(_07615_),
    .A2(_07637_),
    .B1(_07635_),
    .Y(_07638_));
 sky130_fd_sc_hd__and2b_1 _14467_ (.A_N(_07596_),
    .B(_07595_),
    .X(_07639_));
 sky130_fd_sc_hd__xnor2_1 _14468_ (.A(_07579_),
    .B(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__xor2_1 _14469_ (.A(_07615_),
    .B(_07637_),
    .X(_07641_));
 sky130_fd_sc_hd__xnor2_1 _14470_ (.A(_07582_),
    .B(_07592_),
    .Y(_07642_));
 sky130_fd_sc_hd__or2b_1 _14471_ (.A(_07590_),
    .B_N(_07589_),
    .X(_07643_));
 sky130_fd_sc_hd__xor2_1 _14472_ (.A(_07587_),
    .B(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__nor2_1 _14473_ (.A(_07139_),
    .B(_07410_),
    .Y(_07645_));
 sky130_fd_sc_hd__a211oi_1 _14474_ (.A1(_07055_),
    .A2(_07433_),
    .B1(_07588_),
    .C1(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__or2_1 _14475_ (.A(_06869_),
    .B(_07410_),
    .X(_07647_));
 sky130_fd_sc_hd__or3_1 _14476_ (.A(_06844_),
    .B(_06925_),
    .C(_07409_),
    .X(_07648_));
 sky130_fd_sc_hd__a21oi_1 _14477_ (.A1(_07647_),
    .A2(_07648_),
    .B1(_07590_),
    .Y(_07649_));
 sky130_fd_sc_hd__nor2_1 _14478_ (.A(_07453_),
    .B(_07416_),
    .Y(_07650_));
 sky130_fd_sc_hd__xnor2_1 _14479_ (.A(_07620_),
    .B(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__nor2_1 _14480_ (.A(_07649_),
    .B(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__xor2_2 _14481_ (.A(_07625_),
    .B(_07632_),
    .X(_07653_));
 sky130_fd_sc_hd__nor2_1 _14482_ (.A(_07646_),
    .B(_07649_),
    .Y(_07654_));
 sky130_fd_sc_hd__a21o_1 _14483_ (.A1(_07651_),
    .A2(_07654_),
    .B1(_07649_),
    .X(_07655_));
 sky130_fd_sc_hd__xnor2_1 _14484_ (.A(_07644_),
    .B(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__nand2_1 _14485_ (.A(_07653_),
    .B(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__o31a_1 _14486_ (.A1(_07644_),
    .A2(_07646_),
    .A3(_07652_),
    .B1(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__xor2_1 _14487_ (.A(_07642_),
    .B(_07658_),
    .X(_07659_));
 sky130_fd_sc_hd__nor2_1 _14488_ (.A(_07642_),
    .B(_07658_),
    .Y(_07660_));
 sky130_fd_sc_hd__a21oi_1 _14489_ (.A1(_07641_),
    .A2(_07659_),
    .B1(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__xor2_1 _14490_ (.A(_07640_),
    .B(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__nor2_1 _14491_ (.A(_07640_),
    .B(_07661_),
    .Y(_07663_));
 sky130_fd_sc_hd__a21oi_1 _14492_ (.A1(_07638_),
    .A2(_07662_),
    .B1(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__nor2_1 _14493_ (.A(_07610_),
    .B(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__xor2_2 _14494_ (.A(_07556_),
    .B(_07602_),
    .X(_07666_));
 sky130_fd_sc_hd__and2_1 _14495_ (.A(_07665_),
    .B(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__and2_1 _14496_ (.A(_07609_),
    .B(_07667_),
    .X(_07668_));
 sky130_fd_sc_hd__nor2_1 _14497_ (.A(_07609_),
    .B(_07667_),
    .Y(_07669_));
 sky130_fd_sc_hd__nor2_1 _14498_ (.A(_07668_),
    .B(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__inv_2 _14499_ (.A(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__xnor2_1 _14500_ (.A(_07638_),
    .B(_07662_),
    .Y(_07672_));
 sky130_fd_sc_hd__or2_1 _14501_ (.A(_07236_),
    .B(_07415_),
    .X(_07673_));
 sky130_fd_sc_hd__or3b_1 _14502_ (.A(_07673_),
    .B(_07455_),
    .C_N(_07418_),
    .X(_07674_));
 sky130_fd_sc_hd__nor2_1 _14503_ (.A(_07455_),
    .B(_07415_),
    .Y(_07675_));
 sky130_fd_sc_hd__a21o_1 _14504_ (.A1(_06919_),
    .A2(_07418_),
    .B1(_07675_),
    .X(_07676_));
 sky130_fd_sc_hd__nor2_1 _14505_ (.A(_07453_),
    .B(_07413_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand3_1 _14506_ (.A(_07674_),
    .B(_07676_),
    .C(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__xnor2_1 _14507_ (.A(_07626_),
    .B(_07631_),
    .Y(_07679_));
 sky130_fd_sc_hd__a21oi_1 _14508_ (.A1(_07674_),
    .A2(_07678_),
    .B1(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__and3_1 _14509_ (.A(_07674_),
    .B(_07678_),
    .C(_07679_),
    .X(_07681_));
 sky130_fd_sc_hd__or2_1 _14510_ (.A(_07680_),
    .B(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__or2_1 _14511_ (.A(_07152_),
    .B(_07508_),
    .X(_07683_));
 sky130_fd_sc_hd__inv_2 _14512_ (.A(_07683_),
    .Y(_07684_));
 sky130_fd_sc_hd__or2_1 _14513_ (.A(_07427_),
    .B(_07561_),
    .X(_07685_));
 sky130_fd_sc_hd__o22a_1 _14514_ (.A1(_07152_),
    .A2(_07447_),
    .B1(_07508_),
    .B2(_07422_),
    .X(_07686_));
 sky130_fd_sc_hd__a21o_1 _14515_ (.A1(_07628_),
    .A2(_07684_),
    .B1(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__o2bb2a_1 _14516_ (.A1_N(_07628_),
    .A2_N(_07684_),
    .B1(_07685_),
    .B2(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__nor2_1 _14517_ (.A(_07682_),
    .B(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__a21boi_1 _14518_ (.A1(_07562_),
    .A2(_07612_),
    .B1_N(_07510_),
    .Y(_07690_));
 sky130_fd_sc_hd__a21oi_1 _14519_ (.A1(_07563_),
    .A2(_07614_),
    .B1(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__o21a_1 _14520_ (.A1(_07680_),
    .A2(_07689_),
    .B1(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__xnor2_1 _14521_ (.A(_07641_),
    .B(_07659_),
    .Y(_07693_));
 sky130_fd_sc_hd__nor3_1 _14522_ (.A(_07680_),
    .B(_07689_),
    .C(_07691_),
    .Y(_07694_));
 sky130_fd_sc_hd__nor2_1 _14523_ (.A(_07692_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__xnor2_2 _14524_ (.A(_07653_),
    .B(_07656_),
    .Y(_07696_));
 sky130_fd_sc_hd__xor2_1 _14525_ (.A(_07682_),
    .B(_07688_),
    .X(_07697_));
 sky130_fd_sc_hd__a21o_1 _14526_ (.A1(_07674_),
    .A2(_07676_),
    .B1(_07677_),
    .X(_07698_));
 sky130_fd_sc_hd__and2_1 _14527_ (.A(_07678_),
    .B(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__a21oi_1 _14528_ (.A1(_06844_),
    .A2(_07584_),
    .B1(_07410_),
    .Y(_07700_));
 sky130_fd_sc_hd__nand2_1 _14529_ (.A(_07648_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__nand2_1 _14530_ (.A(_06904_),
    .B(_07419_),
    .Y(_07702_));
 sky130_fd_sc_hd__o31ai_2 _14531_ (.A1(_06844_),
    .A2(_07410_),
    .A3(_07702_),
    .B1(_07647_),
    .Y(_07703_));
 sky130_fd_sc_hd__xnor2_2 _14532_ (.A(_07701_),
    .B(_07703_),
    .Y(_07704_));
 sky130_fd_sc_hd__or2b_1 _14533_ (.A(_07701_),
    .B_N(_07703_),
    .X(_07705_));
 sky130_fd_sc_hd__a21bo_1 _14534_ (.A1(_07699_),
    .A2(_07704_),
    .B1_N(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__xnor2_1 _14535_ (.A(_07651_),
    .B(_07654_),
    .Y(_07707_));
 sky130_fd_sc_hd__xnor2_1 _14536_ (.A(_07706_),
    .B(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__nand2_1 _14537_ (.A(_07699_),
    .B(_07704_),
    .Y(_07709_));
 sky130_fd_sc_hd__a21oi_1 _14538_ (.A1(_07705_),
    .A2(_07709_),
    .B1(_07707_),
    .Y(_07710_));
 sky130_fd_sc_hd__a21oi_1 _14539_ (.A1(_07697_),
    .A2(_07708_),
    .B1(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__xor2_1 _14540_ (.A(_07696_),
    .B(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__nor2_1 _14541_ (.A(_07696_),
    .B(_07711_),
    .Y(_07713_));
 sky130_fd_sc_hd__a21oi_1 _14542_ (.A1(_07695_),
    .A2(_07712_),
    .B1(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__xor2_1 _14543_ (.A(_07693_),
    .B(_07714_),
    .X(_07715_));
 sky130_fd_sc_hd__nor2_1 _14544_ (.A(_07693_),
    .B(_07714_),
    .Y(_07716_));
 sky130_fd_sc_hd__a21oi_1 _14545_ (.A1(_07692_),
    .A2(_07715_),
    .B1(_07716_),
    .Y(_07717_));
 sky130_fd_sc_hd__nor2_1 _14546_ (.A(_07672_),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__and2_1 _14547_ (.A(_07610_),
    .B(_07664_),
    .X(_07719_));
 sky130_fd_sc_hd__nor2_1 _14548_ (.A(_07665_),
    .B(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__and2_1 _14549_ (.A(_07718_),
    .B(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__xnor2_1 _14550_ (.A(_07692_),
    .B(_07715_),
    .Y(_07722_));
 sky130_fd_sc_hd__nor2_1 _14551_ (.A(_07236_),
    .B(_07413_),
    .Y(_07723_));
 sky130_fd_sc_hd__nand2_1 _14552_ (.A(_07675_),
    .B(_07723_),
    .Y(_07724_));
 sky130_fd_sc_hd__nor2_1 _14553_ (.A(_07455_),
    .B(_07413_),
    .Y(_07725_));
 sky130_fd_sc_hd__xnor2_1 _14554_ (.A(_07673_),
    .B(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__nor2_1 _14555_ (.A(_07453_),
    .B(_07447_),
    .Y(_07727_));
 sky130_fd_sc_hd__nand2_1 _14556_ (.A(_07726_),
    .B(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__xnor2_1 _14557_ (.A(_07685_),
    .B(_07687_),
    .Y(_07729_));
 sky130_fd_sc_hd__a21o_1 _14558_ (.A1(_07724_),
    .A2(_07728_),
    .B1(_07729_),
    .X(_07730_));
 sky130_fd_sc_hd__nand3_1 _14559_ (.A(_07724_),
    .B(_07728_),
    .C(_07729_),
    .Y(_07731_));
 sky130_fd_sc_hd__nand2_1 _14560_ (.A(_07730_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__clkbuf_4 _14561_ (.A(_07561_),
    .X(_07733_));
 sky130_fd_sc_hd__nor2_1 _14562_ (.A(_07422_),
    .B(_07509_),
    .Y(_07734_));
 sky130_fd_sc_hd__nor2_1 _14563_ (.A(_07152_),
    .B(_07561_),
    .Y(_07735_));
 sky130_fd_sc_hd__o21a_1 _14564_ (.A1(_07422_),
    .A2(_07561_),
    .B1(_07683_),
    .X(_07736_));
 sky130_fd_sc_hd__a21oi_1 _14565_ (.A1(_07734_),
    .A2(_07735_),
    .B1(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__or3b_1 _14566_ (.A(_07427_),
    .B(_07611_),
    .C_N(_07737_),
    .X(_07738_));
 sky130_fd_sc_hd__o31a_1 _14567_ (.A1(_07422_),
    .A2(_07733_),
    .A3(_07683_),
    .B1(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__or2_1 _14568_ (.A(_07732_),
    .B(_07739_),
    .X(_07740_));
 sky130_fd_sc_hd__o22a_1 _14569_ (.A1(_07338_),
    .A2(_07611_),
    .B1(_07733_),
    .B2(_07335_),
    .X(_07741_));
 sky130_fd_sc_hd__a21o_1 _14570_ (.A1(_07562_),
    .A2(_07613_),
    .B1(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__a21oi_2 _14571_ (.A1(_07730_),
    .A2(_07740_),
    .B1(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__xnor2_1 _14572_ (.A(_07695_),
    .B(_07712_),
    .Y(_07744_));
 sky130_fd_sc_hd__and3_1 _14573_ (.A(_07730_),
    .B(_07740_),
    .C(_07742_),
    .X(_07745_));
 sky130_fd_sc_hd__nor2_1 _14574_ (.A(_07743_),
    .B(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__xor2_1 _14575_ (.A(_07697_),
    .B(_07708_),
    .X(_07747_));
 sky130_fd_sc_hd__xor2_1 _14576_ (.A(_07732_),
    .B(_07739_),
    .X(_07748_));
 sky130_fd_sc_hd__xnor2_1 _14577_ (.A(_07699_),
    .B(_07704_),
    .Y(_07749_));
 sky130_fd_sc_hd__or2_1 _14578_ (.A(_07726_),
    .B(_07727_),
    .X(_07750_));
 sky130_fd_sc_hd__and2_1 _14579_ (.A(_07728_),
    .B(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__nor2_1 _14580_ (.A(_06844_),
    .B(_07410_),
    .Y(_07752_));
 sky130_fd_sc_hd__xnor2_1 _14581_ (.A(_07752_),
    .B(_07702_),
    .Y(_07753_));
 sky130_fd_sc_hd__nor2_1 _14582_ (.A(_07584_),
    .B(_07415_),
    .Y(_07754_));
 sky130_fd_sc_hd__a2bb2o_1 _14583_ (.A1_N(_06894_),
    .A2_N(_07410_),
    .B1(_07418_),
    .B2(_06927_),
    .X(_07755_));
 sky130_fd_sc_hd__or4b_1 _14584_ (.A(_06894_),
    .B(_07139_),
    .C(_07409_),
    .D_N(_07418_),
    .X(_07756_));
 sky130_fd_sc_hd__a21boi_1 _14585_ (.A1(_07754_),
    .A2(_07755_),
    .B1_N(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__xnor2_1 _14586_ (.A(_07753_),
    .B(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__and2b_1 _14587_ (.A_N(_07757_),
    .B(_07753_),
    .X(_07759_));
 sky130_fd_sc_hd__a21oi_1 _14588_ (.A1(_07751_),
    .A2(_07758_),
    .B1(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__xor2_1 _14589_ (.A(_07749_),
    .B(_07760_),
    .X(_07761_));
 sky130_fd_sc_hd__nor2_1 _14590_ (.A(_07749_),
    .B(_07760_),
    .Y(_07762_));
 sky130_fd_sc_hd__a21oi_1 _14591_ (.A1(_07748_),
    .A2(_07761_),
    .B1(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__xnor2_1 _14592_ (.A(_07747_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__or2b_1 _14593_ (.A(_07763_),
    .B_N(_07747_),
    .X(_07765_));
 sky130_fd_sc_hd__a21boi_1 _14594_ (.A1(_07746_),
    .A2(_07764_),
    .B1_N(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__xor2_1 _14595_ (.A(_07744_),
    .B(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__nor2_1 _14596_ (.A(_07744_),
    .B(_07766_),
    .Y(_07768_));
 sky130_fd_sc_hd__a21oi_1 _14597_ (.A1(_07743_),
    .A2(_07767_),
    .B1(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__nor2_1 _14598_ (.A(_07722_),
    .B(_07769_),
    .Y(_07770_));
 sky130_fd_sc_hd__xor2_1 _14599_ (.A(_07672_),
    .B(_07717_),
    .X(_07771_));
 sky130_fd_sc_hd__and2_1 _14600_ (.A(_07770_),
    .B(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__xnor2_1 _14601_ (.A(_07743_),
    .B(_07767_),
    .Y(_07773_));
 sky130_fd_sc_hd__nor2_1 _14602_ (.A(_07236_),
    .B(_07447_),
    .Y(_07774_));
 sky130_fd_sc_hd__nand2_1 _14603_ (.A(_07725_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__nor2_1 _14604_ (.A(_06943_),
    .B(_07446_),
    .Y(_07776_));
 sky130_fd_sc_hd__or2_1 _14605_ (.A(_07723_),
    .B(_07776_),
    .X(_07777_));
 sky130_fd_sc_hd__nand2_1 _14606_ (.A(_07775_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__or3_1 _14607_ (.A(_07453_),
    .B(_07509_),
    .C(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__o21bai_1 _14608_ (.A1(_07427_),
    .A2(_07611_),
    .B1_N(_07737_),
    .Y(_07780_));
 sky130_fd_sc_hd__nand2_1 _14609_ (.A(_07738_),
    .B(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__nand3_1 _14610_ (.A(_07775_),
    .B(_07779_),
    .C(_07781_),
    .Y(_07782_));
 sky130_fd_sc_hd__nor2_1 _14611_ (.A(_07422_),
    .B(_07611_),
    .Y(_07783_));
 sky130_fd_sc_hd__and2_1 _14612_ (.A(_07735_),
    .B(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__a21o_1 _14613_ (.A1(_07775_),
    .A2(_07779_),
    .B1(_07781_),
    .X(_07785_));
 sky130_fd_sc_hd__a21boi_1 _14614_ (.A1(_07782_),
    .A2(_07784_),
    .B1_N(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__nor2_1 _14615_ (.A(_07612_),
    .B(_07786_),
    .Y(_07787_));
 sky130_fd_sc_hd__xnor2_1 _14616_ (.A(_07746_),
    .B(_07764_),
    .Y(_07788_));
 sky130_fd_sc_hd__and2_1 _14617_ (.A(_07612_),
    .B(_07786_),
    .X(_07789_));
 sky130_fd_sc_hd__nor2_1 _14618_ (.A(_07787_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__xnor2_1 _14619_ (.A(_07748_),
    .B(_07761_),
    .Y(_07791_));
 sky130_fd_sc_hd__nand2_1 _14620_ (.A(_07785_),
    .B(_07782_),
    .Y(_07792_));
 sky130_fd_sc_hd__xnor2_1 _14621_ (.A(_07792_),
    .B(_07784_),
    .Y(_07793_));
 sky130_fd_sc_hd__xnor2_1 _14622_ (.A(_07751_),
    .B(_07758_),
    .Y(_07794_));
 sky130_fd_sc_hd__nor2_1 _14623_ (.A(_07453_),
    .B(_07509_),
    .Y(_07795_));
 sky130_fd_sc_hd__xnor2_1 _14624_ (.A(_07778_),
    .B(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__and3_1 _14625_ (.A(_07756_),
    .B(_07754_),
    .C(_07755_),
    .X(_07797_));
 sky130_fd_sc_hd__a21oi_1 _14626_ (.A1(_07756_),
    .A2(_07755_),
    .B1(_07754_),
    .Y(_07798_));
 sky130_fd_sc_hd__nor2_1 _14627_ (.A(_07584_),
    .B(_07413_),
    .Y(_07799_));
 sky130_fd_sc_hd__nor2_1 _14628_ (.A(_07139_),
    .B(_07415_),
    .Y(_07800_));
 sky130_fd_sc_hd__a21o_1 _14629_ (.A1(_07055_),
    .A2(_07419_),
    .B1(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__nand3_1 _14630_ (.A(_07055_),
    .B(_07419_),
    .C(_07800_),
    .Y(_07802_));
 sky130_fd_sc_hd__a21boi_1 _14631_ (.A1(_07799_),
    .A2(_07801_),
    .B1_N(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__o21ai_1 _14632_ (.A1(_07797_),
    .A2(_07798_),
    .B1(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__or3_1 _14633_ (.A(_07797_),
    .B(_07798_),
    .C(_07803_),
    .X(_07805_));
 sky130_fd_sc_hd__a21bo_1 _14634_ (.A1(_07796_),
    .A2(_07804_),
    .B1_N(_07805_),
    .X(_07806_));
 sky130_fd_sc_hd__xnor2_1 _14635_ (.A(_07794_),
    .B(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__or2b_1 _14636_ (.A(_07794_),
    .B_N(_07806_),
    .X(_07808_));
 sky130_fd_sc_hd__a21bo_1 _14637_ (.A1(_07793_),
    .A2(_07807_),
    .B1_N(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__xnor2_1 _14638_ (.A(_07791_),
    .B(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__or2b_1 _14639_ (.A(_07791_),
    .B_N(_07809_),
    .X(_07811_));
 sky130_fd_sc_hd__a21boi_1 _14640_ (.A1(_07790_),
    .A2(_07810_),
    .B1_N(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__xor2_1 _14641_ (.A(_07788_),
    .B(_07812_),
    .X(_07813_));
 sky130_fd_sc_hd__nor2_1 _14642_ (.A(_07788_),
    .B(_07812_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21oi_1 _14643_ (.A1(_07787_),
    .A2(_07813_),
    .B1(_07814_),
    .Y(_07815_));
 sky130_fd_sc_hd__nor2_1 _14644_ (.A(_07773_),
    .B(_07815_),
    .Y(_07816_));
 sky130_fd_sc_hd__xor2_1 _14645_ (.A(_07722_),
    .B(_07769_),
    .X(_07817_));
 sky130_fd_sc_hd__and2_1 _14646_ (.A(_07816_),
    .B(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__xor2_1 _14647_ (.A(_07773_),
    .B(_07815_),
    .X(_07819_));
 sky130_fd_sc_hd__nor2_1 _14648_ (.A(_07236_),
    .B(_07509_),
    .Y(_07820_));
 sky130_fd_sc_hd__nand2_1 _14649_ (.A(_07776_),
    .B(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__o21bai_1 _14650_ (.A1(_07455_),
    .A2(_07509_),
    .B1_N(_07774_),
    .Y(_07822_));
 sky130_fd_sc_hd__nand2_1 _14651_ (.A(_07821_),
    .B(_07822_),
    .Y(_07823_));
 sky130_fd_sc_hd__or3_1 _14652_ (.A(_07453_),
    .B(_07733_),
    .C(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__nor2_1 _14653_ (.A(_07735_),
    .B(_07783_),
    .Y(_07825_));
 sky130_fd_sc_hd__or2_1 _14654_ (.A(_07784_),
    .B(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__a21oi_2 _14655_ (.A1(_07821_),
    .A2(_07824_),
    .B1(_07826_),
    .Y(_07827_));
 sky130_fd_sc_hd__xnor2_1 _14656_ (.A(_07793_),
    .B(_07807_),
    .Y(_07828_));
 sky130_fd_sc_hd__and3_1 _14657_ (.A(_07805_),
    .B(_07796_),
    .C(_07804_),
    .X(_07829_));
 sky130_fd_sc_hd__a21oi_1 _14658_ (.A1(_07805_),
    .A2(_07804_),
    .B1(_07796_),
    .Y(_07830_));
 sky130_fd_sc_hd__nor2_1 _14659_ (.A(_07453_),
    .B(_07733_),
    .Y(_07831_));
 sky130_fd_sc_hd__xnor2_1 _14660_ (.A(_07823_),
    .B(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__nand3_1 _14661_ (.A(_07802_),
    .B(_07799_),
    .C(_07801_),
    .Y(_07833_));
 sky130_fd_sc_hd__a21o_1 _14662_ (.A1(_07802_),
    .A2(_07801_),
    .B1(_07799_),
    .X(_07834_));
 sky130_fd_sc_hd__nor2_1 _14663_ (.A(_06894_),
    .B(_07413_),
    .Y(_07835_));
 sky130_fd_sc_hd__nor2_1 _14664_ (.A(_07584_),
    .B(_07447_),
    .Y(_07836_));
 sky130_fd_sc_hd__or2_1 _14665_ (.A(_07139_),
    .B(_07413_),
    .X(_07837_));
 sky130_fd_sc_hd__o21a_1 _14666_ (.A1(_06894_),
    .A2(_07416_),
    .B1(_07837_),
    .X(_07838_));
 sky130_fd_sc_hd__a21oi_1 _14667_ (.A1(_07800_),
    .A2(_07835_),
    .B1(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__a22o_1 _14668_ (.A1(_07800_),
    .A2(_07835_),
    .B1(_07836_),
    .B2(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__a21o_1 _14669_ (.A1(_07833_),
    .A2(_07834_),
    .B1(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__and3_1 _14670_ (.A(_07833_),
    .B(_07834_),
    .C(_07840_),
    .X(_07842_));
 sky130_fd_sc_hd__a21oi_1 _14671_ (.A1(_07832_),
    .A2(_07841_),
    .B1(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__or3_1 _14672_ (.A(_07829_),
    .B(_07830_),
    .C(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__and3_1 _14673_ (.A(_07821_),
    .B(_07824_),
    .C(_07826_),
    .X(_07845_));
 sky130_fd_sc_hd__nor2_1 _14674_ (.A(_07827_),
    .B(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__o21ai_1 _14675_ (.A1(_07829_),
    .A2(_07830_),
    .B1(_07843_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand3_1 _14676_ (.A(_07844_),
    .B(_07846_),
    .C(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__and2_1 _14677_ (.A(_07844_),
    .B(_07848_),
    .X(_07849_));
 sky130_fd_sc_hd__nand2_1 _14678_ (.A(_07828_),
    .B(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__nor2_1 _14679_ (.A(_07828_),
    .B(_07849_),
    .Y(_07851_));
 sky130_fd_sc_hd__a21oi_1 _14680_ (.A1(_07827_),
    .A2(_07850_),
    .B1(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__xnor2_1 _14681_ (.A(_07790_),
    .B(_07810_),
    .Y(_07853_));
 sky130_fd_sc_hd__xor2_1 _14682_ (.A(_07787_),
    .B(_07813_),
    .X(_07854_));
 sky130_fd_sc_hd__nor3b_1 _14683_ (.A(_07852_),
    .B(_07853_),
    .C_N(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__and2_1 _14684_ (.A(_07819_),
    .B(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__xor2_1 _14685_ (.A(_07819_),
    .B(_07855_),
    .X(_07857_));
 sky130_fd_sc_hd__and2b_1 _14686_ (.A_N(_07851_),
    .B(_07850_),
    .X(_07858_));
 sky130_fd_sc_hd__xor2_1 _14687_ (.A(_07827_),
    .B(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__or2_1 _14688_ (.A(_07152_),
    .B(_07611_),
    .X(_07860_));
 sky130_fd_sc_hd__nor2_1 _14689_ (.A(_07455_),
    .B(_07733_),
    .Y(_07861_));
 sky130_fd_sc_hd__xnor2_1 _14690_ (.A(_07820_),
    .B(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__nor2_1 _14691_ (.A(_07453_),
    .B(_07611_),
    .Y(_07863_));
 sky130_fd_sc_hd__and2b_1 _14692_ (.A_N(_07862_),
    .B(_07863_),
    .X(_07864_));
 sky130_fd_sc_hd__a21oi_1 _14693_ (.A1(_07820_),
    .A2(_07861_),
    .B1(_07864_),
    .Y(_07865_));
 sky130_fd_sc_hd__nor2_1 _14694_ (.A(_07860_),
    .B(_07865_),
    .Y(_07866_));
 sky130_fd_sc_hd__a21o_1 _14695_ (.A1(_07844_),
    .A2(_07847_),
    .B1(_07846_),
    .X(_07867_));
 sky130_fd_sc_hd__xnor2_1 _14696_ (.A(_07836_),
    .B(_07839_),
    .Y(_07868_));
 sky130_fd_sc_hd__or2_1 _14697_ (.A(_06894_),
    .B(_07447_),
    .X(_07869_));
 sky130_fd_sc_hd__or2_1 _14698_ (.A(_07584_),
    .B(_07509_),
    .X(_07870_));
 sky130_fd_sc_hd__o22a_1 _14699_ (.A1(_06894_),
    .A2(_07413_),
    .B1(_07447_),
    .B2(_07139_),
    .X(_07871_));
 sky130_fd_sc_hd__o21bai_1 _14700_ (.A1(_07837_),
    .A2(_07869_),
    .B1_N(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__o22a_1 _14701_ (.A1(_07837_),
    .A2(_07869_),
    .B1(_07870_),
    .B2(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__or2_1 _14702_ (.A(_07868_),
    .B(_07873_),
    .X(_07874_));
 sky130_fd_sc_hd__xnor2_1 _14703_ (.A(_07862_),
    .B(_07863_),
    .Y(_07875_));
 sky130_fd_sc_hd__nand2_1 _14704_ (.A(_07868_),
    .B(_07873_),
    .Y(_07876_));
 sky130_fd_sc_hd__and2_1 _14705_ (.A(_07874_),
    .B(_07876_),
    .X(_07877_));
 sky130_fd_sc_hd__nand2_1 _14706_ (.A(_07875_),
    .B(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__and2b_1 _14707_ (.A_N(_07842_),
    .B(_07841_),
    .X(_07879_));
 sky130_fd_sc_hd__xnor2_1 _14708_ (.A(_07832_),
    .B(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__a21o_1 _14709_ (.A1(_07874_),
    .A2(_07878_),
    .B1(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__inv_2 _14710_ (.A(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__and2_1 _14711_ (.A(_07860_),
    .B(_07865_),
    .X(_07883_));
 sky130_fd_sc_hd__nor2_1 _14712_ (.A(_07866_),
    .B(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__nand3_1 _14713_ (.A(_07880_),
    .B(_07874_),
    .C(_07878_),
    .Y(_07885_));
 sky130_fd_sc_hd__and3_1 _14714_ (.A(_07881_),
    .B(_07884_),
    .C(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__a211o_1 _14715_ (.A1(_07848_),
    .A2(_07867_),
    .B1(_07882_),
    .C1(_07886_),
    .X(_07887_));
 sky130_fd_sc_hd__o211ai_1 _14716_ (.A1(_07882_),
    .A2(_07886_),
    .B1(_07848_),
    .C1(_07867_),
    .Y(_07888_));
 sky130_fd_sc_hd__a21bo_1 _14717_ (.A1(_07866_),
    .A2(_07887_),
    .B1_N(_07888_),
    .X(_07889_));
 sky130_fd_sc_hd__xor2_1 _14718_ (.A(_07853_),
    .B(_07852_),
    .X(_07890_));
 sky130_fd_sc_hd__and4_1 _14719_ (.A(_07854_),
    .B(_07859_),
    .C(_07889_),
    .D(_07890_),
    .X(_07891_));
 sky130_fd_sc_hd__xor2_1 _14720_ (.A(_07857_),
    .B(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__nor2_1 _14721_ (.A(_07859_),
    .B(_07889_),
    .Y(_07893_));
 sky130_fd_sc_hd__and3_1 _14722_ (.A(_07866_),
    .B(_07888_),
    .C(_07887_),
    .X(_07894_));
 sky130_fd_sc_hd__a21oi_1 _14723_ (.A1(_07888_),
    .A2(_07887_),
    .B1(_07866_),
    .Y(_07895_));
 sky130_fd_sc_hd__or2_1 _14724_ (.A(_07875_),
    .B(_07877_),
    .X(_07896_));
 sky130_fd_sc_hd__nand2_1 _14725_ (.A(_07878_),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__or2_1 _14726_ (.A(_07139_),
    .B(_07509_),
    .X(_07898_));
 sky130_fd_sc_hd__or2_1 _14727_ (.A(_07869_),
    .B(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__xnor2_1 _14728_ (.A(_07869_),
    .B(_07898_),
    .Y(_07900_));
 sky130_fd_sc_hd__or3_1 _14729_ (.A(_07584_),
    .B(_07733_),
    .C(_07900_),
    .X(_07901_));
 sky130_fd_sc_hd__xnor2_1 _14730_ (.A(_07870_),
    .B(_07872_),
    .Y(_07902_));
 sky130_fd_sc_hd__a21o_1 _14731_ (.A1(_07899_),
    .A2(_07901_),
    .B1(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__or2_1 _14732_ (.A(_07236_),
    .B(_07611_),
    .X(_07904_));
 sky130_fd_sc_hd__nor3_1 _14733_ (.A(_07455_),
    .B(_07733_),
    .C(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__o22a_1 _14734_ (.A1(_07455_),
    .A2(_07611_),
    .B1(_07733_),
    .B2(_07236_),
    .X(_07906_));
 sky130_fd_sc_hd__nor2_1 _14735_ (.A(_07905_),
    .B(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__nand3_1 _14736_ (.A(_07902_),
    .B(_07899_),
    .C(_07901_),
    .Y(_07908_));
 sky130_fd_sc_hd__and2_1 _14737_ (.A(_07903_),
    .B(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__nand2_1 _14738_ (.A(_07907_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__or2_1 _14739_ (.A(_07907_),
    .B(_07909_),
    .X(_07911_));
 sky130_fd_sc_hd__and2_1 _14740_ (.A(_07910_),
    .B(_07911_),
    .X(_07912_));
 sky130_fd_sc_hd__or2_1 _14741_ (.A(_06894_),
    .B(_07509_),
    .X(_07913_));
 sky130_fd_sc_hd__nor2_1 _14742_ (.A(_07584_),
    .B(_07611_),
    .Y(_07914_));
 sky130_fd_sc_hd__nor2_1 _14743_ (.A(_07139_),
    .B(_07561_),
    .Y(_07915_));
 sky130_fd_sc_hd__xnor2_1 _14744_ (.A(_07913_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__and2_1 _14745_ (.A(_07914_),
    .B(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__inv_2 _14746_ (.A(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__o31a_1 _14747_ (.A1(_07139_),
    .A2(_07733_),
    .A3(_07913_),
    .B1(_07918_),
    .X(_07919_));
 sky130_fd_sc_hd__nor2_1 _14748_ (.A(_07584_),
    .B(_07733_),
    .Y(_07920_));
 sky130_fd_sc_hd__xnor2_1 _14749_ (.A(_07920_),
    .B(_07900_),
    .Y(_07921_));
 sky130_fd_sc_hd__nor2_1 _14750_ (.A(_06869_),
    .B(_07917_),
    .Y(_07922_));
 sky130_fd_sc_hd__o211a_1 _14751_ (.A1(_07914_),
    .A2(_07916_),
    .B1(_07922_),
    .C1(_07277_),
    .X(_07923_));
 sky130_fd_sc_hd__and4bb_1 _14752_ (.A_N(_07904_),
    .B_N(_07919_),
    .C(_07921_),
    .D(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__o21bai_1 _14753_ (.A1(_07904_),
    .A2(_07919_),
    .B1_N(_07923_),
    .Y(_07925_));
 sky130_fd_sc_hd__nand2_1 _14754_ (.A(_07904_),
    .B(_07919_),
    .Y(_07926_));
 sky130_fd_sc_hd__a21o_1 _14755_ (.A1(_07921_),
    .A2(_07923_),
    .B1(_07926_),
    .X(_07927_));
 sky130_fd_sc_hd__o221a_1 _14756_ (.A1(_07912_),
    .A2(_07924_),
    .B1(_07925_),
    .B2(_07921_),
    .C1(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__nor2_1 _14757_ (.A(_07905_),
    .B(_07928_),
    .Y(_07929_));
 sky130_fd_sc_hd__a31o_1 _14758_ (.A1(_07897_),
    .A2(_07903_),
    .A3(_07910_),
    .B1(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__a21o_1 _14759_ (.A1(_07903_),
    .A2(_07910_),
    .B1(_07897_),
    .X(_07931_));
 sky130_fd_sc_hd__nand2_1 _14760_ (.A(_07905_),
    .B(_07928_),
    .Y(_07932_));
 sky130_fd_sc_hd__a21oi_1 _14761_ (.A1(_07881_),
    .A2(_07885_),
    .B1(_07884_),
    .Y(_07933_));
 sky130_fd_sc_hd__a311o_1 _14762_ (.A1(_07930_),
    .A2(_07931_),
    .A3(_07932_),
    .B1(_07933_),
    .C1(_07886_),
    .X(_07934_));
 sky130_fd_sc_hd__or3_1 _14763_ (.A(_07894_),
    .B(_07895_),
    .C(_07934_),
    .X(_07935_));
 sky130_fd_sc_hd__and4bb_1 _14764_ (.A_N(_07893_),
    .B_N(_07935_),
    .C(_07854_),
    .D(_07890_),
    .X(_07936_));
 sky130_fd_sc_hd__and2_1 _14765_ (.A(_07857_),
    .B(_07891_),
    .X(_07937_));
 sky130_fd_sc_hd__a21o_1 _14766_ (.A1(_07892_),
    .A2(_07936_),
    .B1(_07937_),
    .X(_07938_));
 sky130_fd_sc_hd__nor2_1 _14767_ (.A(_07816_),
    .B(_07856_),
    .Y(_07939_));
 sky130_fd_sc_hd__xnor2_1 _14768_ (.A(_07817_),
    .B(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__a22o_1 _14769_ (.A1(_07856_),
    .A2(_07817_),
    .B1(_07938_),
    .B2(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__nor2_1 _14770_ (.A(_07770_),
    .B(_07818_),
    .Y(_07942_));
 sky130_fd_sc_hd__xnor2_1 _14771_ (.A(_07771_),
    .B(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__a22o_1 _14772_ (.A1(_07771_),
    .A2(_07818_),
    .B1(_07941_),
    .B2(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__nor3_1 _14773_ (.A(_07718_),
    .B(_07720_),
    .C(_07772_),
    .Y(_07945_));
 sky130_fd_sc_hd__a211oi_1 _14774_ (.A1(_07720_),
    .A2(_07772_),
    .B1(_07945_),
    .C1(_07721_),
    .Y(_07946_));
 sky130_fd_sc_hd__a22o_1 _14775_ (.A1(_07720_),
    .A2(_07772_),
    .B1(_07944_),
    .B2(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__nor2_1 _14776_ (.A(_07665_),
    .B(_07721_),
    .Y(_07948_));
 sky130_fd_sc_hd__xnor2_1 _14777_ (.A(_07666_),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__a22oi_2 _14778_ (.A1(_07666_),
    .A2(_07721_),
    .B1(_07947_),
    .B2(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__o21a_1 _14779_ (.A1(_07606_),
    .A2(_07668_),
    .B1(_07555_),
    .X(_07951_));
 sky130_fd_sc_hd__inv_2 _14780_ (.A(_07951_),
    .Y(_07952_));
 sky130_fd_sc_hd__o31a_2 _14781_ (.A1(_07608_),
    .A2(_07671_),
    .A3(_07950_),
    .B1(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__o21ba_1 _14782_ (.A1(_07553_),
    .A2(_07953_),
    .B1_N(_07550_),
    .X(_07954_));
 sky130_fd_sc_hd__xnor2_2 _14783_ (.A(_07505_),
    .B(_07954_),
    .Y(_07955_));
 sky130_fd_sc_hd__xnor2_1 _14784_ (.A(_07553_),
    .B(_07953_),
    .Y(_07956_));
 sky130_fd_sc_hd__nor2_1 _14785_ (.A(_06646_),
    .B(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__buf_2 _14786_ (.A(_06726_),
    .X(_07958_));
 sky130_fd_sc_hd__a211o_1 _14787_ (.A1(_06646_),
    .A2(_07955_),
    .B1(_07957_),
    .C1(_07958_),
    .X(_07959_));
 sky130_fd_sc_hd__buf_2 _14788_ (.A(_06829_),
    .X(_07960_));
 sky130_fd_sc_hd__inv_2 _14789_ (.A(_07505_),
    .Y(_07961_));
 sky130_fd_sc_hd__o21ai_1 _14790_ (.A1(_07500_),
    .A2(_07550_),
    .B1(_07504_),
    .Y(_07962_));
 sky130_fd_sc_hd__o31ai_4 _14791_ (.A1(_07553_),
    .A2(_07953_),
    .A3(_07961_),
    .B1(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__a2111o_1 _14792_ (.A1(_07062_),
    .A2(_07433_),
    .B1(_07439_),
    .C1(_07430_),
    .D1(_07437_),
    .X(_07964_));
 sky130_fd_sc_hd__nor2_2 _14793_ (.A(_07503_),
    .B(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__xnor2_2 _14794_ (.A(_07963_),
    .B(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__inv_2 _14795_ (.A(_07965_),
    .Y(_07967_));
 sky130_fd_sc_hd__and3_1 _14796_ (.A(_06646_),
    .B(_07963_),
    .C(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__a211o_1 _14797_ (.A1(_07960_),
    .A2(_07966_),
    .B1(_07968_),
    .C1(_06724_),
    .X(_07969_));
 sky130_fd_sc_hd__buf_2 _14798_ (.A(_06705_),
    .X(_07970_));
 sky130_fd_sc_hd__a21o_1 _14799_ (.A1(_07959_),
    .A2(_07969_),
    .B1(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__and2_1 _14800_ (.A(_06672_),
    .B(_06707_),
    .X(_07972_));
 sky130_fd_sc_hd__a21oi_1 _14801_ (.A1(_06849_),
    .A2(_07970_),
    .B1(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__xnor2_1 _14802_ (.A(_07947_),
    .B(_07949_),
    .Y(_07974_));
 sky130_fd_sc_hd__xnor2_1 _14803_ (.A(_07944_),
    .B(_07946_),
    .Y(_07975_));
 sky130_fd_sc_hd__or2_1 _14804_ (.A(_06645_),
    .B(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__o21ai_1 _14805_ (.A1(_06829_),
    .A2(_07974_),
    .B1(_07976_),
    .Y(_07977_));
 sky130_fd_sc_hd__o21ba_1 _14806_ (.A1(_07671_),
    .A2(_07950_),
    .B1_N(_07668_),
    .X(_07978_));
 sky130_fd_sc_hd__xnor2_1 _14807_ (.A(_07607_),
    .B(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__xnor2_1 _14808_ (.A(_07670_),
    .B(_07950_),
    .Y(_07980_));
 sky130_fd_sc_hd__mux2_1 _14809_ (.A0(_07979_),
    .A1(_07980_),
    .S(_06829_),
    .X(_07981_));
 sky130_fd_sc_hd__mux2_1 _14810_ (.A0(_07977_),
    .A1(_07981_),
    .S(_07958_),
    .X(_07982_));
 sky130_fd_sc_hd__xnor2_1 _14811_ (.A(_07892_),
    .B(_07936_),
    .Y(_07983_));
 sky130_fd_sc_hd__or2_1 _14812_ (.A(_07960_),
    .B(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__xnor2_1 _14813_ (.A(_07941_),
    .B(_07943_),
    .Y(_07985_));
 sky130_fd_sc_hd__or2_1 _14814_ (.A(_06829_),
    .B(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__xor2_1 _14815_ (.A(_07938_),
    .B(_07940_),
    .X(_07987_));
 sky130_fd_sc_hd__nand2_1 _14816_ (.A(_06829_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__and2_1 _14817_ (.A(_07986_),
    .B(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__mux2_1 _14818_ (.A0(_07984_),
    .A1(_07989_),
    .S(_07958_),
    .X(_07990_));
 sky130_fd_sc_hd__nor2_1 _14819_ (.A(_07970_),
    .B(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__a21o_1 _14820_ (.A1(_07970_),
    .A2(_07982_),
    .B1(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__a22o_1 _14821_ (.A1(_07971_),
    .A2(_07973_),
    .B1(_07992_),
    .B2(_07972_),
    .X(_07993_));
 sky130_fd_sc_hd__or2_1 _14822_ (.A(_07437_),
    .B(_06640_),
    .X(_07994_));
 sky130_fd_sc_hd__clkbuf_4 _14823_ (.A(_07994_),
    .X(_07995_));
 sky130_fd_sc_hd__buf_2 _14824_ (.A(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__a21o_2 _14825_ (.A1(_06587_),
    .A2(_07993_),
    .B1(_07996_),
    .X(_07997_));
 sky130_fd_sc_hd__and4b_2 _14826_ (.A_N(_04570_),
    .B(_04571_),
    .C(_04568_),
    .D(_06096_),
    .X(_07998_));
 sky130_fd_sc_hd__buf_4 _14827_ (.A(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__mux2_1 _14828_ (.A0(\rbzero.wall_tracer.stepDistY[-11] ),
    .A1(_07997_),
    .S(_07999_),
    .X(_08000_));
 sky130_fd_sc_hd__clkbuf_1 _14829_ (.A(_08000_),
    .X(_00391_));
 sky130_fd_sc_hd__and3_1 _14830_ (.A(_06829_),
    .B(_07963_),
    .C(_07967_),
    .X(_08001_));
 sky130_fd_sc_hd__mux2_1 _14831_ (.A0(_07966_),
    .A1(_07955_),
    .S(_07960_),
    .X(_08002_));
 sky130_fd_sc_hd__mux2_1 _14832_ (.A0(_08001_),
    .A1(_08002_),
    .S(_06724_),
    .X(_08003_));
 sky130_fd_sc_hd__a21o_1 _14833_ (.A1(_06780_),
    .A2(_08003_),
    .B1(_07972_),
    .X(_08004_));
 sky130_fd_sc_hd__and2_1 _14834_ (.A(_06645_),
    .B(_07987_),
    .X(_08005_));
 sky130_fd_sc_hd__o21bai_1 _14835_ (.A1(_06646_),
    .A2(_07983_),
    .B1_N(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__nor2_1 _14836_ (.A(_06829_),
    .B(_07975_),
    .Y(_08007_));
 sky130_fd_sc_hd__nor2_1 _14837_ (.A(_06646_),
    .B(_07985_),
    .Y(_08008_));
 sky130_fd_sc_hd__or2_1 _14838_ (.A(_08007_),
    .B(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__nor2_1 _14839_ (.A(_06645_),
    .B(_07974_),
    .Y(_08010_));
 sky130_fd_sc_hd__and2_1 _14840_ (.A(_06645_),
    .B(_07980_),
    .X(_08011_));
 sky130_fd_sc_hd__or2_1 _14841_ (.A(_08010_),
    .B(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__xnor2_1 _14842_ (.A(_07552_),
    .B(_07953_),
    .Y(_08013_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(_08013_),
    .A1(_07979_),
    .S(_06829_),
    .X(_08014_));
 sky130_fd_sc_hd__mux4_2 _14844_ (.A0(_08006_),
    .A1(_08009_),
    .A2(_08012_),
    .A3(_08014_),
    .S0(_07958_),
    .S1(_06705_),
    .X(_08015_));
 sky130_fd_sc_hd__or2_1 _14845_ (.A(_06719_),
    .B(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__a31o_2 _14846_ (.A1(_06587_),
    .A2(_08004_),
    .A3(_08016_),
    .B1(_07996_),
    .X(_08017_));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(\rbzero.wall_tracer.stepDistY[-10] ),
    .A1(_08017_),
    .S(_07999_),
    .X(_08018_));
 sky130_fd_sc_hd__clkbuf_1 _14848_ (.A(_08018_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _14849_ (.A0(_07966_),
    .A1(_07955_),
    .S(_06646_),
    .X(_08019_));
 sky130_fd_sc_hd__or3_1 _14850_ (.A(_07437_),
    .B(_06835_),
    .C(_07968_),
    .X(_08020_));
 sky130_fd_sc_hd__o211a_1 _14851_ (.A1(_06731_),
    .A2(_08019_),
    .B1(_08020_),
    .C1(_06730_),
    .X(_08021_));
 sky130_fd_sc_hd__mux2_1 _14852_ (.A0(_08013_),
    .A1(_07979_),
    .S(_06646_),
    .X(_08022_));
 sky130_fd_sc_hd__nor2_1 _14853_ (.A(_07960_),
    .B(_07974_),
    .Y(_08023_));
 sky130_fd_sc_hd__a21o_1 _14854_ (.A1(_07960_),
    .A2(_07980_),
    .B1(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__and2_1 _14855_ (.A(_06835_),
    .B(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__buf_2 _14856_ (.A(_06730_),
    .X(_08026_));
 sky130_fd_sc_hd__a211o_1 _14857_ (.A1(_06731_),
    .A2(_08022_),
    .B1(_08025_),
    .C1(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__nand2_1 _14858_ (.A(_07986_),
    .B(_07976_),
    .Y(_08028_));
 sky130_fd_sc_hd__or2_1 _14859_ (.A(_06685_),
    .B(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__nand2_1 _14860_ (.A(_06587_),
    .B(_06729_),
    .Y(_08030_));
 sky130_fd_sc_hd__a31oi_1 _14861_ (.A1(_06690_),
    .A2(_07988_),
    .A3(_07984_),
    .B1(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__a31o_1 _14862_ (.A1(_08027_),
    .A2(_08029_),
    .A3(_08031_),
    .B1(_07995_),
    .X(_08032_));
 sky130_fd_sc_hd__a21o_1 _14863_ (.A1(_06558_),
    .A2(_08021_),
    .B1(_08032_),
    .X(_08033_));
 sky130_fd_sc_hd__mux2_1 _14864_ (.A0(\rbzero.wall_tracer.stepDistY[-9] ),
    .A1(_08033_),
    .S(_07999_),
    .X(_08034_));
 sky130_fd_sc_hd__clkbuf_1 _14865_ (.A(_08034_),
    .X(_00393_));
 sky130_fd_sc_hd__buf_2 _14866_ (.A(_06731_),
    .X(_08035_));
 sky130_fd_sc_hd__nor2_1 _14867_ (.A(_07960_),
    .B(_07956_),
    .Y(_08036_));
 sky130_fd_sc_hd__a21oi_1 _14868_ (.A1(_07960_),
    .A2(_07955_),
    .B1(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__a21oi_1 _14869_ (.A1(_07960_),
    .A2(_07979_),
    .B1(_08011_),
    .Y(_08038_));
 sky130_fd_sc_hd__and2_1 _14870_ (.A(_06835_),
    .B(_08038_),
    .X(_08039_));
 sky130_fd_sc_hd__a211o_1 _14871_ (.A1(_08035_),
    .A2(_08037_),
    .B1(_08039_),
    .C1(_08026_),
    .X(_08040_));
 sky130_fd_sc_hd__nor2_1 _14872_ (.A(_08010_),
    .B(_08007_),
    .Y(_08041_));
 sky130_fd_sc_hd__nor2_1 _14873_ (.A(_08008_),
    .B(_08005_),
    .Y(_08042_));
 sky130_fd_sc_hd__o221a_1 _14874_ (.A1(_06685_),
    .A2(_08041_),
    .B1(_08042_),
    .B2(_06721_),
    .C1(_06729_),
    .X(_08043_));
 sky130_fd_sc_hd__a21o_1 _14875_ (.A1(_06646_),
    .A2(_07966_),
    .B1(_08001_),
    .X(_08044_));
 sky130_fd_sc_hd__a21oi_1 _14876_ (.A1(_06690_),
    .A2(_08044_),
    .B1(_06729_),
    .Y(_08045_));
 sky130_fd_sc_hd__a21oi_1 _14877_ (.A1(_08040_),
    .A2(_08043_),
    .B1(_08045_),
    .Y(_08046_));
 sky130_fd_sc_hd__nand2_1 _14878_ (.A(_07958_),
    .B(_08006_),
    .Y(_08047_));
 sky130_fd_sc_hd__nor2_1 _14879_ (.A(_06780_),
    .B(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__a21o_1 _14880_ (.A1(_06832_),
    .A2(_08048_),
    .B1(_07996_),
    .X(_08049_));
 sky130_fd_sc_hd__a21o_2 _14881_ (.A1(_06587_),
    .A2(_08046_),
    .B1(_08049_),
    .X(_08050_));
 sky130_fd_sc_hd__mux2_1 _14882_ (.A0(\rbzero.wall_tracer.stepDistY[-8] ),
    .A1(_08050_),
    .S(_07999_),
    .X(_08051_));
 sky130_fd_sc_hd__clkbuf_1 _14883_ (.A(_08051_),
    .X(_00394_));
 sky130_fd_sc_hd__or2_1 _14884_ (.A(_07437_),
    .B(_07968_),
    .X(_08052_));
 sky130_fd_sc_hd__and2_1 _14885_ (.A(_06690_),
    .B(_08052_),
    .X(_08053_));
 sky130_fd_sc_hd__mux2_1 _14886_ (.A0(_08028_),
    .A1(_08024_),
    .S(_08035_),
    .X(_08054_));
 sky130_fd_sc_hd__a21oi_1 _14887_ (.A1(_08026_),
    .A2(_08054_),
    .B1(_06696_),
    .Y(_08055_));
 sky130_fd_sc_hd__xnor2_1 _14888_ (.A(_07963_),
    .B(_07967_),
    .Y(_08056_));
 sky130_fd_sc_hd__xnor2_1 _14889_ (.A(_07961_),
    .B(_07954_),
    .Y(_08057_));
 sky130_fd_sc_hd__mux2_1 _14890_ (.A0(_08056_),
    .A1(_08057_),
    .S(_06646_),
    .X(_08058_));
 sky130_fd_sc_hd__nor2_1 _14891_ (.A(_08035_),
    .B(_08022_),
    .Y(_08059_));
 sky130_fd_sc_hd__a211o_1 _14892_ (.A1(_08035_),
    .A2(_08058_),
    .B1(_08059_),
    .C1(_08026_),
    .X(_08060_));
 sky130_fd_sc_hd__a2bb2o_1 _14893_ (.A1_N(_06729_),
    .A2_N(_08053_),
    .B1(_08055_),
    .B2(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__nor2_4 _14894_ (.A(_07437_),
    .B(_06640_),
    .Y(_08062_));
 sky130_fd_sc_hd__o31a_1 _14895_ (.A1(_06587_),
    .A2(_06780_),
    .A3(_07990_),
    .B1(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__o21ai_4 _14896_ (.A1(_06650_),
    .A2(_08061_),
    .B1(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__mux2_1 _14897_ (.A0(\rbzero.wall_tracer.stepDistY[-7] ),
    .A1(_08064_),
    .S(_07999_),
    .X(_08065_));
 sky130_fd_sc_hd__clkbuf_1 _14898_ (.A(_08065_),
    .X(_00395_));
 sky130_fd_sc_hd__a211o_1 _14899_ (.A1(_07960_),
    .A2(_07955_),
    .B1(_08036_),
    .C1(_06731_),
    .X(_08066_));
 sky130_fd_sc_hd__o21a_1 _14900_ (.A1(_06835_),
    .A2(_08044_),
    .B1(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__mux2_1 _14901_ (.A0(_08041_),
    .A1(_08038_),
    .S(_08035_),
    .X(_08068_));
 sky130_fd_sc_hd__nand2_1 _14902_ (.A(_08026_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__nor2_2 _14903_ (.A(_06650_),
    .B(_06696_),
    .Y(_08070_));
 sky130_fd_sc_hd__o211a_1 _14904_ (.A1(_08026_),
    .A2(_08067_),
    .B1(_08069_),
    .C1(_08070_),
    .X(_08071_));
 sky130_fd_sc_hd__mux2_1 _14905_ (.A0(_08006_),
    .A1(_08009_),
    .S(_07958_),
    .X(_08072_));
 sky130_fd_sc_hd__and3_1 _14906_ (.A(_07970_),
    .B(_06832_),
    .C(_08072_),
    .X(_08073_));
 sky130_fd_sc_hd__or3_2 _14907_ (.A(_07996_),
    .B(_08071_),
    .C(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__mux2_1 _14908_ (.A0(\rbzero.wall_tracer.stepDistY[-6] ),
    .A1(_08074_),
    .S(_07999_),
    .X(_08075_));
 sky130_fd_sc_hd__clkbuf_1 _14909_ (.A(_08075_),
    .X(_00396_));
 sky130_fd_sc_hd__nand2_1 _14910_ (.A(_08035_),
    .B(_07968_),
    .Y(_08076_));
 sky130_fd_sc_hd__o211a_1 _14911_ (.A1(_08035_),
    .A2(_08058_),
    .B1(_08076_),
    .C1(_06661_),
    .X(_08077_));
 sky130_fd_sc_hd__a211o_1 _14912_ (.A1(_08035_),
    .A2(_08022_),
    .B1(_08025_),
    .C1(_06661_),
    .X(_08078_));
 sky130_fd_sc_hd__nand2_1 _14913_ (.A(_08070_),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__clkinv_2 _14914_ (.A(_07989_),
    .Y(_08080_));
 sky130_fd_sc_hd__mux2_1 _14915_ (.A0(_08080_),
    .A1(_07977_),
    .S(_06726_),
    .X(_08081_));
 sky130_fd_sc_hd__nand2_1 _14916_ (.A(_06705_),
    .B(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__o31a_1 _14917_ (.A1(_06730_),
    .A2(_06724_),
    .A3(_07984_),
    .B1(_08082_),
    .X(_08083_));
 sky130_fd_sc_hd__o21ai_1 _14918_ (.A1(_06744_),
    .A2(_08083_),
    .B1(_08062_),
    .Y(_08084_));
 sky130_fd_sc_hd__o21bai_4 _14919_ (.A1(_08077_),
    .A2(_08079_),
    .B1_N(_08084_),
    .Y(_08085_));
 sky130_fd_sc_hd__mux2_1 _14920_ (.A0(\rbzero.wall_tracer.stepDistY[-5] ),
    .A1(_08085_),
    .S(_07999_),
    .X(_08086_));
 sky130_fd_sc_hd__clkbuf_1 _14921_ (.A(_08086_),
    .X(_00397_));
 sky130_fd_sc_hd__a21o_1 _14922_ (.A1(_08035_),
    .A2(_08037_),
    .B1(_08039_),
    .X(_08087_));
 sky130_fd_sc_hd__a21oi_1 _14923_ (.A1(_06835_),
    .A2(_08044_),
    .B1(_08026_),
    .Y(_08088_));
 sky130_fd_sc_hd__a211o_1 _14924_ (.A1(_08026_),
    .A2(_08087_),
    .B1(_08088_),
    .C1(_08030_),
    .X(_08089_));
 sky130_fd_sc_hd__or2_1 _14925_ (.A(_07958_),
    .B(_08009_),
    .X(_08090_));
 sky130_fd_sc_hd__o21ai_1 _14926_ (.A1(_06724_),
    .A2(_08012_),
    .B1(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__mux2_1 _14927_ (.A0(_08047_),
    .A1(_08091_),
    .S(_07970_),
    .X(_08092_));
 sky130_fd_sc_hd__or2_1 _14928_ (.A(_06744_),
    .B(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__nand3_2 _14929_ (.A(_08062_),
    .B(_08089_),
    .C(_08093_),
    .Y(_08094_));
 sky130_fd_sc_hd__mux2_1 _14930_ (.A0(\rbzero.wall_tracer.stepDistY[-4] ),
    .A1(_08094_),
    .S(_07999_),
    .X(_08095_));
 sky130_fd_sc_hd__clkbuf_1 _14931_ (.A(_08095_),
    .X(_00398_));
 sky130_fd_sc_hd__a21oi_1 _14932_ (.A1(_08035_),
    .A2(_08058_),
    .B1(_08059_),
    .Y(_08096_));
 sky130_fd_sc_hd__a21o_1 _14933_ (.A1(_06835_),
    .A2(_08052_),
    .B1(_08026_),
    .X(_08097_));
 sky130_fd_sc_hd__o211ai_4 _14934_ (.A1(_06661_),
    .A2(_08096_),
    .B1(_08097_),
    .C1(_08070_),
    .Y(_08098_));
 sky130_fd_sc_hd__nand2_1 _14935_ (.A(_06832_),
    .B(_07992_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand3_4 _14936_ (.A(_08062_),
    .B(_08098_),
    .C(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__mux2_1 _14937_ (.A0(\rbzero.wall_tracer.stepDistY[-3] ),
    .A1(_08100_),
    .S(_07999_),
    .X(_08101_));
 sky130_fd_sc_hd__clkbuf_1 _14938_ (.A(_08101_),
    .X(_00399_));
 sky130_fd_sc_hd__o211a_1 _14939_ (.A1(_06835_),
    .A2(_08044_),
    .B1(_08066_),
    .C1(_06730_),
    .X(_08102_));
 sky130_fd_sc_hd__a21o_1 _14940_ (.A1(_06832_),
    .A2(_08015_),
    .B1(_07995_),
    .X(_08103_));
 sky130_fd_sc_hd__a21o_4 _14941_ (.A1(_08070_),
    .A2(_08102_),
    .B1(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__mux2_1 _14942_ (.A0(\rbzero.wall_tracer.stepDistY[-2] ),
    .A1(_08104_),
    .S(_07999_),
    .X(_08105_));
 sky130_fd_sc_hd__clkbuf_1 _14943_ (.A(_08105_),
    .X(_00400_));
 sky130_fd_sc_hd__or2_1 _14944_ (.A(_07958_),
    .B(_07981_),
    .X(_08106_));
 sky130_fd_sc_hd__a211o_1 _14945_ (.A1(_06646_),
    .A2(_07955_),
    .B1(_07957_),
    .C1(_06724_),
    .X(_08107_));
 sky130_fd_sc_hd__and2_1 _14946_ (.A(_06780_),
    .B(_08081_),
    .X(_08108_));
 sky130_fd_sc_hd__a311o_1 _14947_ (.A1(_06705_),
    .A2(_08106_),
    .A3(_08107_),
    .B1(_08108_),
    .C1(_07972_),
    .X(_08109_));
 sky130_fd_sc_hd__a22o_1 _14948_ (.A1(_06729_),
    .A2(_08021_),
    .B1(_08109_),
    .B2(_06832_),
    .X(_08110_));
 sky130_fd_sc_hd__or2_4 _14949_ (.A(_07995_),
    .B(_08110_),
    .X(_08111_));
 sky130_fd_sc_hd__buf_4 _14950_ (.A(_07998_),
    .X(_08112_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(\rbzero.wall_tracer.stepDistY[-1] ),
    .A1(_08111_),
    .S(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__clkbuf_1 _14952_ (.A(_08113_),
    .X(_00401_));
 sky130_fd_sc_hd__mux4_2 _14953_ (.A0(_08002_),
    .A1(_08012_),
    .A2(_08014_),
    .A3(_08009_),
    .S0(_06780_),
    .S1(_06724_),
    .X(_08114_));
 sky130_fd_sc_hd__a21o_1 _14954_ (.A1(_06720_),
    .A2(_08048_),
    .B1(_07995_),
    .X(_08115_));
 sky130_fd_sc_hd__a31o_1 _14955_ (.A1(_06729_),
    .A2(_06690_),
    .A3(_08044_),
    .B1(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__a21o_4 _14956_ (.A1(_06832_),
    .A2(_08114_),
    .B1(_08116_),
    .X(_08117_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(\rbzero.wall_tracer.stepDistY[0] ),
    .A1(_08117_),
    .S(_08112_),
    .X(_08118_));
 sky130_fd_sc_hd__clkbuf_1 _14958_ (.A(_08118_),
    .X(_00402_));
 sky130_fd_sc_hd__and2_1 _14959_ (.A(_07959_),
    .B(_07969_),
    .X(_08119_));
 sky130_fd_sc_hd__mux2_1 _14960_ (.A0(_08119_),
    .A1(_07982_),
    .S(_06780_),
    .X(_08120_));
 sky130_fd_sc_hd__a221o_4 _14961_ (.A1(_06729_),
    .A2(_08053_),
    .B1(_08120_),
    .B2(_06832_),
    .C1(_07995_),
    .X(_08121_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(\rbzero.wall_tracer.stepDistY[1] ),
    .A1(_08121_),
    .S(_08112_),
    .X(_08122_));
 sky130_fd_sc_hd__clkbuf_1 _14963_ (.A(_08122_),
    .X(_00403_));
 sky130_fd_sc_hd__and2_1 _14964_ (.A(_07970_),
    .B(_08072_),
    .X(_08123_));
 sky130_fd_sc_hd__mux2_1 _14965_ (.A0(_08012_),
    .A1(_08014_),
    .S(_07958_),
    .X(_08124_));
 sky130_fd_sc_hd__mux2_1 _14966_ (.A0(_08003_),
    .A1(_08124_),
    .S(_06780_),
    .X(_08125_));
 sky130_fd_sc_hd__a221o_4 _14967_ (.A1(_06720_),
    .A2(_08123_),
    .B1(_08125_),
    .B2(_06832_),
    .C1(_07995_),
    .X(_08126_));
 sky130_fd_sc_hd__mux2_1 _14968_ (.A0(\rbzero.wall_tracer.stepDistY[2] ),
    .A1(_08126_),
    .S(_08112_),
    .X(_08127_));
 sky130_fd_sc_hd__clkbuf_1 _14969_ (.A(_08127_),
    .X(_00404_));
 sky130_fd_sc_hd__a21o_1 _14970_ (.A1(_07960_),
    .A2(_07966_),
    .B1(_07968_),
    .X(_08128_));
 sky130_fd_sc_hd__a21o_1 _14971_ (.A1(_06724_),
    .A2(_08128_),
    .B1(_06780_),
    .X(_08129_));
 sky130_fd_sc_hd__and2_1 _14972_ (.A(_08106_),
    .B(_08107_),
    .X(_08130_));
 sky130_fd_sc_hd__or2_1 _14973_ (.A(_07970_),
    .B(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__nand2_1 _14974_ (.A(_06610_),
    .B(_06612_),
    .Y(_08132_));
 sky130_fd_sc_hd__o21ai_1 _14975_ (.A1(_08132_),
    .A2(_08083_),
    .B1(_08062_),
    .Y(_08133_));
 sky130_fd_sc_hd__a31o_2 _14976_ (.A1(_06832_),
    .A2(_08129_),
    .A3(_08131_),
    .B1(_08133_),
    .X(_08134_));
 sky130_fd_sc_hd__mux2_1 _14977_ (.A0(\rbzero.wall_tracer.stepDistY[3] ),
    .A1(_08134_),
    .S(_08112_),
    .X(_08135_));
 sky130_fd_sc_hd__clkbuf_1 _14978_ (.A(_08135_),
    .X(_00405_));
 sky130_fd_sc_hd__or2_1 _14979_ (.A(_07958_),
    .B(_08014_),
    .X(_08136_));
 sky130_fd_sc_hd__o211a_1 _14980_ (.A1(_06724_),
    .A2(_08002_),
    .B1(_08136_),
    .C1(_06780_),
    .X(_08137_));
 sky130_fd_sc_hd__a311o_1 _14981_ (.A1(_06835_),
    .A2(_07970_),
    .A3(_08001_),
    .B1(_08137_),
    .C1(_07972_),
    .X(_08138_));
 sky130_fd_sc_hd__nand2_1 _14982_ (.A(_07972_),
    .B(_08092_),
    .Y(_08139_));
 sky130_fd_sc_hd__a31o_2 _14983_ (.A1(_06650_),
    .A2(_08138_),
    .A3(_08139_),
    .B1(_07996_),
    .X(_08140_));
 sky130_fd_sc_hd__mux2_1 _14984_ (.A0(\rbzero.wall_tracer.stepDistY[4] ),
    .A1(_08140_),
    .S(_08112_),
    .X(_08141_));
 sky130_fd_sc_hd__clkbuf_1 _14985_ (.A(_08141_),
    .X(_00406_));
 sky130_fd_sc_hd__a221o_2 _14986_ (.A1(_06718_),
    .A2(_08119_),
    .B1(_07992_),
    .B2(_06720_),
    .C1(_07995_),
    .X(_08142_));
 sky130_fd_sc_hd__mux2_1 _14987_ (.A0(\rbzero.wall_tracer.stepDistY[5] ),
    .A1(_08142_),
    .S(_08112_),
    .X(_08143_));
 sky130_fd_sc_hd__clkbuf_1 _14988_ (.A(_08143_),
    .X(_00407_));
 sky130_fd_sc_hd__a21o_1 _14989_ (.A1(_06720_),
    .A2(_08015_),
    .B1(_07995_),
    .X(_08144_));
 sky130_fd_sc_hd__a21o_1 _14990_ (.A1(_06718_),
    .A2(_08003_),
    .B1(_08144_),
    .X(_08145_));
 sky130_fd_sc_hd__mux2_1 _14991_ (.A0(\rbzero.wall_tracer.stepDistY[6] ),
    .A1(_08145_),
    .S(_08112_),
    .X(_08146_));
 sky130_fd_sc_hd__clkbuf_1 _14992_ (.A(_08146_),
    .X(_00408_));
 sky130_fd_sc_hd__a211o_1 _14993_ (.A1(_07970_),
    .A2(_08130_),
    .B1(_08108_),
    .C1(_06719_),
    .X(_08147_));
 sky130_fd_sc_hd__a31o_1 _14994_ (.A1(_06724_),
    .A2(_06718_),
    .A3(_08128_),
    .B1(_06720_),
    .X(_08148_));
 sky130_fd_sc_hd__a21o_1 _14995_ (.A1(_08147_),
    .A2(_08148_),
    .B1(_07996_),
    .X(_08149_));
 sky130_fd_sc_hd__mux2_1 _14996_ (.A0(\rbzero.wall_tracer.stepDistY[7] ),
    .A1(_08149_),
    .S(_08112_),
    .X(_08150_));
 sky130_fd_sc_hd__clkbuf_1 _14997_ (.A(_08150_),
    .X(_00409_));
 sky130_fd_sc_hd__a41o_1 _14998_ (.A1(_06650_),
    .A2(_08026_),
    .A3(_06835_),
    .A4(_08001_),
    .B1(_06720_),
    .X(_08151_));
 sky130_fd_sc_hd__o21a_1 _14999_ (.A1(_06719_),
    .A2(_08114_),
    .B1(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__or2_1 _15000_ (.A(_07996_),
    .B(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__mux2_1 _15001_ (.A0(\rbzero.wall_tracer.stepDistY[8] ),
    .A1(_08153_),
    .S(_08112_),
    .X(_08154_));
 sky130_fd_sc_hd__clkbuf_1 _15002_ (.A(_08154_),
    .X(_00410_));
 sky130_fd_sc_hd__a21o_1 _15003_ (.A1(_06720_),
    .A2(_08120_),
    .B1(_07996_),
    .X(_08155_));
 sky130_fd_sc_hd__mux2_1 _15004_ (.A0(\rbzero.wall_tracer.stepDistY[9] ),
    .A1(_08155_),
    .S(_07998_),
    .X(_08156_));
 sky130_fd_sc_hd__clkbuf_1 _15005_ (.A(_08156_),
    .X(_00411_));
 sky130_fd_sc_hd__and3_1 _15006_ (.A(_08062_),
    .B(_06720_),
    .C(_08125_),
    .X(_08157_));
 sky130_fd_sc_hd__mux2_1 _15007_ (.A0(\rbzero.wall_tracer.stepDistY[10] ),
    .A1(_08157_),
    .S(_07998_),
    .X(_08158_));
 sky130_fd_sc_hd__clkbuf_1 _15008_ (.A(_08158_),
    .X(_00412_));
 sky130_fd_sc_hd__nand2_1 _15009_ (.A(_06094_),
    .B(_06281_),
    .Y(_08159_));
 sky130_fd_sc_hd__clkbuf_4 _15010_ (.A(_08159_),
    .X(_08160_));
 sky130_fd_sc_hd__buf_2 _15011_ (.A(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__buf_4 _15012_ (.A(_06178_),
    .X(_08162_));
 sky130_fd_sc_hd__mux2_1 _15013_ (.A0(\rbzero.wall_tracer.trackDistY[-11] ),
    .A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .S(_08162_),
    .X(_08163_));
 sky130_fd_sc_hd__buf_4 _15014_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_08164_));
 sky130_fd_sc_hd__and2_2 _15015_ (.A(_06094_),
    .B(_06281_),
    .X(_08165_));
 sky130_fd_sc_hd__buf_2 _15016_ (.A(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__or2_1 _15017_ (.A(_08164_),
    .B(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__clkbuf_4 _15018_ (.A(_04576_),
    .X(_01633_));
 sky130_fd_sc_hd__o211a_1 _15019_ (.A1(_08161_),
    .A2(_08163_),
    .B1(_08167_),
    .C1(_01633_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _15020_ (.A0(\rbzero.wall_tracer.trackDistY[-10] ),
    .A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .S(_08162_),
    .X(_08168_));
 sky130_fd_sc_hd__inv_2 _15021_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .Y(_08169_));
 sky130_fd_sc_hd__nand2_1 _15022_ (.A(_08169_),
    .B(_08160_),
    .Y(_08170_));
 sky130_fd_sc_hd__o211a_1 _15023_ (.A1(_08161_),
    .A2(_08168_),
    .B1(_08170_),
    .C1(_01633_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _15024_ (.A0(\rbzero.wall_tracer.trackDistY[-9] ),
    .A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .S(_08162_),
    .X(_08171_));
 sky130_fd_sc_hd__or2_1 _15025_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(_08166_),
    .X(_08172_));
 sky130_fd_sc_hd__o211a_1 _15026_ (.A1(_08161_),
    .A2(_08171_),
    .B1(_08172_),
    .C1(_01633_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _15027_ (.A0(\rbzero.wall_tracer.trackDistY[-8] ),
    .A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .S(_08162_),
    .X(_08173_));
 sky130_fd_sc_hd__or2_1 _15028_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_08166_),
    .X(_08174_));
 sky130_fd_sc_hd__o211a_1 _15029_ (.A1(_08161_),
    .A2(_08173_),
    .B1(_08174_),
    .C1(_01633_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _15030_ (.A0(\rbzero.wall_tracer.trackDistY[-7] ),
    .A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .S(_08162_),
    .X(_08175_));
 sky130_fd_sc_hd__or2_1 _15031_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(_08166_),
    .X(_08176_));
 sky130_fd_sc_hd__o211a_1 _15032_ (.A1(_08161_),
    .A2(_08175_),
    .B1(_08176_),
    .C1(_01633_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _15033_ (.A0(\rbzero.wall_tracer.trackDistY[-6] ),
    .A1(\rbzero.wall_tracer.trackDistX[-6] ),
    .S(_08162_),
    .X(_08177_));
 sky130_fd_sc_hd__or2_1 _15034_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(_08166_),
    .X(_08178_));
 sky130_fd_sc_hd__o211a_1 _15035_ (.A1(_08161_),
    .A2(_08177_),
    .B1(_08178_),
    .C1(_01633_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _15036_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .S(_08162_),
    .X(_08179_));
 sky130_fd_sc_hd__or2_1 _15037_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_08166_),
    .X(_08180_));
 sky130_fd_sc_hd__o211a_1 _15038_ (.A1(_08161_),
    .A2(_08179_),
    .B1(_08180_),
    .C1(_01633_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _15039_ (.A0(\rbzero.wall_tracer.trackDistY[-4] ),
    .A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .S(_08162_),
    .X(_08181_));
 sky130_fd_sc_hd__inv_2 _15040_ (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .Y(_08182_));
 sky130_fd_sc_hd__nand2_1 _15041_ (.A(_08182_),
    .B(_08160_),
    .Y(_08183_));
 sky130_fd_sc_hd__o211a_1 _15042_ (.A1(_08161_),
    .A2(_08181_),
    .B1(_08183_),
    .C1(_01633_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _15043_ (.A0(\rbzero.wall_tracer.trackDistY[-3] ),
    .A1(\rbzero.wall_tracer.trackDistX[-3] ),
    .S(_08162_),
    .X(_08184_));
 sky130_fd_sc_hd__or2_1 _15044_ (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .B(_08166_),
    .X(_08185_));
 sky130_fd_sc_hd__buf_2 _15045_ (.A(_04576_),
    .X(_08186_));
 sky130_fd_sc_hd__o211a_1 _15046_ (.A1(_08161_),
    .A2(_08184_),
    .B1(_08185_),
    .C1(_08186_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _15047_ (.A0(\rbzero.wall_tracer.trackDistY[-2] ),
    .A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .S(_08162_),
    .X(_08187_));
 sky130_fd_sc_hd__or2_1 _15048_ (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .B(_08166_),
    .X(_08188_));
 sky130_fd_sc_hd__o211a_1 _15049_ (.A1(_08161_),
    .A2(_08187_),
    .B1(_08188_),
    .C1(_08186_),
    .X(_00422_));
 sky130_fd_sc_hd__buf_2 _15050_ (.A(_08159_),
    .X(_08189_));
 sky130_fd_sc_hd__clkbuf_4 _15051_ (.A(_06178_),
    .X(_08190_));
 sky130_fd_sc_hd__mux2_1 _15052_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .S(_08190_),
    .X(_08191_));
 sky130_fd_sc_hd__or2_1 _15053_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(_08166_),
    .X(_08192_));
 sky130_fd_sc_hd__o211a_1 _15054_ (.A1(_08189_),
    .A2(_08191_),
    .B1(_08192_),
    .C1(_08186_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _15055_ (.A0(\rbzero.wall_tracer.trackDistY[0] ),
    .A1(\rbzero.wall_tracer.trackDistX[0] ),
    .S(_08190_),
    .X(_08193_));
 sky130_fd_sc_hd__inv_2 _15056_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .Y(_08194_));
 sky130_fd_sc_hd__nand2_1 _15057_ (.A(_08194_),
    .B(_08160_),
    .Y(_08195_));
 sky130_fd_sc_hd__o211a_1 _15058_ (.A1(_08189_),
    .A2(_08193_),
    .B1(_08195_),
    .C1(_08186_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _15059_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(\rbzero.wall_tracer.trackDistX[1] ),
    .S(_08190_),
    .X(_08196_));
 sky130_fd_sc_hd__nand2_1 _15060_ (.A(_06461_),
    .B(_08160_),
    .Y(_08197_));
 sky130_fd_sc_hd__o211a_1 _15061_ (.A1(_08189_),
    .A2(_08196_),
    .B1(_08197_),
    .C1(_08186_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _15062_ (.A0(\rbzero.wall_tracer.trackDistY[2] ),
    .A1(\rbzero.wall_tracer.trackDistX[2] ),
    .S(_08190_),
    .X(_08198_));
 sky130_fd_sc_hd__or2_1 _15063_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08166_),
    .X(_08199_));
 sky130_fd_sc_hd__o211a_1 _15064_ (.A1(_08189_),
    .A2(_08198_),
    .B1(_08199_),
    .C1(_08186_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _15065_ (.A0(\rbzero.wall_tracer.trackDistY[3] ),
    .A1(\rbzero.wall_tracer.trackDistX[3] ),
    .S(_08190_),
    .X(_08200_));
 sky130_fd_sc_hd__clkinv_2 _15066_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .Y(_08201_));
 sky130_fd_sc_hd__nand2_1 _15067_ (.A(_08201_),
    .B(_08160_),
    .Y(_08202_));
 sky130_fd_sc_hd__o211a_1 _15068_ (.A1(_08189_),
    .A2(_08200_),
    .B1(_08202_),
    .C1(_08186_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _15069_ (.A0(\rbzero.wall_tracer.trackDistY[4] ),
    .A1(\rbzero.wall_tracer.trackDistX[4] ),
    .S(_08190_),
    .X(_08203_));
 sky130_fd_sc_hd__or2_1 _15070_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08165_),
    .X(_08204_));
 sky130_fd_sc_hd__o211a_1 _15071_ (.A1(_08189_),
    .A2(_08203_),
    .B1(_08204_),
    .C1(_08186_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _15072_ (.A0(\rbzero.wall_tracer.trackDistY[5] ),
    .A1(\rbzero.wall_tracer.trackDistX[5] ),
    .S(_08190_),
    .X(_08205_));
 sky130_fd_sc_hd__or2_1 _15073_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08165_),
    .X(_08206_));
 sky130_fd_sc_hd__o211a_1 _15074_ (.A1(_08189_),
    .A2(_08205_),
    .B1(_08206_),
    .C1(_08186_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _15075_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(\rbzero.wall_tracer.trackDistX[6] ),
    .S(_08190_),
    .X(_08207_));
 sky130_fd_sc_hd__or2_1 _15076_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08165_),
    .X(_08208_));
 sky130_fd_sc_hd__o211a_1 _15077_ (.A1(_08189_),
    .A2(_08207_),
    .B1(_08208_),
    .C1(_08186_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _15078_ (.A0(\rbzero.wall_tracer.trackDistY[7] ),
    .A1(\rbzero.wall_tracer.trackDistX[7] ),
    .S(_08190_),
    .X(_08209_));
 sky130_fd_sc_hd__or2_1 _15079_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08165_),
    .X(_08210_));
 sky130_fd_sc_hd__buf_4 _15080_ (.A(_04576_),
    .X(_08211_));
 sky130_fd_sc_hd__o211a_1 _15081_ (.A1(_08189_),
    .A2(_08209_),
    .B1(_08210_),
    .C1(_08211_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _15082_ (.A0(\rbzero.wall_tracer.trackDistY[8] ),
    .A1(\rbzero.wall_tracer.trackDistX[8] ),
    .S(_08190_),
    .X(_08212_));
 sky130_fd_sc_hd__or2_1 _15083_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08165_),
    .X(_08213_));
 sky130_fd_sc_hd__o211a_1 _15084_ (.A1(_08189_),
    .A2(_08212_),
    .B1(_08213_),
    .C1(_08211_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _15085_ (.A0(\rbzero.wall_tracer.trackDistY[9] ),
    .A1(\rbzero.wall_tracer.trackDistX[9] ),
    .S(_06178_),
    .X(_08214_));
 sky130_fd_sc_hd__or2_1 _15086_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_08165_),
    .X(_08215_));
 sky130_fd_sc_hd__o211a_1 _15087_ (.A1(_08160_),
    .A2(_08214_),
    .B1(_08215_),
    .C1(_08211_),
    .X(_00433_));
 sky130_fd_sc_hd__o21a_1 _15088_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(_06177_),
    .B1(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_08216_));
 sky130_fd_sc_hd__inv_2 _15089_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_1 _15090_ (.A(_08217_),
    .B(_08160_),
    .Y(_08218_));
 sky130_fd_sc_hd__o211a_1 _15091_ (.A1(_08160_),
    .A2(_08216_),
    .B1(_08218_),
    .C1(_08211_),
    .X(_00434_));
 sky130_fd_sc_hd__and4b_2 _15092_ (.A_N(_04571_),
    .B(_04568_),
    .C(_04572_),
    .D(_04570_),
    .X(_08219_));
 sky130_fd_sc_hd__buf_4 _15093_ (.A(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__mux2_1 _15094_ (.A0(\rbzero.wall_tracer.stepDistX[-11] ),
    .A1(_07997_),
    .S(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__clkbuf_1 _15095_ (.A(_08221_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _15096_ (.A0(\rbzero.wall_tracer.stepDistX[-10] ),
    .A1(_08017_),
    .S(_08220_),
    .X(_08222_));
 sky130_fd_sc_hd__clkbuf_1 _15097_ (.A(_08222_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _15098_ (.A0(\rbzero.wall_tracer.stepDistX[-9] ),
    .A1(_08033_),
    .S(_08220_),
    .X(_08223_));
 sky130_fd_sc_hd__clkbuf_1 _15099_ (.A(_08223_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _15100_ (.A0(\rbzero.wall_tracer.stepDistX[-8] ),
    .A1(_08050_),
    .S(_08220_),
    .X(_08224_));
 sky130_fd_sc_hd__clkbuf_1 _15101_ (.A(_08224_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _15102_ (.A0(\rbzero.wall_tracer.stepDistX[-7] ),
    .A1(_08064_),
    .S(_08220_),
    .X(_08225_));
 sky130_fd_sc_hd__clkbuf_1 _15103_ (.A(_08225_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _15104_ (.A0(\rbzero.wall_tracer.stepDistX[-6] ),
    .A1(_08074_),
    .S(_08220_),
    .X(_08226_));
 sky130_fd_sc_hd__clkbuf_1 _15105_ (.A(_08226_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _15106_ (.A0(\rbzero.wall_tracer.stepDistX[-5] ),
    .A1(_08085_),
    .S(_08220_),
    .X(_08227_));
 sky130_fd_sc_hd__clkbuf_1 _15107_ (.A(_08227_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _15108_ (.A0(\rbzero.wall_tracer.stepDistX[-4] ),
    .A1(_08094_),
    .S(_08220_),
    .X(_08228_));
 sky130_fd_sc_hd__clkbuf_1 _15109_ (.A(_08228_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _15110_ (.A0(\rbzero.wall_tracer.stepDistX[-3] ),
    .A1(_08100_),
    .S(_08220_),
    .X(_08229_));
 sky130_fd_sc_hd__clkbuf_1 _15111_ (.A(_08229_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _15112_ (.A0(\rbzero.wall_tracer.stepDistX[-2] ),
    .A1(_08104_),
    .S(_08220_),
    .X(_08230_));
 sky130_fd_sc_hd__clkbuf_1 _15113_ (.A(_08230_),
    .X(_00444_));
 sky130_fd_sc_hd__buf_4 _15114_ (.A(_08219_),
    .X(_08231_));
 sky130_fd_sc_hd__mux2_1 _15115_ (.A0(\rbzero.wall_tracer.stepDistX[-1] ),
    .A1(_08111_),
    .S(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__clkbuf_1 _15116_ (.A(_08232_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _15117_ (.A0(\rbzero.wall_tracer.stepDistX[0] ),
    .A1(_08117_),
    .S(_08231_),
    .X(_08233_));
 sky130_fd_sc_hd__clkbuf_1 _15118_ (.A(_08233_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _15119_ (.A0(\rbzero.wall_tracer.stepDistX[1] ),
    .A1(_08121_),
    .S(_08231_),
    .X(_08234_));
 sky130_fd_sc_hd__clkbuf_1 _15120_ (.A(_08234_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _15121_ (.A0(\rbzero.wall_tracer.stepDistX[2] ),
    .A1(_08126_),
    .S(_08231_),
    .X(_08235_));
 sky130_fd_sc_hd__clkbuf_1 _15122_ (.A(_08235_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _15123_ (.A0(\rbzero.wall_tracer.stepDistX[3] ),
    .A1(_08134_),
    .S(_08231_),
    .X(_08236_));
 sky130_fd_sc_hd__clkbuf_1 _15124_ (.A(_08236_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _15125_ (.A0(\rbzero.wall_tracer.stepDistX[4] ),
    .A1(_08140_),
    .S(_08231_),
    .X(_08237_));
 sky130_fd_sc_hd__clkbuf_1 _15126_ (.A(_08237_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _15127_ (.A0(\rbzero.wall_tracer.stepDistX[5] ),
    .A1(_08142_),
    .S(_08231_),
    .X(_08238_));
 sky130_fd_sc_hd__clkbuf_1 _15128_ (.A(_08238_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _15129_ (.A0(\rbzero.wall_tracer.stepDistX[6] ),
    .A1(_08145_),
    .S(_08231_),
    .X(_08239_));
 sky130_fd_sc_hd__clkbuf_1 _15130_ (.A(_08239_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _15131_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_08149_),
    .S(_08231_),
    .X(_08240_));
 sky130_fd_sc_hd__clkbuf_1 _15132_ (.A(_08240_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _15133_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_08153_),
    .S(_08231_),
    .X(_08241_));
 sky130_fd_sc_hd__clkbuf_1 _15134_ (.A(_08241_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _15135_ (.A0(\rbzero.wall_tracer.stepDistX[9] ),
    .A1(_08155_),
    .S(_08219_),
    .X(_08242_));
 sky130_fd_sc_hd__clkbuf_1 _15136_ (.A(_08242_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _15137_ (.A0(\rbzero.wall_tracer.stepDistX[10] ),
    .A1(_08157_),
    .S(_08219_),
    .X(_08243_));
 sky130_fd_sc_hd__clkbuf_1 _15138_ (.A(_08243_),
    .X(_00456_));
 sky130_fd_sc_hd__buf_4 _15139_ (.A(_04108_),
    .X(_08244_));
 sky130_fd_sc_hd__clkbuf_8 _15140_ (.A(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__buf_4 _15141_ (.A(_08245_),
    .X(_08246_));
 sky130_fd_sc_hd__and2_1 _15142_ (.A(_08246_),
    .B(_05181_),
    .X(_08247_));
 sky130_fd_sc_hd__clkbuf_1 _15143_ (.A(_08247_),
    .X(_00457_));
 sky130_fd_sc_hd__nor2_1 _15144_ (.A(net64),
    .B(_05409_),
    .Y(_00458_));
 sky130_fd_sc_hd__and2_1 _15145_ (.A(_08246_),
    .B(_05493_),
    .X(_08248_));
 sky130_fd_sc_hd__clkbuf_1 _15146_ (.A(_08248_),
    .X(_00459_));
 sky130_fd_sc_hd__buf_4 _15147_ (.A(_08245_),
    .X(_08249_));
 sky130_fd_sc_hd__and2_1 _15148_ (.A(_08249_),
    .B(_05573_),
    .X(_08250_));
 sky130_fd_sc_hd__clkbuf_1 _15149_ (.A(_08250_),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _15150_ (.A(_08249_),
    .B(_05647_),
    .X(_08251_));
 sky130_fd_sc_hd__clkbuf_1 _15151_ (.A(_08251_),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _15152_ (.A(_08249_),
    .B(_05725_),
    .X(_08252_));
 sky130_fd_sc_hd__clkbuf_1 _15153_ (.A(_08252_),
    .X(_00462_));
 sky130_fd_sc_hd__clkinv_2 _15154_ (.A(_06283_),
    .Y(_08253_));
 sky130_fd_sc_hd__nor2_1 _15155_ (.A(_06218_),
    .B(_06265_),
    .Y(_08254_));
 sky130_fd_sc_hd__inv_2 _15156_ (.A(_06280_),
    .Y(_08255_));
 sky130_fd_sc_hd__a22o_1 _15157_ (.A1(\rbzero.mapdyw[0] ),
    .A2(_08254_),
    .B1(_08255_),
    .B2(_06248_),
    .X(_08256_));
 sky130_fd_sc_hd__mux2_1 _15158_ (.A0(_08256_),
    .A1(\rbzero.mapdxw[0] ),
    .S(_06228_),
    .X(_08257_));
 sky130_fd_sc_hd__and2_2 _15159_ (.A(_04568_),
    .B(_06282_),
    .X(_08258_));
 sky130_fd_sc_hd__a22o_1 _15160_ (.A1(_04592_),
    .A2(_08253_),
    .B1(_08257_),
    .B2(_08258_),
    .X(_00463_));
 sky130_fd_sc_hd__a22o_1 _15161_ (.A1(\rbzero.mapdyw[1] ),
    .A2(_08254_),
    .B1(_08255_),
    .B2(_06256_),
    .X(_08259_));
 sky130_fd_sc_hd__mux2_1 _15162_ (.A0(_08259_),
    .A1(\rbzero.mapdxw[1] ),
    .S(_06228_),
    .X(_08260_));
 sky130_fd_sc_hd__a22o_1 _15163_ (.A1(\rbzero.wall_hot[1] ),
    .A2(_08253_),
    .B1(_08258_),
    .B2(_08260_),
    .X(_00464_));
 sky130_fd_sc_hd__clkbuf_4 _15164_ (.A(_04566_),
    .X(_08261_));
 sky130_fd_sc_hd__buf_4 _15165_ (.A(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__buf_4 _15166_ (.A(_04618_),
    .X(_08263_));
 sky130_fd_sc_hd__nor2_1 _15167_ (.A(_06178_),
    .B(_08159_),
    .Y(_08264_));
 sky130_fd_sc_hd__a21oi_1 _15168_ (.A1(_08263_),
    .A2(_08160_),
    .B1(_08264_),
    .Y(_08265_));
 sky130_fd_sc_hd__nor2_1 _15169_ (.A(_08262_),
    .B(_08265_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _15170_ (.A(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .Y(_08266_));
 sky130_fd_sc_hd__nor2_1 _15171_ (.A(_04564_),
    .B(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__buf_4 _15172_ (.A(_08267_),
    .X(_08268_));
 sky130_fd_sc_hd__clkbuf_4 _15173_ (.A(_08268_),
    .X(_08269_));
 sky130_fd_sc_hd__buf_4 _15174_ (.A(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__and2b_1 _15175_ (.A_N(_08263_),
    .B(\rbzero.debug_overlay.playerY[-6] ),
    .X(_08271_));
 sky130_fd_sc_hd__a21oi_1 _15176_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_08263_),
    .B1(_08271_),
    .Y(_08272_));
 sky130_fd_sc_hd__or2_1 _15177_ (.A(\rbzero.trace_state[0] ),
    .B(_06097_),
    .X(_08273_));
 sky130_fd_sc_hd__buf_6 _15178_ (.A(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__xor2_2 _15179_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(\rbzero.debug_overlay.playerX[-9] ),
    .X(_08275_));
 sky130_fd_sc_hd__or3_1 _15180_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .B(_06491_),
    .C(_06514_),
    .X(_08276_));
 sky130_fd_sc_hd__nand2_1 _15181_ (.A(_06424_),
    .B(_06500_),
    .Y(_08277_));
 sky130_fd_sc_hd__and4bb_1 _15182_ (.A_N(\rbzero.wall_tracer.rayAddendX[-2] ),
    .B_N(_08276_),
    .C(_08277_),
    .D(_06507_),
    .X(_08278_));
 sky130_fd_sc_hd__and4_1 _15183_ (.A(_06477_),
    .B(_06482_),
    .C(_06486_),
    .D(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__and4bb_1 _15184_ (.A_N(_06521_),
    .B_N(_06473_),
    .C(_08279_),
    .D(_06528_),
    .X(_08280_));
 sky130_fd_sc_hd__a31o_2 _15185_ (.A1(_06466_),
    .A2(_06454_),
    .A3(_08280_),
    .B1(_06552_),
    .X(_08281_));
 sky130_fd_sc_hd__mux2_2 _15186_ (.A0(_08275_),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__xor2_1 _15187_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(\rbzero.debug_overlay.playerY[-9] ),
    .X(_08283_));
 sky130_fd_sc_hd__mux2_1 _15188_ (.A0(_08283_),
    .A1(\rbzero.debug_overlay.playerY[-8] ),
    .S(_06370_),
    .X(_08284_));
 sky130_fd_sc_hd__and2_2 _15189_ (.A(\rbzero.trace_state[1] ),
    .B(_06096_),
    .X(_08285_));
 sky130_fd_sc_hd__or2_1 _15190_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__nand2_4 _15191_ (.A(\rbzero.trace_state[0] ),
    .B(_08285_),
    .Y(_08287_));
 sky130_fd_sc_hd__mux2_1 _15192_ (.A0(_08284_),
    .A1(_08286_),
    .S(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__o21ai_4 _15193_ (.A1(_08274_),
    .A2(_08282_),
    .B1(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__buf_2 _15194_ (.A(_08289_),
    .X(_08290_));
 sky130_fd_sc_hd__buf_6 _15195_ (.A(_08274_),
    .X(_08291_));
 sky130_fd_sc_hd__buf_6 _15196_ (.A(_08291_),
    .X(_08292_));
 sky130_fd_sc_hd__and3_2 _15197_ (.A(_04570_),
    .B(\rbzero.trace_state[0] ),
    .C(_06096_),
    .X(_08293_));
 sky130_fd_sc_hd__buf_4 _15198_ (.A(_08293_),
    .X(_08294_));
 sky130_fd_sc_hd__o31a_4 _15199_ (.A1(_07995_),
    .A2(_08104_),
    .A3(_08110_),
    .B1(_08117_),
    .X(_08295_));
 sky130_fd_sc_hd__nor4_1 _15200_ (.A(_07996_),
    .B(_08104_),
    .C(_08110_),
    .D(_08117_),
    .Y(_08296_));
 sky130_fd_sc_hd__or2_1 _15201_ (.A(_04564_),
    .B(_08266_),
    .X(_08297_));
 sky130_fd_sc_hd__buf_4 _15202_ (.A(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__o21ai_1 _15203_ (.A1(_08295_),
    .A2(_08296_),
    .B1(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__nand2_1 _15204_ (.A(_04617_),
    .B(_06521_),
    .Y(_08300_));
 sky130_fd_sc_hd__o211a_1 _15205_ (.A1(_04617_),
    .A2(_06346_),
    .B1(_08268_),
    .C1(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__nor2_1 _15206_ (.A(_08294_),
    .B(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__a22o_4 _15207_ (.A1(\rbzero.wall_tracer.stepDistY[0] ),
    .A2(_08294_),
    .B1(_08299_),
    .B2(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__and2_1 _15208_ (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .B(_06099_),
    .X(_08304_));
 sky130_fd_sc_hd__a21oi_2 _15209_ (.A1(_08292_),
    .A2(_08303_),
    .B1(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__nor2_1 _15210_ (.A(_08290_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__or3_1 _15211_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(\rbzero.debug_overlay.playerX[-8] ),
    .C(\rbzero.debug_overlay.playerX[-9] ),
    .X(_08307_));
 sky130_fd_sc_hd__o21ai_1 _15212_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(\rbzero.debug_overlay.playerX[-9] ),
    .B1(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_08308_));
 sky130_fd_sc_hd__and2_1 _15213_ (.A(_08307_),
    .B(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__mux2_2 _15214_ (.A0(_08309_),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_08281_),
    .X(_08310_));
 sky130_fd_sc_hd__or3_1 _15215_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(\rbzero.debug_overlay.playerY[-8] ),
    .C(\rbzero.debug_overlay.playerY[-9] ),
    .X(_08311_));
 sky130_fd_sc_hd__o21ai_1 _15216_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(\rbzero.debug_overlay.playerY[-9] ),
    .B1(\rbzero.debug_overlay.playerY[-7] ),
    .Y(_08312_));
 sky130_fd_sc_hd__and2_1 _15217_ (.A(_08311_),
    .B(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__mux2_1 _15218_ (.A0(_08313_),
    .A1(\rbzero.debug_overlay.playerY[-7] ),
    .S(_06370_),
    .X(_08314_));
 sky130_fd_sc_hd__or2_1 _15219_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(_08285_),
    .X(_08315_));
 sky130_fd_sc_hd__mux2_1 _15220_ (.A0(_08314_),
    .A1(_08315_),
    .S(_08287_),
    .X(_08316_));
 sky130_fd_sc_hd__o21ai_4 _15221_ (.A1(_08274_),
    .A2(_08310_),
    .B1(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__clkbuf_4 _15222_ (.A(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__buf_6 _15223_ (.A(_06097_),
    .X(_08319_));
 sky130_fd_sc_hd__xor2_1 _15224_ (.A(_08104_),
    .B(_08111_),
    .X(_08320_));
 sky130_fd_sc_hd__nor2_1 _15225_ (.A(_04616_),
    .B(_06349_),
    .Y(_08321_));
 sky130_fd_sc_hd__a211o_1 _15226_ (.A1(_04617_),
    .A2(_06528_),
    .B1(_08298_),
    .C1(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__o21ai_4 _15227_ (.A1(_08268_),
    .A2(_08320_),
    .B1(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__buf_4 _15228_ (.A(_08285_),
    .X(_08324_));
 sky130_fd_sc_hd__and3_2 _15229_ (.A(\rbzero.trace_state[0] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .C(_08324_),
    .X(_08325_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .B(_06099_),
    .Y(_08326_));
 sky130_fd_sc_hd__inv_2 _15231_ (.A(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__a211oi_4 _15232_ (.A1(_08319_),
    .A2(_08323_),
    .B1(_08325_),
    .C1(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__nor2_1 _15233_ (.A(_08318_),
    .B(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__xnor2_1 _15234_ (.A(_08306_),
    .B(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__or2_1 _15235_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08307_),
    .X(_08331_));
 sky130_fd_sc_hd__nand2_1 _15236_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08307_),
    .Y(_08332_));
 sky130_fd_sc_hd__and2_1 _15237_ (.A(_08331_),
    .B(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__clkbuf_4 _15238_ (.A(_08281_),
    .X(_08334_));
 sky130_fd_sc_hd__mux2_1 _15239_ (.A0(_08333_),
    .A1(\rbzero.debug_overlay.playerX[-6] ),
    .S(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__or2_1 _15240_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08311_),
    .X(_08336_));
 sky130_fd_sc_hd__nand2_1 _15241_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08311_),
    .Y(_08337_));
 sky130_fd_sc_hd__and2_1 _15242_ (.A(_08336_),
    .B(_08337_),
    .X(_08338_));
 sky130_fd_sc_hd__mux2_1 _15243_ (.A0(_08338_),
    .A1(\rbzero.debug_overlay.playerY[-6] ),
    .S(_06370_),
    .X(_08339_));
 sky130_fd_sc_hd__or2_1 _15244_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(_08324_),
    .X(_08340_));
 sky130_fd_sc_hd__buf_4 _15245_ (.A(_08287_),
    .X(_08341_));
 sky130_fd_sc_hd__mux2_1 _15246_ (.A0(_08339_),
    .A1(_08340_),
    .S(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__o21ai_4 _15247_ (.A1(_08291_),
    .A2(_08335_),
    .B1(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__clkbuf_4 _15248_ (.A(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__nand2_1 _15249_ (.A(_04616_),
    .B(_06473_),
    .Y(_08345_));
 sky130_fd_sc_hd__o211a_1 _15250_ (.A1(_04616_),
    .A2(_06367_),
    .B1(_08268_),
    .C1(_08345_),
    .X(_08346_));
 sky130_fd_sc_hd__a211oi_4 _15251_ (.A1(_08104_),
    .A2(_08298_),
    .B1(_08346_),
    .C1(_08324_),
    .Y(_08347_));
 sky130_fd_sc_hd__a21oi_1 _15252_ (.A1(\rbzero.wall_tracer.stepDistY[-2] ),
    .A2(_08293_),
    .B1(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__clkbuf_4 _15253_ (.A(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__a21boi_2 _15254_ (.A1(\rbzero.wall_tracer.stepDistX[-2] ),
    .A2(_06099_),
    .B1_N(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__buf_2 _15255_ (.A(_08350_),
    .X(_08351_));
 sky130_fd_sc_hd__nor2_1 _15256_ (.A(_08344_),
    .B(_08351_),
    .Y(_08352_));
 sky130_fd_sc_hd__xnor2_1 _15257_ (.A(_08330_),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__buf_4 _15258_ (.A(_08324_),
    .X(_08354_));
 sky130_fd_sc_hd__buf_6 _15259_ (.A(_08298_),
    .X(_08355_));
 sky130_fd_sc_hd__xnor2_1 _15260_ (.A(_08121_),
    .B(_08295_),
    .Y(_08356_));
 sky130_fd_sc_hd__nand2_1 _15261_ (.A(_04618_),
    .B(_06466_),
    .Y(_08357_));
 sky130_fd_sc_hd__o211a_1 _15262_ (.A1(_04618_),
    .A2(_06336_),
    .B1(_08269_),
    .C1(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__a21oi_2 _15263_ (.A1(_08355_),
    .A2(_08356_),
    .B1(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__buf_2 _15264_ (.A(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__a22o_1 _15265_ (.A1(\rbzero.wall_tracer.stepDistX[1] ),
    .A2(_06099_),
    .B1(_08294_),
    .B2(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_08361_));
 sky130_fd_sc_hd__o21ba_2 _15266_ (.A1(_08354_),
    .A2(_08360_),
    .B1_N(_08361_),
    .X(_08362_));
 sky130_fd_sc_hd__clkinv_2 _15267_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_08363_));
 sky130_fd_sc_hd__nor2_2 _15268_ (.A(_08363_),
    .B(_08341_),
    .Y(_08364_));
 sky130_fd_sc_hd__a221oi_4 _15269_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08319_),
    .B1(_06099_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__clkbuf_4 _15270_ (.A(_08365_),
    .X(_08366_));
 sky130_fd_sc_hd__nor2_1 _15271_ (.A(_08362_),
    .B(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__or4_2 _15272_ (.A(_08121_),
    .B(_08126_),
    .C(_08134_),
    .D(_08295_),
    .X(_08368_));
 sky130_fd_sc_hd__o31ai_1 _15273_ (.A1(_08121_),
    .A2(_08126_),
    .A3(_08295_),
    .B1(_08134_),
    .Y(_08369_));
 sky130_fd_sc_hd__mux2_2 _15274_ (.A0(_06329_),
    .A1(_06443_),
    .S(_04617_),
    .X(_08370_));
 sky130_fd_sc_hd__a21o_1 _15275_ (.A1(_08269_),
    .A2(_08370_),
    .B1(_08294_),
    .X(_08371_));
 sky130_fd_sc_hd__a31o_1 _15276_ (.A1(_08355_),
    .A2(_08368_),
    .A3(_08369_),
    .B1(_08371_),
    .X(_08372_));
 sky130_fd_sc_hd__nand2_1 _15277_ (.A(_08164_),
    .B(_08319_),
    .Y(_08373_));
 sky130_fd_sc_hd__buf_2 _15278_ (.A(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__nor2_1 _15279_ (.A(_08372_),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__nor2_1 _15280_ (.A(_04618_),
    .B(_06332_),
    .Y(_08376_));
 sky130_fd_sc_hd__a211o_2 _15281_ (.A1(_04618_),
    .A2(_06454_),
    .B1(_08355_),
    .C1(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__or3_1 _15282_ (.A(_08121_),
    .B(_08126_),
    .C(_08295_),
    .X(_08378_));
 sky130_fd_sc_hd__o21ai_1 _15283_ (.A1(_08121_),
    .A2(_08295_),
    .B1(_08126_),
    .Y(_08379_));
 sky130_fd_sc_hd__a21o_1 _15284_ (.A1(_08378_),
    .A2(_08379_),
    .B1(_08269_),
    .X(_08380_));
 sky130_fd_sc_hd__nand2_1 _15285_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_06097_),
    .Y(_08381_));
 sky130_fd_sc_hd__buf_2 _15286_ (.A(_08381_),
    .X(_08382_));
 sky130_fd_sc_hd__clkbuf_4 _15287_ (.A(_08382_),
    .X(_08383_));
 sky130_fd_sc_hd__a21oi_1 _15288_ (.A1(_08377_),
    .A2(_08380_),
    .B1(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__xnor2_1 _15289_ (.A(_08375_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__xnor2_2 _15290_ (.A(_08367_),
    .B(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__clkbuf_4 _15291_ (.A(_08305_),
    .X(_08387_));
 sky130_fd_sc_hd__nor2_1 _15292_ (.A(_08387_),
    .B(_08366_),
    .Y(_08388_));
 sky130_fd_sc_hd__nor2_1 _15293_ (.A(_08354_),
    .B(_08360_),
    .Y(_08389_));
 sky130_fd_sc_hd__clkbuf_4 _15294_ (.A(_08354_),
    .X(_08390_));
 sky130_fd_sc_hd__a21oi_2 _15295_ (.A1(_08377_),
    .A2(_08380_),
    .B1(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__and2_1 _15296_ (.A(_08164_),
    .B(_08341_),
    .X(_08392_));
 sky130_fd_sc_hd__a22o_1 _15297_ (.A1(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A2(_08389_),
    .B1(_08391_),
    .B2(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__or2_2 _15298_ (.A(_08354_),
    .B(_08359_),
    .X(_08394_));
 sky130_fd_sc_hd__a21o_2 _15299_ (.A1(_08377_),
    .A2(_08380_),
    .B1(_08354_),
    .X(_08395_));
 sky130_fd_sc_hd__nand2_2 _15300_ (.A(_08164_),
    .B(_08287_),
    .Y(_08396_));
 sky130_fd_sc_hd__or4_2 _15301_ (.A(_08169_),
    .B(_08394_),
    .C(_08395_),
    .D(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__a21boi_1 _15302_ (.A1(_08388_),
    .A2(_08393_),
    .B1_N(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__xnor2_1 _15303_ (.A(_08386_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__xnor2_1 _15304_ (.A(_08353_),
    .B(_08399_),
    .Y(_08400_));
 sky130_fd_sc_hd__nand3_1 _15305_ (.A(_08397_),
    .B(_08388_),
    .C(_08393_),
    .Y(_08401_));
 sky130_fd_sc_hd__a21o_1 _15306_ (.A1(_08397_),
    .A2(_08393_),
    .B1(_08388_),
    .X(_08402_));
 sky130_fd_sc_hd__nor2_4 _15307_ (.A(_06099_),
    .B(_08396_),
    .Y(_08403_));
 sky130_fd_sc_hd__nor2_4 _15308_ (.A(_08169_),
    .B(_08354_),
    .Y(_08404_));
 sky130_fd_sc_hd__o2bb2a_1 _15309_ (.A1_N(_08303_),
    .A2_N(_08404_),
    .B1(_08359_),
    .B2(_08374_),
    .X(_08405_));
 sky130_fd_sc_hd__a41o_1 _15310_ (.A1(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A2(_08303_),
    .A3(_08389_),
    .A4(_08403_),
    .B1(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__buf_2 _15311_ (.A(_08328_),
    .X(_08407_));
 sky130_fd_sc_hd__or2_1 _15312_ (.A(_08407_),
    .B(_08366_),
    .X(_08408_));
 sky130_fd_sc_hd__nand2_1 _15313_ (.A(_08303_),
    .B(_08404_),
    .Y(_08409_));
 sky130_fd_sc_hd__or3_1 _15314_ (.A(_08360_),
    .B(_08374_),
    .C(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__o21ai_1 _15315_ (.A1(_08406_),
    .A2(_08408_),
    .B1(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__a21o_1 _15316_ (.A1(_08401_),
    .A2(_08402_),
    .B1(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__clkbuf_4 _15317_ (.A(_08290_),
    .X(_08413_));
 sky130_fd_sc_hd__or2_1 _15318_ (.A(_08318_),
    .B(_08351_),
    .X(_08414_));
 sky130_fd_sc_hd__or3_1 _15319_ (.A(_08413_),
    .B(_08328_),
    .C(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__o21ai_1 _15320_ (.A1(_08413_),
    .A2(_08407_),
    .B1(_08414_),
    .Y(_08416_));
 sky130_fd_sc_hd__nand2_1 _15321_ (.A(_08415_),
    .B(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__a31o_1 _15322_ (.A1(_08062_),
    .A2(_08098_),
    .A3(_08099_),
    .B1(_08268_),
    .X(_08418_));
 sky130_fd_sc_hd__nand2_1 _15323_ (.A(\rbzero.side_hot ),
    .B(_06477_),
    .Y(_08419_));
 sky130_fd_sc_hd__o211a_1 _15324_ (.A1(_04616_),
    .A2(_06342_),
    .B1(_08267_),
    .C1(_08419_),
    .X(_08420_));
 sky130_fd_sc_hd__nor2_1 _15325_ (.A(_08285_),
    .B(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__a2bb2o_4 _15326_ (.A1_N(\rbzero.wall_tracer.stepDistY[-3] ),
    .A2_N(_08287_),
    .B1(_08418_),
    .B2(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__o21bai_4 _15327_ (.A1(\rbzero.wall_tracer.stepDistX[-3] ),
    .A2(_08274_),
    .B1_N(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__buf_2 _15328_ (.A(_08423_),
    .X(_08424_));
 sky130_fd_sc_hd__nor2_1 _15329_ (.A(_08424_),
    .B(_08344_),
    .Y(_08425_));
 sky130_fd_sc_hd__xnor2_1 _15330_ (.A(_08417_),
    .B(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__nand3_1 _15331_ (.A(_08401_),
    .B(_08402_),
    .C(_08411_),
    .Y(_08427_));
 sky130_fd_sc_hd__a21boi_1 _15332_ (.A1(_08412_),
    .A2(_08426_),
    .B1_N(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__nor2_1 _15333_ (.A(_08400_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__and2_1 _15334_ (.A(_08400_),
    .B(_08428_),
    .X(_08430_));
 sky130_fd_sc_hd__nor2_1 _15335_ (.A(_08429_),
    .B(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__a31o_1 _15336_ (.A1(_08062_),
    .A2(_08089_),
    .A3(_08093_),
    .B1(_08268_),
    .X(_08432_));
 sky130_fd_sc_hd__nand2_1 _15337_ (.A(_04616_),
    .B(_06482_),
    .Y(_08433_));
 sky130_fd_sc_hd__o211a_1 _15338_ (.A1(_04616_),
    .A2(_06350_),
    .B1(_08268_),
    .C1(_08433_),
    .X(_08434_));
 sky130_fd_sc_hd__nor2_1 _15339_ (.A(_08324_),
    .B(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__a2bb2o_1 _15340_ (.A1_N(\rbzero.wall_tracer.stepDistY[-4] ),
    .A2_N(_08287_),
    .B1(_08432_),
    .B2(_08435_),
    .X(_08436_));
 sky130_fd_sc_hd__o21bai_4 _15341_ (.A1(\rbzero.wall_tracer.stepDistX[-4] ),
    .A2(_08274_),
    .B1_N(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__inv_2 _15342_ (.A(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_08438_));
 sky130_fd_sc_hd__nand2_1 _15343_ (.A(_04616_),
    .B(_06486_),
    .Y(_08439_));
 sky130_fd_sc_hd__o211a_1 _15344_ (.A1(_04616_),
    .A2(_06352_),
    .B1(_08268_),
    .C1(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__a21oi_2 _15345_ (.A1(_08085_),
    .A2(_08298_),
    .B1(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__nor2_1 _15346_ (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(_08274_),
    .Y(_08442_));
 sky130_fd_sc_hd__a221o_2 _15347_ (.A1(_08438_),
    .A2(_08293_),
    .B1(_08441_),
    .B2(_06097_),
    .C1(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__buf_2 _15348_ (.A(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__xor2_1 _15349_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_08331_),
    .X(_08445_));
 sky130_fd_sc_hd__mux2_1 _15350_ (.A0(_08445_),
    .A1(\rbzero.debug_overlay.playerX[-5] ),
    .S(_08281_),
    .X(_08446_));
 sky130_fd_sc_hd__xor2_1 _15351_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_08336_),
    .X(_08447_));
 sky130_fd_sc_hd__mux2_1 _15352_ (.A0(_08447_),
    .A1(\rbzero.debug_overlay.playerY[-5] ),
    .S(_06370_),
    .X(_08448_));
 sky130_fd_sc_hd__or2_1 _15353_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_08324_),
    .X(_08449_));
 sky130_fd_sc_hd__mux2_1 _15354_ (.A0(_08448_),
    .A1(_08449_),
    .S(_08341_),
    .X(_08450_));
 sky130_fd_sc_hd__o21ai_4 _15355_ (.A1(_08291_),
    .A2(_08446_),
    .B1(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__clkbuf_4 _15356_ (.A(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__or3_1 _15357_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(\rbzero.debug_overlay.playerX[-5] ),
    .C(_08331_),
    .X(_08453_));
 sky130_fd_sc_hd__o21ai_1 _15358_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_08331_),
    .B1(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_08454_));
 sky130_fd_sc_hd__nand2_1 _15359_ (.A(_08453_),
    .B(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__inv_2 _15360_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_08456_));
 sky130_fd_sc_hd__mux2_1 _15361_ (.A0(_08455_),
    .A1(_08456_),
    .S(_08281_),
    .X(_08457_));
 sky130_fd_sc_hd__or3_1 _15362_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .C(_08336_),
    .X(_08458_));
 sky130_fd_sc_hd__o21ai_1 _15363_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_08336_),
    .B1(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_08459_));
 sky130_fd_sc_hd__nand2_1 _15364_ (.A(_08458_),
    .B(_08459_),
    .Y(_08460_));
 sky130_fd_sc_hd__inv_2 _15365_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_08461_));
 sky130_fd_sc_hd__mux2_1 _15366_ (.A0(_08460_),
    .A1(_08461_),
    .S(_06370_),
    .X(_08462_));
 sky130_fd_sc_hd__mux2_1 _15367_ (.A0(_08182_),
    .A1(_08462_),
    .S(_08293_),
    .X(_08463_));
 sky130_fd_sc_hd__mux2_4 _15368_ (.A0(_08457_),
    .A1(_08463_),
    .S(_08274_),
    .X(_08464_));
 sky130_fd_sc_hd__buf_2 _15369_ (.A(_08464_),
    .X(_08465_));
 sky130_fd_sc_hd__or4_1 _15370_ (.A(_08437_),
    .B(_08444_),
    .C(_08452_),
    .D(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__nor2_1 _15371_ (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .B(_08291_),
    .Y(_08467_));
 sky130_fd_sc_hd__o31ai_2 _15372_ (.A1(_07996_),
    .A2(_08071_),
    .A3(_08073_),
    .B1(_08298_),
    .Y(_08468_));
 sky130_fd_sc_hd__mux2_1 _15373_ (.A0(_06356_),
    .A1(_06514_),
    .S(_04617_),
    .X(_08469_));
 sky130_fd_sc_hd__a21oi_1 _15374_ (.A1(_08269_),
    .A2(_08469_),
    .B1(_08324_),
    .Y(_08470_));
 sky130_fd_sc_hd__a2bb2o_2 _15375_ (.A1_N(\rbzero.wall_tracer.stepDistY[-6] ),
    .A2_N(_08341_),
    .B1(_08468_),
    .B2(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__or2_2 _15376_ (.A(_08467_),
    .B(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__buf_2 _15377_ (.A(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__or2_1 _15378_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08453_),
    .X(_08474_));
 sky130_fd_sc_hd__nand2_1 _15379_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08453_),
    .Y(_08475_));
 sky130_fd_sc_hd__and2_1 _15380_ (.A(_08474_),
    .B(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__mux2_2 _15381_ (.A0(_08476_),
    .A1(\rbzero.debug_overlay.playerX[-3] ),
    .S(_08334_),
    .X(_08477_));
 sky130_fd_sc_hd__or2_1 _15382_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08458_),
    .X(_08478_));
 sky130_fd_sc_hd__nand2_1 _15383_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08458_),
    .Y(_08479_));
 sky130_fd_sc_hd__and2_1 _15384_ (.A(_08478_),
    .B(_08479_),
    .X(_08480_));
 sky130_fd_sc_hd__mux2_1 _15385_ (.A0(_08480_),
    .A1(\rbzero.debug_overlay.playerY[-3] ),
    .S(_06370_),
    .X(_08481_));
 sky130_fd_sc_hd__or2_1 _15386_ (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .B(_08354_),
    .X(_08482_));
 sky130_fd_sc_hd__mux2_1 _15387_ (.A0(_08481_),
    .A1(_08482_),
    .S(_08341_),
    .X(_08483_));
 sky130_fd_sc_hd__o21ai_4 _15388_ (.A1(_08292_),
    .A2(_08477_),
    .B1(_08483_),
    .Y(_08484_));
 sky130_fd_sc_hd__buf_2 _15389_ (.A(_08484_),
    .X(_08485_));
 sky130_fd_sc_hd__buf_2 _15390_ (.A(_08437_),
    .X(_08486_));
 sky130_fd_sc_hd__buf_4 _15391_ (.A(_08465_),
    .X(_08487_));
 sky130_fd_sc_hd__o22ai_1 _15392_ (.A1(_08486_),
    .A2(_08452_),
    .B1(_08487_),
    .B2(_08444_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand2_1 _15393_ (.A(_08466_),
    .B(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__or3_1 _15394_ (.A(_08473_),
    .B(_08485_),
    .C(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__nand2_1 _15395_ (.A(_08466_),
    .B(_08490_),
    .Y(_08491_));
 sky130_fd_sc_hd__clkbuf_4 _15396_ (.A(_08344_),
    .X(_08492_));
 sky130_fd_sc_hd__o31a_1 _15397_ (.A1(_08424_),
    .A2(_08492_),
    .A3(_08417_),
    .B1(_08415_),
    .X(_08493_));
 sky130_fd_sc_hd__or4_1 _15398_ (.A(_08424_),
    .B(_08486_),
    .C(_08452_),
    .D(_08465_),
    .X(_08494_));
 sky130_fd_sc_hd__clkbuf_4 _15399_ (.A(_08452_),
    .X(_08495_));
 sky130_fd_sc_hd__o22ai_1 _15400_ (.A1(_08424_),
    .A2(_08495_),
    .B1(_08487_),
    .B2(_08486_),
    .Y(_08496_));
 sky130_fd_sc_hd__or4bb_1 _15401_ (.A(_08444_),
    .B(_08485_),
    .C_N(_08494_),
    .D_N(_08496_),
    .X(_08497_));
 sky130_fd_sc_hd__a2bb2o_1 _15402_ (.A1_N(_08444_),
    .A2_N(_08485_),
    .B1(_08494_),
    .B2(_08496_),
    .X(_08498_));
 sky130_fd_sc_hd__nand2_1 _15403_ (.A(_08497_),
    .B(_08498_),
    .Y(_08499_));
 sky130_fd_sc_hd__xnor2_1 _15404_ (.A(_08493_),
    .B(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__xnor2_1 _15405_ (.A(_08491_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__xnor2_1 _15406_ (.A(_08431_),
    .B(_08501_),
    .Y(_08502_));
 sky130_fd_sc_hd__nand2_1 _15407_ (.A(_08427_),
    .B(_08412_),
    .Y(_08503_));
 sky130_fd_sc_hd__xor2_2 _15408_ (.A(_08503_),
    .B(_08426_),
    .X(_08504_));
 sky130_fd_sc_hd__nor2_1 _15409_ (.A(_08328_),
    .B(_08366_),
    .Y(_08505_));
 sky130_fd_sc_hd__xnor2_1 _15410_ (.A(_08406_),
    .B(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__a22o_1 _15411_ (.A1(_08303_),
    .A2(_08403_),
    .B1(_08404_),
    .B2(_08323_),
    .X(_08507_));
 sky130_fd_sc_hd__nor2_1 _15412_ (.A(_08350_),
    .B(_08365_),
    .Y(_08508_));
 sky130_fd_sc_hd__a21oi_4 _15413_ (.A1(_08319_),
    .A2(_08323_),
    .B1(_08325_),
    .Y(_08509_));
 sky130_fd_sc_hd__or3_1 _15414_ (.A(_08509_),
    .B(_08396_),
    .C(_08409_),
    .X(_08510_));
 sky130_fd_sc_hd__a21boi_2 _15415_ (.A1(_08507_),
    .A2(_08508_),
    .B1_N(_08510_),
    .Y(_08511_));
 sky130_fd_sc_hd__xnor2_1 _15416_ (.A(_08506_),
    .B(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__nor2_1 _15417_ (.A(_08423_),
    .B(_08317_),
    .Y(_08513_));
 sky130_fd_sc_hd__nor2_1 _15418_ (.A(_08290_),
    .B(_08350_),
    .Y(_08514_));
 sky130_fd_sc_hd__xnor2_1 _15419_ (.A(_08513_),
    .B(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__or3_1 _15420_ (.A(_08486_),
    .B(_08344_),
    .C(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__o21ai_1 _15421_ (.A1(_08486_),
    .A2(_08344_),
    .B1(_08515_),
    .Y(_08517_));
 sky130_fd_sc_hd__and2_1 _15422_ (.A(_08516_),
    .B(_08517_),
    .X(_08518_));
 sky130_fd_sc_hd__or2b_1 _15423_ (.A(_08511_),
    .B_N(_08506_),
    .X(_08519_));
 sky130_fd_sc_hd__a21boi_1 _15424_ (.A1(_08512_),
    .A2(_08518_),
    .B1_N(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__xor2_1 _15425_ (.A(_08504_),
    .B(_08520_),
    .X(_08521_));
 sky130_fd_sc_hd__o22ai_1 _15426_ (.A1(_08444_),
    .A2(_08452_),
    .B1(_08473_),
    .B2(_08465_),
    .Y(_08522_));
 sky130_fd_sc_hd__or2_2 _15427_ (.A(\rbzero.wall_tracer.stepDistY[-7] ),
    .B(_08341_),
    .X(_08523_));
 sky130_fd_sc_hd__nand2_1 _15428_ (.A(_04617_),
    .B(_06507_),
    .Y(_08524_));
 sky130_fd_sc_hd__o211a_1 _15429_ (.A1(_04617_),
    .A2(_06360_),
    .B1(_08268_),
    .C1(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__a211o_2 _15430_ (.A1(_08064_),
    .A2(_08298_),
    .B1(_08525_),
    .C1(_08354_),
    .X(_08526_));
 sky130_fd_sc_hd__o211ai_4 _15431_ (.A1(\rbzero.wall_tracer.stepDistX[-7] ),
    .A2(_08291_),
    .B1(_08523_),
    .C1(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__clkbuf_4 _15432_ (.A(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__nor2_1 _15433_ (.A(_08528_),
    .B(_08485_),
    .Y(_08529_));
 sky130_fd_sc_hd__or4_1 _15434_ (.A(_08443_),
    .B(_08451_),
    .C(_08472_),
    .D(_08465_),
    .X(_08530_));
 sky130_fd_sc_hd__a21bo_1 _15435_ (.A1(_08522_),
    .A2(_08529_),
    .B1_N(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__nand2_1 _15436_ (.A(_08513_),
    .B(_08514_),
    .Y(_08532_));
 sky130_fd_sc_hd__clkbuf_4 _15437_ (.A(_08485_),
    .X(_08533_));
 sky130_fd_sc_hd__o21ai_1 _15438_ (.A1(_08473_),
    .A2(_08533_),
    .B1(_08489_),
    .Y(_08534_));
 sky130_fd_sc_hd__nand2_1 _15439_ (.A(_08490_),
    .B(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__a21o_1 _15440_ (.A1(_08532_),
    .A2(_08516_),
    .B1(_08535_),
    .X(_08536_));
 sky130_fd_sc_hd__nand3_1 _15441_ (.A(_08532_),
    .B(_08516_),
    .C(_08535_),
    .Y(_08537_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(_08536_),
    .B(_08537_),
    .Y(_08538_));
 sky130_fd_sc_hd__xnor2_1 _15443_ (.A(_08531_),
    .B(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__nor2_1 _15444_ (.A(_08504_),
    .B(_08520_),
    .Y(_08540_));
 sky130_fd_sc_hd__a21oi_1 _15445_ (.A1(_08521_),
    .A2(_08539_),
    .B1(_08540_),
    .Y(_08541_));
 sky130_fd_sc_hd__xor2_1 _15446_ (.A(_08502_),
    .B(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__buf_6 _15447_ (.A(_08319_),
    .X(_08543_));
 sky130_fd_sc_hd__nand2_4 _15448_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__clkbuf_4 _15449_ (.A(_08544_),
    .X(_08545_));
 sky130_fd_sc_hd__mux2_1 _15450_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(_04617_),
    .X(_08546_));
 sky130_fd_sc_hd__a21o_1 _15451_ (.A1(_08269_),
    .A2(_08546_),
    .B1(_08294_),
    .X(_08547_));
 sky130_fd_sc_hd__a21o_2 _15452_ (.A1(_07997_),
    .A2(_08298_),
    .B1(_08547_),
    .X(_08548_));
 sky130_fd_sc_hd__o211ai_4 _15453_ (.A1(\rbzero.wall_tracer.stepDistY[-11] ),
    .A2(_08319_),
    .B1(_08291_),
    .C1(_08548_),
    .Y(_08549_));
 sky130_fd_sc_hd__clkbuf_4 _15454_ (.A(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__mux2_1 _15455_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(_04616_),
    .X(_08551_));
 sky130_fd_sc_hd__or2_1 _15456_ (.A(_08298_),
    .B(_08551_),
    .X(_08552_));
 sky130_fd_sc_hd__o211a_4 _15457_ (.A1(_08017_),
    .A2(_08268_),
    .B1(_08552_),
    .C1(_08341_),
    .X(_08553_));
 sky130_fd_sc_hd__buf_4 _15458_ (.A(_08341_),
    .X(_08554_));
 sky130_fd_sc_hd__nand2_1 _15459_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__nor2_2 _15460_ (.A(_06101_),
    .B(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__nand2_1 _15461_ (.A(_08553_),
    .B(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__or3_2 _15462_ (.A(_08545_),
    .B(_08550_),
    .C(_08557_),
    .X(_08558_));
 sky130_fd_sc_hd__a21o_1 _15463_ (.A1(\rbzero.wall_tracer.stepDistY[-10] ),
    .A2(_08324_),
    .B1(_06098_),
    .X(_08559_));
 sky130_fd_sc_hd__nor2_2 _15464_ (.A(_08553_),
    .B(_08559_),
    .Y(_08560_));
 sky130_fd_sc_hd__clkbuf_4 _15465_ (.A(_08560_),
    .X(_08561_));
 sky130_fd_sc_hd__a2bb2o_1 _15466_ (.A1_N(_08545_),
    .A2_N(_08561_),
    .B1(_08548_),
    .B2(_08556_),
    .X(_08562_));
 sky130_fd_sc_hd__or2_1 _15467_ (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .B(_08291_),
    .X(_08563_));
 sky130_fd_sc_hd__or2_1 _15468_ (.A(\rbzero.wall_tracer.stepDistY[-8] ),
    .B(_08341_),
    .X(_08564_));
 sky130_fd_sc_hd__mux2_1 _15469_ (.A0(_06358_),
    .A1(_06491_),
    .S(_04617_),
    .X(_08565_));
 sky130_fd_sc_hd__a21o_1 _15470_ (.A1(_08269_),
    .A2(_08565_),
    .B1(_08324_),
    .X(_08566_));
 sky130_fd_sc_hd__a21o_2 _15471_ (.A1(_08050_),
    .A2(_08298_),
    .B1(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__nand3_1 _15472_ (.A(_08563_),
    .B(_08564_),
    .C(_08567_),
    .Y(_08568_));
 sky130_fd_sc_hd__clkbuf_4 _15473_ (.A(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__or3_4 _15474_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .B(\rbzero.debug_overlay.playerX[-2] ),
    .C(_08474_),
    .X(_08570_));
 sky130_fd_sc_hd__o21ai_1 _15475_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_08474_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_08571_));
 sky130_fd_sc_hd__nand2_2 _15476_ (.A(_08570_),
    .B(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__mux2_1 _15477_ (.A0(_08572_),
    .A1(_04862_),
    .S(_08334_),
    .X(_08573_));
 sky130_fd_sc_hd__or3_4 _15478_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .C(_08478_),
    .X(_08574_));
 sky130_fd_sc_hd__o21ai_1 _15479_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_08478_),
    .B1(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_08575_));
 sky130_fd_sc_hd__and2_1 _15480_ (.A(_08574_),
    .B(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__mux2_1 _15481_ (.A0(_08576_),
    .A1(\rbzero.debug_overlay.playerY[-1] ),
    .S(_06370_),
    .X(_08577_));
 sky130_fd_sc_hd__nand2_1 _15482_ (.A(_08294_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__a21oi_1 _15483_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_08319_),
    .B1(_06099_),
    .Y(_08579_));
 sky130_fd_sc_hd__a22o_4 _15484_ (.A1(_06099_),
    .A2(_08573_),
    .B1(_08578_),
    .B2(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__xor2_1 _15485_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_08478_),
    .X(_08581_));
 sky130_fd_sc_hd__mux2_1 _15486_ (.A0(_08581_),
    .A1(\rbzero.debug_overlay.playerY[-2] ),
    .S(_06370_),
    .X(_08582_));
 sky130_fd_sc_hd__mux2_1 _15487_ (.A0(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A1(_08582_),
    .S(_08294_),
    .X(_08583_));
 sky130_fd_sc_hd__xnor2_2 _15488_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_08474_),
    .Y(_08584_));
 sky130_fd_sc_hd__or2_1 _15489_ (.A(_08334_),
    .B(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__a21oi_1 _15490_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_08334_),
    .B1(_08291_),
    .Y(_08586_));
 sky130_fd_sc_hd__a2bb2o_4 _15491_ (.A1_N(_06100_),
    .A2_N(_08583_),
    .B1(_08585_),
    .B2(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__or2_1 _15492_ (.A(_08528_),
    .B(_08587_),
    .X(_08588_));
 sky130_fd_sc_hd__or3_1 _15493_ (.A(_08569_),
    .B(_08580_),
    .C(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__clkbuf_4 _15494_ (.A(_08580_),
    .X(_08590_));
 sky130_fd_sc_hd__o21ai_1 _15495_ (.A1(_08569_),
    .A2(_08590_),
    .B1(_08588_),
    .Y(_08591_));
 sky130_fd_sc_hd__nand2_1 _15496_ (.A(_08589_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__nor2_1 _15497_ (.A(\rbzero.wall_tracer.stepDistX[-9] ),
    .B(_08274_),
    .Y(_08593_));
 sky130_fd_sc_hd__nand2_1 _15498_ (.A(\rbzero.side_hot ),
    .B(_08277_),
    .Y(_08594_));
 sky130_fd_sc_hd__o211a_1 _15499_ (.A1(\rbzero.side_hot ),
    .A2(_06361_),
    .B1(_08267_),
    .C1(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__a211o_1 _15500_ (.A1(_08033_),
    .A2(_08297_),
    .B1(_08595_),
    .C1(_08324_),
    .X(_08596_));
 sky130_fd_sc_hd__o21ai_2 _15501_ (.A1(\rbzero.wall_tracer.stepDistY[-9] ),
    .A2(_08287_),
    .B1(_08596_),
    .Y(_08597_));
 sky130_fd_sc_hd__or2_1 _15502_ (.A(_08593_),
    .B(_08597_),
    .X(_08598_));
 sky130_fd_sc_hd__clkbuf_4 _15503_ (.A(_08598_),
    .X(_08599_));
 sky130_fd_sc_hd__o32a_1 _15504_ (.A1(_06370_),
    .A2(_08554_),
    .A3(_08574_),
    .B1(_08354_),
    .B2(_08194_),
    .X(_08600_));
 sky130_fd_sc_hd__o31a_4 _15505_ (.A1(_08292_),
    .A2(_08334_),
    .A3(_08570_),
    .B1(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__buf_2 _15506_ (.A(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__or2_1 _15507_ (.A(_08599_),
    .B(_08602_),
    .X(_08603_));
 sky130_fd_sc_hd__xnor2_1 _15508_ (.A(_08592_),
    .B(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__or2_1 _15509_ (.A(_08569_),
    .B(_08587_),
    .X(_08605_));
 sky130_fd_sc_hd__or2_1 _15510_ (.A(_08580_),
    .B(_08599_),
    .X(_08606_));
 sky130_fd_sc_hd__o22ai_4 _15511_ (.A1(\rbzero.wall_tracer.stepDistX[-10] ),
    .A2(_08291_),
    .B1(_08553_),
    .B2(_08559_),
    .Y(_08607_));
 sky130_fd_sc_hd__nor2_1 _15512_ (.A(_08601_),
    .B(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__xor2_1 _15513_ (.A(_08605_),
    .B(_08606_),
    .X(_08609_));
 sky130_fd_sc_hd__a2bb2oi_1 _15514_ (.A1_N(_08605_),
    .A2_N(_08606_),
    .B1(_08608_),
    .B2(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__nor2_1 _15515_ (.A(_08604_),
    .B(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__and2_1 _15516_ (.A(_08604_),
    .B(_08610_),
    .X(_08612_));
 sky130_fd_sc_hd__nor2_1 _15517_ (.A(_08611_),
    .B(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__a31o_1 _15518_ (.A1(_08558_),
    .A2(_08562_),
    .A3(_08613_),
    .B1(_08611_),
    .X(_08614_));
 sky130_fd_sc_hd__or2b_1 _15519_ (.A(_08538_),
    .B_N(_08531_),
    .X(_08615_));
 sky130_fd_sc_hd__clkbuf_4 _15520_ (.A(_08597_),
    .X(_08616_));
 sky130_fd_sc_hd__nor2_1 _15521_ (.A(_08544_),
    .B(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__xnor2_1 _15522_ (.A(_08557_),
    .B(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__nand2_1 _15523_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08543_),
    .Y(_08619_));
 sky130_fd_sc_hd__buf_2 _15524_ (.A(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__nor2_1 _15525_ (.A(_08549_),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__nand2_1 _15526_ (.A(_08618_),
    .B(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__or2_1 _15527_ (.A(_08618_),
    .B(_08621_),
    .X(_08623_));
 sky130_fd_sc_hd__and2_1 _15528_ (.A(_08622_),
    .B(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__or2_1 _15529_ (.A(_08569_),
    .B(_08601_),
    .X(_08625_));
 sky130_fd_sc_hd__o22ai_1 _15530_ (.A1(_08473_),
    .A2(_08587_),
    .B1(_08580_),
    .B2(_08528_),
    .Y(_08626_));
 sky130_fd_sc_hd__or3_1 _15531_ (.A(_08473_),
    .B(_08580_),
    .C(_08588_),
    .X(_08627_));
 sky130_fd_sc_hd__nand3b_1 _15532_ (.A_N(_08625_),
    .B(_08626_),
    .C(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__a21bo_1 _15533_ (.A1(_08627_),
    .A2(_08626_),
    .B1_N(_08625_),
    .X(_08629_));
 sky130_fd_sc_hd__nand2_1 _15534_ (.A(_08628_),
    .B(_08629_),
    .Y(_08630_));
 sky130_fd_sc_hd__o31a_1 _15535_ (.A1(_08592_),
    .A2(_08599_),
    .A3(_08602_),
    .B1(_08589_),
    .X(_08631_));
 sky130_fd_sc_hd__xor2_1 _15536_ (.A(_08630_),
    .B(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__nand2_1 _15537_ (.A(_08624_),
    .B(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__or2_1 _15538_ (.A(_08624_),
    .B(_08632_),
    .X(_08634_));
 sky130_fd_sc_hd__nand2_1 _15539_ (.A(_08633_),
    .B(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__a21o_1 _15540_ (.A1(_08536_),
    .A2(_08615_),
    .B1(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__nand3_1 _15541_ (.A(_08536_),
    .B(_08615_),
    .C(_08635_),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_1 _15542_ (.A(_08636_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__xnor2_1 _15543_ (.A(_08614_),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__xnor2_1 _15544_ (.A(_08542_),
    .B(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__xnor2_1 _15545_ (.A(_08521_),
    .B(_08539_),
    .Y(_08641_));
 sky130_fd_sc_hd__xnor2_1 _15546_ (.A(_08512_),
    .B(_08518_),
    .Y(_08642_));
 sky130_fd_sc_hd__o31a_1 _15547_ (.A1(_08509_),
    .A2(_08396_),
    .A3(_08409_),
    .B1(_08507_),
    .X(_08643_));
 sky130_fd_sc_hd__xnor2_2 _15548_ (.A(_08643_),
    .B(_08508_),
    .Y(_08644_));
 sky130_fd_sc_hd__or4bb_1 _15549_ (.A(_08381_),
    .B(_08348_),
    .C_N(_08323_),
    .D_N(_08392_),
    .X(_08645_));
 sky130_fd_sc_hd__nor2_1 _15550_ (.A(_08169_),
    .B(_08294_),
    .Y(_08646_));
 sky130_fd_sc_hd__a22o_1 _15551_ (.A1(_08323_),
    .A2(_08403_),
    .B1(_08646_),
    .B2(_08347_),
    .X(_08647_));
 sky130_fd_sc_hd__or4bb_1 _15552_ (.A(_08423_),
    .B(_08365_),
    .C_N(_08645_),
    .D_N(_08647_),
    .X(_08648_));
 sky130_fd_sc_hd__and2_1 _15553_ (.A(_08645_),
    .B(_08648_),
    .X(_08649_));
 sky130_fd_sc_hd__xor2_1 _15554_ (.A(_08644_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__or4_1 _15555_ (.A(_08423_),
    .B(_08317_),
    .C(_08289_),
    .D(_08437_),
    .X(_08651_));
 sky130_fd_sc_hd__o22ai_1 _15556_ (.A1(_08423_),
    .A2(_08290_),
    .B1(_08437_),
    .B2(_08317_),
    .Y(_08652_));
 sky130_fd_sc_hd__nand2_1 _15557_ (.A(_08651_),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__or3_1 _15558_ (.A(_08653_),
    .B(_08343_),
    .C(_08443_),
    .X(_08654_));
 sky130_fd_sc_hd__o21ai_1 _15559_ (.A1(_08343_),
    .A2(_08444_),
    .B1(_08653_),
    .Y(_08655_));
 sky130_fd_sc_hd__and2_1 _15560_ (.A(_08654_),
    .B(_08655_),
    .X(_08656_));
 sky130_fd_sc_hd__nor2_1 _15561_ (.A(_08644_),
    .B(_08649_),
    .Y(_08657_));
 sky130_fd_sc_hd__a21o_1 _15562_ (.A1(_08650_),
    .A2(_08656_),
    .B1(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__xnor2_1 _15563_ (.A(_08642_),
    .B(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__o22a_1 _15564_ (.A1(_08451_),
    .A2(_08472_),
    .B1(_08464_),
    .B2(_08527_),
    .X(_08660_));
 sky130_fd_sc_hd__or2_1 _15565_ (.A(_08484_),
    .B(_08569_),
    .X(_08661_));
 sky130_fd_sc_hd__or4_1 _15566_ (.A(_08495_),
    .B(_08473_),
    .C(_08487_),
    .D(_08528_),
    .X(_08662_));
 sky130_fd_sc_hd__o21ai_1 _15567_ (.A1(_08660_),
    .A2(_08661_),
    .B1(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__nand2_1 _15568_ (.A(_08530_),
    .B(_08522_),
    .Y(_08664_));
 sky130_fd_sc_hd__xor2_1 _15569_ (.A(_08664_),
    .B(_08529_),
    .X(_08665_));
 sky130_fd_sc_hd__a21o_1 _15570_ (.A1(_08651_),
    .A2(_08654_),
    .B1(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__nand3_1 _15571_ (.A(_08651_),
    .B(_08654_),
    .C(_08665_),
    .Y(_08667_));
 sky130_fd_sc_hd__nand2_1 _15572_ (.A(_08666_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__xnor2_1 _15573_ (.A(_08663_),
    .B(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__and2b_1 _15574_ (.A_N(_08642_),
    .B(_08658_),
    .X(_08670_));
 sky130_fd_sc_hd__a21oi_1 _15575_ (.A1(_08659_),
    .A2(_08669_),
    .B1(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__xor2_1 _15576_ (.A(_08641_),
    .B(_08671_),
    .X(_08672_));
 sky130_fd_sc_hd__xnor2_1 _15577_ (.A(_08608_),
    .B(_08609_),
    .Y(_08673_));
 sky130_fd_sc_hd__buf_4 _15578_ (.A(_08587_),
    .X(_08674_));
 sky130_fd_sc_hd__buf_2 _15579_ (.A(_08607_),
    .X(_08675_));
 sky130_fd_sc_hd__a21boi_2 _15580_ (.A1(\rbzero.wall_tracer.stepDistX[-11] ),
    .A2(_06100_),
    .B1_N(_08549_),
    .Y(_08676_));
 sky130_fd_sc_hd__or2_1 _15581_ (.A(_08601_),
    .B(_08676_),
    .X(_08677_));
 sky130_fd_sc_hd__o22ai_1 _15582_ (.A1(_08587_),
    .A2(_08599_),
    .B1(_08607_),
    .B2(_08580_),
    .Y(_08678_));
 sky130_fd_sc_hd__o31a_1 _15583_ (.A1(_08587_),
    .A2(_08606_),
    .A3(_08607_),
    .B1(_08678_),
    .X(_08679_));
 sky130_fd_sc_hd__or2b_1 _15584_ (.A(_08677_),
    .B_N(_08679_),
    .X(_08680_));
 sky130_fd_sc_hd__o31a_1 _15585_ (.A1(_08674_),
    .A2(_08606_),
    .A3(_08675_),
    .B1(_08680_),
    .X(_08681_));
 sky130_fd_sc_hd__xor2_1 _15586_ (.A(_08673_),
    .B(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__or3b_2 _15587_ (.A(_08545_),
    .B(_08550_),
    .C_N(_08682_),
    .X(_08683_));
 sky130_fd_sc_hd__o21ai_1 _15588_ (.A1(_08673_),
    .A2(_08681_),
    .B1(_08683_),
    .Y(_08684_));
 sky130_fd_sc_hd__a21bo_1 _15589_ (.A1(_08663_),
    .A2(_08667_),
    .B1_N(_08666_),
    .X(_08685_));
 sky130_fd_sc_hd__nand2_1 _15590_ (.A(_08558_),
    .B(_08562_),
    .Y(_08686_));
 sky130_fd_sc_hd__xor2_1 _15591_ (.A(_08686_),
    .B(_08613_),
    .X(_08687_));
 sky130_fd_sc_hd__xor2_1 _15592_ (.A(_08685_),
    .B(_08687_),
    .X(_08688_));
 sky130_fd_sc_hd__xnor2_1 _15593_ (.A(_08684_),
    .B(_08688_),
    .Y(_08689_));
 sky130_fd_sc_hd__nand2_1 _15594_ (.A(_08672_),
    .B(_08689_),
    .Y(_08690_));
 sky130_fd_sc_hd__o21a_1 _15595_ (.A1(_08641_),
    .A2(_08671_),
    .B1(_08690_),
    .X(_08691_));
 sky130_fd_sc_hd__xor2_1 _15596_ (.A(_08640_),
    .B(_08691_),
    .X(_08692_));
 sky130_fd_sc_hd__or2b_1 _15597_ (.A(_08687_),
    .B_N(_08685_),
    .X(_08693_));
 sky130_fd_sc_hd__or2b_1 _15598_ (.A(_08688_),
    .B_N(_08684_),
    .X(_08694_));
 sky130_fd_sc_hd__a21oi_2 _15599_ (.A1(_08693_),
    .A2(_08694_),
    .B1(_08558_),
    .Y(_08695_));
 sky130_fd_sc_hd__and3_1 _15600_ (.A(_08558_),
    .B(_08693_),
    .C(_08694_),
    .X(_08696_));
 sky130_fd_sc_hd__nor2_1 _15601_ (.A(_08695_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__xnor2_1 _15602_ (.A(_08692_),
    .B(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__or2_1 _15603_ (.A(_08672_),
    .B(_08689_),
    .X(_08699_));
 sky130_fd_sc_hd__nand2_1 _15604_ (.A(_08690_),
    .B(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__xnor2_1 _15605_ (.A(_08659_),
    .B(_08669_),
    .Y(_08701_));
 sky130_fd_sc_hd__xnor2_1 _15606_ (.A(_08650_),
    .B(_08656_),
    .Y(_08702_));
 sky130_fd_sc_hd__a2bb2o_1 _15607_ (.A1_N(_08423_),
    .A2_N(_08365_),
    .B1(_08645_),
    .B2(_08647_),
    .X(_08703_));
 sky130_fd_sc_hd__or4_1 _15608_ (.A(_08422_),
    .B(_08348_),
    .C(_08396_),
    .D(_08382_),
    .X(_08704_));
 sky130_fd_sc_hd__o22ai_1 _15609_ (.A1(_08349_),
    .A2(_08396_),
    .B1(_08382_),
    .B2(_08422_),
    .Y(_08705_));
 sky130_fd_sc_hd__or4bb_1 _15610_ (.A(_08437_),
    .B(_08365_),
    .C_N(_08704_),
    .D_N(_08705_),
    .X(_08706_));
 sky130_fd_sc_hd__nand2_1 _15611_ (.A(_08704_),
    .B(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__nand3_1 _15612_ (.A(_08648_),
    .B(_08703_),
    .C(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__or2_1 _15613_ (.A(_08343_),
    .B(_08472_),
    .X(_08709_));
 sky130_fd_sc_hd__nor2_1 _15614_ (.A(_08289_),
    .B(_08443_),
    .Y(_08710_));
 sky130_fd_sc_hd__or3b_1 _15615_ (.A(_08317_),
    .B(_08437_),
    .C_N(_08710_),
    .X(_08711_));
 sky130_fd_sc_hd__a22o_1 _15616_ (.A1(_08438_),
    .A2(_08294_),
    .B1(_08441_),
    .B2(_06097_),
    .X(_08712_));
 sky130_fd_sc_hd__nor2_1 _15617_ (.A(_08442_),
    .B(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__inv_2 _15618_ (.A(_08317_),
    .Y(_08714_));
 sky130_fd_sc_hd__a2bb2o_1 _15619_ (.A1_N(_08289_),
    .A2_N(_08437_),
    .B1(_08713_),
    .B2(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__and2_1 _15620_ (.A(_08711_),
    .B(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__xnor2_1 _15621_ (.A(_08709_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__a21o_1 _15622_ (.A1(_08648_),
    .A2(_08703_),
    .B1(_08707_),
    .X(_08718_));
 sky130_fd_sc_hd__nand3_1 _15623_ (.A(_08708_),
    .B(_08717_),
    .C(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__and2_1 _15624_ (.A(_08708_),
    .B(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__xor2_1 _15625_ (.A(_08702_),
    .B(_08720_),
    .X(_08721_));
 sky130_fd_sc_hd__nor2_1 _15626_ (.A(_08464_),
    .B(_08527_),
    .Y(_08722_));
 sky130_fd_sc_hd__and4b_1 _15627_ (.A_N(_08451_),
    .B(_08563_),
    .C(_08564_),
    .D(_08567_),
    .X(_08723_));
 sky130_fd_sc_hd__nor2_1 _15628_ (.A(_08484_),
    .B(_08599_),
    .Y(_08724_));
 sky130_fd_sc_hd__o22a_1 _15629_ (.A1(_08451_),
    .A2(_08527_),
    .B1(_08568_),
    .B2(_08464_),
    .X(_08725_));
 sky130_fd_sc_hd__a21oi_1 _15630_ (.A1(_08722_),
    .A2(_08723_),
    .B1(_08725_),
    .Y(_08726_));
 sky130_fd_sc_hd__a22o_1 _15631_ (.A1(_08722_),
    .A2(_08723_),
    .B1(_08724_),
    .B2(_08726_),
    .X(_08727_));
 sky130_fd_sc_hd__or2b_1 _15632_ (.A(_08709_),
    .B_N(_08716_),
    .X(_08728_));
 sky130_fd_sc_hd__nor4_1 _15633_ (.A(_08451_),
    .B(_08472_),
    .C(_08464_),
    .D(_08527_),
    .Y(_08729_));
 sky130_fd_sc_hd__nor2_1 _15634_ (.A(_08729_),
    .B(_08660_),
    .Y(_08730_));
 sky130_fd_sc_hd__xor2_1 _15635_ (.A(_08730_),
    .B(_08661_),
    .X(_08731_));
 sky130_fd_sc_hd__a21o_1 _15636_ (.A1(_08711_),
    .A2(_08728_),
    .B1(_08731_),
    .X(_08732_));
 sky130_fd_sc_hd__nand3_1 _15637_ (.A(_08711_),
    .B(_08728_),
    .C(_08731_),
    .Y(_08733_));
 sky130_fd_sc_hd__nand2_1 _15638_ (.A(_08732_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__xnor2_1 _15639_ (.A(_08727_),
    .B(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__nor2_1 _15640_ (.A(_08702_),
    .B(_08720_),
    .Y(_08736_));
 sky130_fd_sc_hd__a21oi_1 _15641_ (.A1(_08721_),
    .A2(_08735_),
    .B1(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__nor2_1 _15642_ (.A(_08701_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__and2_1 _15643_ (.A(_08701_),
    .B(_08737_),
    .X(_08739_));
 sky130_fd_sc_hd__nor2_1 _15644_ (.A(_08738_),
    .B(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__nor2_1 _15645_ (.A(_08674_),
    .B(_08675_),
    .Y(_08741_));
 sky130_fd_sc_hd__clkbuf_4 _15646_ (.A(_08676_),
    .X(_08742_));
 sky130_fd_sc_hd__nor2_1 _15647_ (.A(_08590_),
    .B(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__nand2_1 _15648_ (.A(_08741_),
    .B(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__xnor2_1 _15649_ (.A(_08677_),
    .B(_08679_),
    .Y(_08745_));
 sky130_fd_sc_hd__or2b_1 _15650_ (.A(_08744_),
    .B_N(_08745_),
    .X(_08746_));
 sky130_fd_sc_hd__a21bo_1 _15651_ (.A1(_08727_),
    .A2(_08733_),
    .B1_N(_08732_),
    .X(_08747_));
 sky130_fd_sc_hd__a31o_1 _15652_ (.A1(\rbzero.wall_tracer.visualWallDist[1] ),
    .A2(_08543_),
    .A3(_08548_),
    .B1(_08682_),
    .X(_08748_));
 sky130_fd_sc_hd__nand2_1 _15653_ (.A(_08683_),
    .B(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__xnor2_2 _15654_ (.A(_08747_),
    .B(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__xnor2_1 _15655_ (.A(_08746_),
    .B(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__a21oi_1 _15656_ (.A1(_08740_),
    .A2(_08751_),
    .B1(_08738_),
    .Y(_08752_));
 sky130_fd_sc_hd__xnor2_2 _15657_ (.A(_08700_),
    .B(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__and3_1 _15658_ (.A(_08741_),
    .B(_08743_),
    .C(_08745_),
    .X(_08754_));
 sky130_fd_sc_hd__a32oi_4 _15659_ (.A1(_08683_),
    .A2(_08747_),
    .A3(_08748_),
    .B1(_08750_),
    .B2(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__or2_1 _15660_ (.A(_08700_),
    .B(_08752_),
    .X(_08756_));
 sky130_fd_sc_hd__o21a_1 _15661_ (.A1(_08753_),
    .A2(_08755_),
    .B1(_08756_),
    .X(_08757_));
 sky130_fd_sc_hd__nor2_1 _15662_ (.A(_08698_),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__and2_1 _15663_ (.A(_08698_),
    .B(_08757_),
    .X(_08759_));
 sky130_fd_sc_hd__or2_1 _15664_ (.A(_08758_),
    .B(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__xnor2_1 _15665_ (.A(_08724_),
    .B(_08726_),
    .Y(_08761_));
 sky130_fd_sc_hd__nor2_1 _15666_ (.A(_08317_),
    .B(_08473_),
    .Y(_08762_));
 sky130_fd_sc_hd__or3_1 _15667_ (.A(_08317_),
    .B(_08467_),
    .C(_08471_),
    .X(_08763_));
 sky130_fd_sc_hd__xnor2_1 _15668_ (.A(_08710_),
    .B(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__nor2_1 _15669_ (.A(_08343_),
    .B(_08528_),
    .Y(_08765_));
 sky130_fd_sc_hd__a22o_1 _15670_ (.A1(_08710_),
    .A2(_08762_),
    .B1(_08764_),
    .B2(_08765_),
    .X(_08766_));
 sky130_fd_sc_hd__or2b_1 _15671_ (.A(_08761_),
    .B_N(_08766_),
    .X(_08767_));
 sky130_fd_sc_hd__xor2_1 _15672_ (.A(_08766_),
    .B(_08761_),
    .X(_08768_));
 sky130_fd_sc_hd__nor2_1 _15673_ (.A(_08485_),
    .B(_08607_),
    .Y(_08769_));
 sky130_fd_sc_hd__or3_1 _15674_ (.A(_08464_),
    .B(_08593_),
    .C(_08616_),
    .X(_08770_));
 sky130_fd_sc_hd__xnor2_1 _15675_ (.A(_08723_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__or3_1 _15676_ (.A(_08452_),
    .B(_08569_),
    .C(_08770_),
    .X(_08772_));
 sky130_fd_sc_hd__a21bo_1 _15677_ (.A1(_08769_),
    .A2(_08771_),
    .B1_N(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__or2b_1 _15678_ (.A(_08768_),
    .B_N(_08773_),
    .X(_08774_));
 sky130_fd_sc_hd__a21o_1 _15679_ (.A1(_08741_),
    .A2(_08743_),
    .B1(_08745_),
    .X(_08775_));
 sky130_fd_sc_hd__nand2_1 _15680_ (.A(_08746_),
    .B(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__a21oi_2 _15681_ (.A1(_08767_),
    .A2(_08774_),
    .B1(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__xnor2_1 _15682_ (.A(_08740_),
    .B(_08751_),
    .Y(_08778_));
 sky130_fd_sc_hd__xnor2_1 _15683_ (.A(_08721_),
    .B(_08735_),
    .Y(_08779_));
 sky130_fd_sc_hd__a21o_1 _15684_ (.A1(_08708_),
    .A2(_08718_),
    .B1(_08717_),
    .X(_08780_));
 sky130_fd_sc_hd__a2bb2o_1 _15685_ (.A1_N(_08437_),
    .A2_N(_08365_),
    .B1(_08704_),
    .B2(_08705_),
    .X(_08781_));
 sky130_fd_sc_hd__a221o_4 _15686_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08319_),
    .B1(_06099_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08364_),
    .X(_08782_));
 sky130_fd_sc_hd__clkbuf_4 _15687_ (.A(_08436_),
    .X(_08783_));
 sky130_fd_sc_hd__o22ai_2 _15688_ (.A1(_08422_),
    .A2(_08373_),
    .B1(_08382_),
    .B2(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__and4bb_1 _15689_ (.A_N(_08422_),
    .B_N(_08783_),
    .C(_08403_),
    .D(_08404_),
    .X(_08785_));
 sky130_fd_sc_hd__a31o_1 _15690_ (.A1(_08713_),
    .A2(_08782_),
    .A3(_08784_),
    .B1(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__nand3_1 _15691_ (.A(_08706_),
    .B(_08781_),
    .C(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__xor2_1 _15692_ (.A(_08765_),
    .B(_08764_),
    .X(_08788_));
 sky130_fd_sc_hd__a21o_1 _15693_ (.A1(_08706_),
    .A2(_08781_),
    .B1(_08786_),
    .X(_08789_));
 sky130_fd_sc_hd__nand3_1 _15694_ (.A(_08787_),
    .B(_08788_),
    .C(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__nand2_1 _15695_ (.A(_08787_),
    .B(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__nand3_1 _15696_ (.A(_08719_),
    .B(_08780_),
    .C(_08791_),
    .Y(_08792_));
 sky130_fd_sc_hd__xnor2_1 _15697_ (.A(_08773_),
    .B(_08768_),
    .Y(_08793_));
 sky130_fd_sc_hd__a21o_1 _15698_ (.A1(_08719_),
    .A2(_08780_),
    .B1(_08791_),
    .X(_08794_));
 sky130_fd_sc_hd__nand3_1 _15699_ (.A(_08792_),
    .B(_08793_),
    .C(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__and2_1 _15700_ (.A(_08792_),
    .B(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__xor2_1 _15701_ (.A(_08779_),
    .B(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__and3_1 _15702_ (.A(_08767_),
    .B(_08774_),
    .C(_08776_),
    .X(_08798_));
 sky130_fd_sc_hd__nor2_1 _15703_ (.A(_08777_),
    .B(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__nor2_1 _15704_ (.A(_08779_),
    .B(_08796_),
    .Y(_08800_));
 sky130_fd_sc_hd__a21oi_1 _15705_ (.A1(_08797_),
    .A2(_08799_),
    .B1(_08800_),
    .Y(_08801_));
 sky130_fd_sc_hd__xor2_1 _15706_ (.A(_08778_),
    .B(_08801_),
    .X(_08802_));
 sky130_fd_sc_hd__xnor2_1 _15707_ (.A(_08777_),
    .B(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__nor2_1 _15708_ (.A(_08290_),
    .B(_08528_),
    .Y(_08804_));
 sky130_fd_sc_hd__or3_1 _15709_ (.A(_08289_),
    .B(_08467_),
    .C(_08471_),
    .X(_08805_));
 sky130_fd_sc_hd__o2111a_1 _15710_ (.A1(\rbzero.wall_tracer.stepDistX[-7] ),
    .A2(_08291_),
    .B1(_08714_),
    .C1(_08523_),
    .D1(_08526_),
    .X(_08806_));
 sky130_fd_sc_hd__xnor2_1 _15711_ (.A(_08805_),
    .B(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__nor2_1 _15712_ (.A(_08343_),
    .B(_08569_),
    .Y(_08808_));
 sky130_fd_sc_hd__a22o_1 _15713_ (.A1(_08762_),
    .A2(_08804_),
    .B1(_08807_),
    .B2(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__or2_1 _15714_ (.A(_08484_),
    .B(_08607_),
    .X(_08810_));
 sky130_fd_sc_hd__xnor2_1 _15715_ (.A(_08810_),
    .B(_08771_),
    .Y(_08811_));
 sky130_fd_sc_hd__nand2_1 _15716_ (.A(_08809_),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__xnor2_1 _15717_ (.A(_08809_),
    .B(_08811_),
    .Y(_08813_));
 sky130_fd_sc_hd__or3_1 _15718_ (.A(_08451_),
    .B(_08607_),
    .C(_08770_),
    .X(_08814_));
 sky130_fd_sc_hd__o22ai_1 _15719_ (.A1(_08451_),
    .A2(_08599_),
    .B1(_08607_),
    .B2(_08465_),
    .Y(_08815_));
 sky130_fd_sc_hd__or4bb_1 _15720_ (.A(_08484_),
    .B(_08676_),
    .C_N(_08814_),
    .D_N(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__nand2_1 _15721_ (.A(_08814_),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__or2b_1 _15722_ (.A(_08813_),
    .B_N(_08817_),
    .X(_08818_));
 sky130_fd_sc_hd__or2_1 _15723_ (.A(_08741_),
    .B(_08743_),
    .X(_08819_));
 sky130_fd_sc_hd__nand2_1 _15724_ (.A(_08744_),
    .B(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__a21oi_1 _15725_ (.A1(_08812_),
    .A2(_08818_),
    .B1(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__xnor2_1 _15726_ (.A(_08797_),
    .B(_08799_),
    .Y(_08822_));
 sky130_fd_sc_hd__a21o_1 _15727_ (.A1(_08792_),
    .A2(_08794_),
    .B1(_08793_),
    .X(_08823_));
 sky130_fd_sc_hd__a21o_1 _15728_ (.A1(_08787_),
    .A2(_08789_),
    .B1(_08788_),
    .X(_08824_));
 sky130_fd_sc_hd__xor2_1 _15729_ (.A(_08808_),
    .B(_08807_),
    .X(_08825_));
 sky130_fd_sc_hd__or4b_1 _15730_ (.A(_08443_),
    .B(_08365_),
    .C(_08785_),
    .D_N(_08784_),
    .X(_08826_));
 sky130_fd_sc_hd__or4_1 _15731_ (.A(_08422_),
    .B(_08783_),
    .C(_08373_),
    .D(_08382_),
    .X(_08827_));
 sky130_fd_sc_hd__a22o_1 _15732_ (.A1(_08713_),
    .A2(_08782_),
    .B1(_08827_),
    .B2(_08784_),
    .X(_08828_));
 sky130_fd_sc_hd__clkbuf_4 _15733_ (.A(_08712_),
    .X(_08829_));
 sky130_fd_sc_hd__o22a_1 _15734_ (.A1(_08783_),
    .A2(_08373_),
    .B1(_08382_),
    .B2(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__or4_1 _15735_ (.A(_08783_),
    .B(_08712_),
    .C(_08373_),
    .D(_08382_),
    .X(_08831_));
 sky130_fd_sc_hd__o31ai_1 _15736_ (.A1(_08472_),
    .A2(_08365_),
    .A3(_08830_),
    .B1(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__a21o_1 _15737_ (.A1(_08826_),
    .A2(_08828_),
    .B1(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__and3_1 _15738_ (.A(_08826_),
    .B(_08828_),
    .C(_08832_),
    .X(_08834_));
 sky130_fd_sc_hd__a21o_1 _15739_ (.A1(_08825_),
    .A2(_08833_),
    .B1(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__nand3_1 _15740_ (.A(_08790_),
    .B(_08824_),
    .C(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__xnor2_1 _15741_ (.A(_08817_),
    .B(_08813_),
    .Y(_08837_));
 sky130_fd_sc_hd__a21o_1 _15742_ (.A1(_08790_),
    .A2(_08824_),
    .B1(_08835_),
    .X(_08838_));
 sky130_fd_sc_hd__nand3_1 _15743_ (.A(_08836_),
    .B(_08837_),
    .C(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__nand2_1 _15744_ (.A(_08836_),
    .B(_08839_),
    .Y(_08840_));
 sky130_fd_sc_hd__a21o_1 _15745_ (.A1(_08795_),
    .A2(_08823_),
    .B1(_08840_),
    .X(_08841_));
 sky130_fd_sc_hd__and3_1 _15746_ (.A(_08812_),
    .B(_08818_),
    .C(_08820_),
    .X(_08842_));
 sky130_fd_sc_hd__nor2_1 _15747_ (.A(_08821_),
    .B(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__nand3_1 _15748_ (.A(_08795_),
    .B(_08823_),
    .C(_08840_),
    .Y(_08844_));
 sky130_fd_sc_hd__a21boi_1 _15749_ (.A1(_08841_),
    .A2(_08843_),
    .B1_N(_08844_),
    .Y(_08845_));
 sky130_fd_sc_hd__xor2_1 _15750_ (.A(_08822_),
    .B(_08845_),
    .X(_08846_));
 sky130_fd_sc_hd__nor2_1 _15751_ (.A(_08822_),
    .B(_08845_),
    .Y(_08847_));
 sky130_fd_sc_hd__a21oi_1 _15752_ (.A1(_08821_),
    .A2(_08846_),
    .B1(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__nor2_1 _15753_ (.A(_08803_),
    .B(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__xnor2_2 _15754_ (.A(_08753_),
    .B(_08755_),
    .Y(_08850_));
 sky130_fd_sc_hd__nor2_1 _15755_ (.A(_08778_),
    .B(_08801_),
    .Y(_08851_));
 sky130_fd_sc_hd__a21oi_2 _15756_ (.A1(_08777_),
    .A2(_08802_),
    .B1(_08851_),
    .Y(_08852_));
 sky130_fd_sc_hd__xor2_2 _15757_ (.A(_08850_),
    .B(_08852_),
    .X(_08853_));
 sky130_fd_sc_hd__nand2_1 _15758_ (.A(_08849_),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__xnor2_1 _15759_ (.A(_08821_),
    .B(_08846_),
    .Y(_08855_));
 sky130_fd_sc_hd__buf_4 _15760_ (.A(_08674_),
    .X(_08856_));
 sky130_fd_sc_hd__or2_1 _15761_ (.A(_08856_),
    .B(_08742_),
    .X(_08857_));
 sky130_fd_sc_hd__clkbuf_4 _15762_ (.A(_08487_),
    .X(_08858_));
 sky130_fd_sc_hd__nor2_1 _15763_ (.A(_08317_),
    .B(_08569_),
    .Y(_08859_));
 sky130_fd_sc_hd__xor2_1 _15764_ (.A(_08804_),
    .B(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(_08343_),
    .B(_08599_),
    .Y(_08861_));
 sky130_fd_sc_hd__a22o_1 _15766_ (.A1(_08804_),
    .A2(_08859_),
    .B1(_08860_),
    .B2(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__a2bb2o_1 _15767_ (.A1_N(_08484_),
    .A2_N(_08676_),
    .B1(_08814_),
    .B2(_08815_),
    .X(_08863_));
 sky130_fd_sc_hd__and2_1 _15768_ (.A(_08816_),
    .B(_08863_),
    .X(_08864_));
 sky130_fd_sc_hd__nand2_1 _15769_ (.A(_08862_),
    .B(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__or2_1 _15770_ (.A(_08862_),
    .B(_08864_),
    .X(_08866_));
 sky130_fd_sc_hd__nand2_1 _15771_ (.A(_08865_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__clkbuf_4 _15772_ (.A(_08495_),
    .X(_08868_));
 sky130_fd_sc_hd__or2_1 _15773_ (.A(_08868_),
    .B(_08742_),
    .X(_08869_));
 sky130_fd_sc_hd__o41a_1 _15774_ (.A1(_08858_),
    .A2(_08675_),
    .A3(_08867_),
    .A4(_08869_),
    .B1(_08865_),
    .X(_08870_));
 sky130_fd_sc_hd__nor2_1 _15775_ (.A(_08857_),
    .B(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__and3_1 _15776_ (.A(_08844_),
    .B(_08841_),
    .C(_08843_),
    .X(_08872_));
 sky130_fd_sc_hd__a21oi_1 _15777_ (.A1(_08844_),
    .A2(_08841_),
    .B1(_08843_),
    .Y(_08873_));
 sky130_fd_sc_hd__or2_1 _15778_ (.A(_08872_),
    .B(_08873_),
    .X(_08874_));
 sky130_fd_sc_hd__and2_1 _15779_ (.A(_08857_),
    .B(_08870_),
    .X(_08875_));
 sky130_fd_sc_hd__nor2_1 _15780_ (.A(_08871_),
    .B(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__a21o_1 _15781_ (.A1(_08836_),
    .A2(_08838_),
    .B1(_08837_),
    .X(_08877_));
 sky130_fd_sc_hd__nand2_1 _15782_ (.A(_08839_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__inv_2 _15783_ (.A(_08834_),
    .Y(_08879_));
 sky130_fd_sc_hd__nand3_1 _15784_ (.A(_08879_),
    .B(_08825_),
    .C(_08833_),
    .Y(_08880_));
 sky130_fd_sc_hd__a21o_1 _15785_ (.A1(_08879_),
    .A2(_08833_),
    .B1(_08825_),
    .X(_08881_));
 sky130_fd_sc_hd__xor2_1 _15786_ (.A(_08861_),
    .B(_08860_),
    .X(_08882_));
 sky130_fd_sc_hd__or2_1 _15787_ (.A(_08472_),
    .B(_08365_),
    .X(_08883_));
 sky130_fd_sc_hd__nor2_1 _15788_ (.A(_08783_),
    .B(_08382_),
    .Y(_08884_));
 sky130_fd_sc_hd__nor2_1 _15789_ (.A(_08829_),
    .B(_08374_),
    .Y(_08885_));
 sky130_fd_sc_hd__a21o_1 _15790_ (.A1(_08884_),
    .A2(_08885_),
    .B1(_08830_),
    .X(_08886_));
 sky130_fd_sc_hd__xnor2_1 _15791_ (.A(_08883_),
    .B(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__clkbuf_4 _15792_ (.A(_08471_),
    .X(_08888_));
 sky130_fd_sc_hd__nor2_1 _15793_ (.A(_08888_),
    .B(_08382_),
    .Y(_08889_));
 sky130_fd_sc_hd__nor2_1 _15794_ (.A(_08885_),
    .B(_08889_),
    .Y(_08890_));
 sky130_fd_sc_hd__or4_1 _15795_ (.A(_08829_),
    .B(_08471_),
    .C(_08374_),
    .D(_08382_),
    .X(_08891_));
 sky130_fd_sc_hd__o31a_1 _15796_ (.A1(_08528_),
    .A2(_08365_),
    .A3(_08890_),
    .B1(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__nor2_1 _15797_ (.A(_08887_),
    .B(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__and2_1 _15798_ (.A(_08887_),
    .B(_08892_),
    .X(_08894_));
 sky130_fd_sc_hd__nor2_1 _15799_ (.A(_08893_),
    .B(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__a21o_1 _15800_ (.A1(_08882_),
    .A2(_08895_),
    .B1(_08893_),
    .X(_08896_));
 sky130_fd_sc_hd__nor2_1 _15801_ (.A(_08495_),
    .B(_08675_),
    .Y(_08897_));
 sky130_fd_sc_hd__nor2_1 _15802_ (.A(_08487_),
    .B(_08742_),
    .Y(_08898_));
 sky130_fd_sc_hd__and2_1 _15803_ (.A(_08897_),
    .B(_08898_),
    .X(_08899_));
 sky130_fd_sc_hd__xnor2_1 _15804_ (.A(_08867_),
    .B(_08899_),
    .Y(_08900_));
 sky130_fd_sc_hd__nand2_1 _15805_ (.A(_08880_),
    .B(_08881_),
    .Y(_08901_));
 sky130_fd_sc_hd__xnor2_1 _15806_ (.A(_08901_),
    .B(_08896_),
    .Y(_08902_));
 sky130_fd_sc_hd__a32o_1 _15807_ (.A1(_08880_),
    .A2(_08881_),
    .A3(_08896_),
    .B1(_08900_),
    .B2(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__xnor2_1 _15808_ (.A(_08878_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__and3_1 _15809_ (.A(_08839_),
    .B(_08877_),
    .C(_08903_),
    .X(_08905_));
 sky130_fd_sc_hd__a21oi_1 _15810_ (.A1(_08876_),
    .A2(_08904_),
    .B1(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__xor2_1 _15811_ (.A(_08874_),
    .B(_08906_),
    .X(_08907_));
 sky130_fd_sc_hd__nor2_1 _15812_ (.A(_08874_),
    .B(_08906_),
    .Y(_08908_));
 sky130_fd_sc_hd__a21oi_1 _15813_ (.A1(_08871_),
    .A2(_08907_),
    .B1(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__nor2_1 _15814_ (.A(_08855_),
    .B(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__xor2_1 _15815_ (.A(_08803_),
    .B(_08848_),
    .X(_08911_));
 sky130_fd_sc_hd__and2_1 _15816_ (.A(_08910_),
    .B(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__xor2_1 _15817_ (.A(_08855_),
    .B(_08909_),
    .X(_08913_));
 sky130_fd_sc_hd__xor2_1 _15818_ (.A(_08871_),
    .B(_08907_),
    .X(_08914_));
 sky130_fd_sc_hd__xnor2_1 _15819_ (.A(_08900_),
    .B(_08902_),
    .Y(_08915_));
 sky130_fd_sc_hd__xnor2_1 _15820_ (.A(_08882_),
    .B(_08895_),
    .Y(_08916_));
 sky130_fd_sc_hd__nor2_1 _15821_ (.A(_08528_),
    .B(_08366_),
    .Y(_08917_));
 sky130_fd_sc_hd__o21a_1 _15822_ (.A1(_08885_),
    .A2(_08889_),
    .B1(_08891_),
    .X(_08918_));
 sky130_fd_sc_hd__xnor2_1 _15823_ (.A(_08917_),
    .B(_08918_),
    .Y(_08919_));
 sky130_fd_sc_hd__or2_1 _15824_ (.A(_08569_),
    .B(_08366_),
    .X(_08920_));
 sky130_fd_sc_hd__nand2_1 _15825_ (.A(_08523_),
    .B(_08526_),
    .Y(_08921_));
 sky130_fd_sc_hd__clkbuf_4 _15826_ (.A(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__o22a_1 _15827_ (.A1(_08888_),
    .A2(_08374_),
    .B1(_08383_),
    .B2(_08922_),
    .X(_08923_));
 sky130_fd_sc_hd__or3b_1 _15828_ (.A(_08921_),
    .B(_08374_),
    .C_N(_08889_),
    .X(_08924_));
 sky130_fd_sc_hd__o21a_1 _15829_ (.A1(_08920_),
    .A2(_08923_),
    .B1(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__nor2_1 _15830_ (.A(_08919_),
    .B(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__and2_1 _15831_ (.A(_08919_),
    .B(_08925_),
    .X(_08927_));
 sky130_fd_sc_hd__nor2_1 _15832_ (.A(_08926_),
    .B(_08927_),
    .Y(_08928_));
 sky130_fd_sc_hd__or2_1 _15833_ (.A(_08344_),
    .B(_08675_),
    .X(_08929_));
 sky130_fd_sc_hd__or2_1 _15834_ (.A(_08290_),
    .B(_08569_),
    .X(_08930_));
 sky130_fd_sc_hd__or2_1 _15835_ (.A(_08318_),
    .B(_08599_),
    .X(_08931_));
 sky130_fd_sc_hd__xor2_1 _15836_ (.A(_08930_),
    .B(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__xnor2_1 _15837_ (.A(_08929_),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__a21oi_1 _15838_ (.A1(_08928_),
    .A2(_08933_),
    .B1(_08926_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand2_1 _15839_ (.A(_08916_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__or2_1 _15840_ (.A(_08930_),
    .B(_08931_),
    .X(_08936_));
 sky130_fd_sc_hd__or2b_1 _15841_ (.A(_08929_),
    .B_N(_08932_),
    .X(_08937_));
 sky130_fd_sc_hd__xnor2_1 _15842_ (.A(_08897_),
    .B(_08898_),
    .Y(_08938_));
 sky130_fd_sc_hd__a21oi_1 _15843_ (.A1(_08936_),
    .A2(_08937_),
    .B1(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__and3_1 _15844_ (.A(_08936_),
    .B(_08937_),
    .C(_08938_),
    .X(_08940_));
 sky130_fd_sc_hd__nor2_1 _15845_ (.A(_08939_),
    .B(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__nor2_1 _15846_ (.A(_08916_),
    .B(_08934_),
    .Y(_08942_));
 sky130_fd_sc_hd__a21oi_1 _15847_ (.A1(_08935_),
    .A2(_08941_),
    .B1(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__or2_1 _15848_ (.A(_08915_),
    .B(_08943_),
    .X(_08944_));
 sky130_fd_sc_hd__xor2_1 _15849_ (.A(_08915_),
    .B(_08943_),
    .X(_08945_));
 sky130_fd_sc_hd__nand2_1 _15850_ (.A(_08939_),
    .B(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__xnor2_1 _15851_ (.A(_08876_),
    .B(_08904_),
    .Y(_08947_));
 sky130_fd_sc_hd__a21o_1 _15852_ (.A1(_08944_),
    .A2(_08946_),
    .B1(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__inv_2 _15853_ (.A(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__and2_1 _15854_ (.A(_08914_),
    .B(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__and2_1 _15855_ (.A(_08913_),
    .B(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__xor2_1 _15856_ (.A(_08913_),
    .B(_08950_),
    .X(_08952_));
 sky130_fd_sc_hd__nand2_1 _15857_ (.A(_08947_),
    .B(_08944_),
    .Y(_08953_));
 sky130_fd_sc_hd__and2b_1 _15858_ (.A_N(_08942_),
    .B(_08935_),
    .X(_08954_));
 sky130_fd_sc_hd__xnor2_1 _15859_ (.A(_08954_),
    .B(_08941_),
    .Y(_08955_));
 sky130_fd_sc_hd__xnor2_1 _15860_ (.A(_08928_),
    .B(_08933_),
    .Y(_08956_));
 sky130_fd_sc_hd__o22ai_1 _15861_ (.A1(_08413_),
    .A2(_08599_),
    .B1(_08607_),
    .B2(_08318_),
    .Y(_08957_));
 sky130_fd_sc_hd__o31a_1 _15862_ (.A1(_08413_),
    .A2(_08675_),
    .A3(_08931_),
    .B1(_08957_),
    .X(_08958_));
 sky130_fd_sc_hd__or3b_1 _15863_ (.A(_08492_),
    .B(_08742_),
    .C_N(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__o21bai_1 _15864_ (.A1(_08492_),
    .A2(_08742_),
    .B1_N(_08958_),
    .Y(_08960_));
 sky130_fd_sc_hd__and2_1 _15865_ (.A(_08959_),
    .B(_08960_),
    .X(_08961_));
 sky130_fd_sc_hd__clkinv_2 _15866_ (.A(_08922_),
    .Y(_08962_));
 sky130_fd_sc_hd__a31oi_1 _15867_ (.A1(_08962_),
    .A2(_08403_),
    .A3(_08889_),
    .B1(_08923_),
    .Y(_08963_));
 sky130_fd_sc_hd__xor2_1 _15868_ (.A(_08920_),
    .B(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__clkbuf_4 _15869_ (.A(_08366_),
    .X(_08965_));
 sky130_fd_sc_hd__or2_1 _15870_ (.A(_08599_),
    .B(_08965_),
    .X(_08966_));
 sky130_fd_sc_hd__nand2_4 _15871_ (.A(_08564_),
    .B(_08567_),
    .Y(_08967_));
 sky130_fd_sc_hd__or2_1 _15872_ (.A(_08967_),
    .B(_08374_),
    .X(_08968_));
 sky130_fd_sc_hd__or3_1 _15873_ (.A(_08922_),
    .B(_08383_),
    .C(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__o22ai_1 _15874_ (.A1(_08922_),
    .A2(_08374_),
    .B1(_08383_),
    .B2(_08967_),
    .Y(_08970_));
 sky130_fd_sc_hd__nand2_1 _15875_ (.A(_08969_),
    .B(_08970_),
    .Y(_08971_));
 sky130_fd_sc_hd__o21a_1 _15876_ (.A1(_08966_),
    .A2(_08971_),
    .B1(_08969_),
    .X(_08972_));
 sky130_fd_sc_hd__nand2_1 _15877_ (.A(_08964_),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__nor2_1 _15878_ (.A(_08964_),
    .B(_08972_),
    .Y(_08974_));
 sky130_fd_sc_hd__a21oi_1 _15879_ (.A1(_08961_),
    .A2(_08973_),
    .B1(_08974_),
    .Y(_08975_));
 sky130_fd_sc_hd__xor2_1 _15880_ (.A(_08956_),
    .B(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__buf_4 _15881_ (.A(_08290_),
    .X(_08977_));
 sky130_fd_sc_hd__o31a_1 _15882_ (.A1(_08977_),
    .A2(_08675_),
    .A3(_08931_),
    .B1(_08959_),
    .X(_08978_));
 sky130_fd_sc_hd__xor2_1 _15883_ (.A(_08869_),
    .B(_08978_),
    .X(_08979_));
 sky130_fd_sc_hd__nand2_1 _15884_ (.A(_08976_),
    .B(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__o21a_1 _15885_ (.A1(_08956_),
    .A2(_08975_),
    .B1(_08980_),
    .X(_08981_));
 sky130_fd_sc_hd__or2_1 _15886_ (.A(_08955_),
    .B(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__xnor2_1 _15887_ (.A(_08955_),
    .B(_08981_),
    .Y(_08983_));
 sky130_fd_sc_hd__or3_1 _15888_ (.A(_08869_),
    .B(_08978_),
    .C(_08983_),
    .X(_08984_));
 sky130_fd_sc_hd__or2_1 _15889_ (.A(_08939_),
    .B(_08945_),
    .X(_08985_));
 sky130_fd_sc_hd__nand2_1 _15890_ (.A(_08946_),
    .B(_08985_),
    .Y(_08986_));
 sky130_fd_sc_hd__a21oi_1 _15891_ (.A1(_08982_),
    .A2(_08984_),
    .B1(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__and4_1 _15892_ (.A(_08914_),
    .B(_08948_),
    .C(_08953_),
    .D(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__xor2_1 _15893_ (.A(_08952_),
    .B(_08988_),
    .X(_08989_));
 sky130_fd_sc_hd__o21ai_1 _15894_ (.A1(_08869_),
    .A2(_08978_),
    .B1(_08983_),
    .Y(_08990_));
 sky130_fd_sc_hd__or2_1 _15895_ (.A(_08976_),
    .B(_08979_),
    .X(_08991_));
 sky130_fd_sc_hd__nand2_1 _15896_ (.A(_08980_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__and2b_1 _15897_ (.A_N(_08974_),
    .B(_08973_),
    .X(_08993_));
 sky130_fd_sc_hd__xnor2_1 _15898_ (.A(_08961_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__xnor2_1 _15899_ (.A(_08966_),
    .B(_08971_),
    .Y(_08995_));
 sky130_fd_sc_hd__nor2_1 _15900_ (.A(_08675_),
    .B(_08965_),
    .Y(_08996_));
 sky130_fd_sc_hd__nor2_1 _15901_ (.A(_08616_),
    .B(_08383_),
    .Y(_08997_));
 sky130_fd_sc_hd__xnor2_1 _15902_ (.A(_08968_),
    .B(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__nand2_1 _15903_ (.A(_08996_),
    .B(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__o31a_1 _15904_ (.A1(_08616_),
    .A2(_08383_),
    .A3(_08968_),
    .B1(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__xor2_1 _15905_ (.A(_08995_),
    .B(_09000_),
    .X(_09001_));
 sky130_fd_sc_hd__clkbuf_4 _15906_ (.A(_08318_),
    .X(_09002_));
 sky130_fd_sc_hd__or2_1 _15907_ (.A(_08413_),
    .B(_08742_),
    .X(_09003_));
 sky130_fd_sc_hd__or3_1 _15908_ (.A(_09002_),
    .B(_08675_),
    .C(_09003_),
    .X(_09004_));
 sky130_fd_sc_hd__o22ai_1 _15909_ (.A1(_08977_),
    .A2(_08675_),
    .B1(_08742_),
    .B2(_09002_),
    .Y(_09005_));
 sky130_fd_sc_hd__and2_1 _15910_ (.A(_09004_),
    .B(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__nand2_1 _15911_ (.A(_09001_),
    .B(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__o21a_1 _15912_ (.A1(_08995_),
    .A2(_09000_),
    .B1(_09007_),
    .X(_09008_));
 sky130_fd_sc_hd__or2_1 _15913_ (.A(_08994_),
    .B(_09008_),
    .X(_09009_));
 sky130_fd_sc_hd__nor2_1 _15914_ (.A(_08616_),
    .B(_08374_),
    .Y(_09010_));
 sky130_fd_sc_hd__nor2_1 _15915_ (.A(_08560_),
    .B(_08383_),
    .Y(_09011_));
 sky130_fd_sc_hd__xor2_1 _15916_ (.A(_09010_),
    .B(_09011_),
    .X(_09012_));
 sky130_fd_sc_hd__o21ba_1 _15917_ (.A1(_08742_),
    .A2(_08965_),
    .B1_N(_09012_),
    .X(_09013_));
 sky130_fd_sc_hd__and3b_1 _15918_ (.A_N(_08742_),
    .B(_08782_),
    .C(_09012_),
    .X(_09014_));
 sky130_fd_sc_hd__or4b_1 _15919_ (.A(_08396_),
    .B(_09013_),
    .C(_09014_),
    .D_N(_09011_),
    .X(_09015_));
 sky130_fd_sc_hd__xnor2_1 _15920_ (.A(_08996_),
    .B(_08998_),
    .Y(_09016_));
 sky130_fd_sc_hd__a21oi_1 _15921_ (.A1(_09010_),
    .A2(_09011_),
    .B1(_09014_),
    .Y(_09017_));
 sky130_fd_sc_hd__xnor2_1 _15922_ (.A(_09016_),
    .B(_09017_),
    .Y(_09018_));
 sky130_fd_sc_hd__or2_1 _15923_ (.A(_09003_),
    .B(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__nand2_1 _15924_ (.A(_09003_),
    .B(_09018_),
    .Y(_09020_));
 sky130_fd_sc_hd__nand2_1 _15925_ (.A(_09019_),
    .B(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__or2_1 _15926_ (.A(_09001_),
    .B(_09006_),
    .X(_09022_));
 sky130_fd_sc_hd__and2_1 _15927_ (.A(_09007_),
    .B(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__o21ai_1 _15928_ (.A1(_09016_),
    .A2(_09017_),
    .B1(_09019_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand2_1 _15929_ (.A(_09023_),
    .B(_09024_),
    .Y(_09025_));
 sky130_fd_sc_hd__o31a_1 _15930_ (.A1(_08550_),
    .A2(_09015_),
    .A3(_09021_),
    .B1(_09025_),
    .X(_09026_));
 sky130_fd_sc_hd__xnor2_1 _15931_ (.A(_08994_),
    .B(_09008_),
    .Y(_09027_));
 sky130_fd_sc_hd__or2_1 _15932_ (.A(_09004_),
    .B(_09027_),
    .X(_09028_));
 sky130_fd_sc_hd__nand2_1 _15933_ (.A(_09004_),
    .B(_09027_),
    .Y(_09029_));
 sky130_fd_sc_hd__o211ai_1 _15934_ (.A1(_09023_),
    .A2(_09024_),
    .B1(_09028_),
    .C1(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__a21o_1 _15935_ (.A1(_09009_),
    .A2(_09028_),
    .B1(_08992_),
    .X(_09031_));
 sky130_fd_sc_hd__o21a_1 _15936_ (.A1(_09026_),
    .A2(_09030_),
    .B1(_09031_),
    .X(_09032_));
 sky130_fd_sc_hd__a21oi_1 _15937_ (.A1(_08992_),
    .A2(_09009_),
    .B1(_09032_),
    .Y(_09033_));
 sky130_fd_sc_hd__and4_1 _15938_ (.A(_08948_),
    .B(_08984_),
    .C(_08990_),
    .D(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__or2b_1 _15939_ (.A(_08953_),
    .B_N(_08946_),
    .X(_09035_));
 sky130_fd_sc_hd__xor2_1 _15940_ (.A(_08986_),
    .B(_08982_),
    .X(_09036_));
 sky130_fd_sc_hd__and4_1 _15941_ (.A(_08914_),
    .B(_09034_),
    .C(_09035_),
    .D(_09036_),
    .X(_09037_));
 sky130_fd_sc_hd__and2_1 _15942_ (.A(_08952_),
    .B(_08988_),
    .X(_09038_));
 sky130_fd_sc_hd__a21o_1 _15943_ (.A1(_08989_),
    .A2(_09037_),
    .B1(_09038_),
    .X(_09039_));
 sky130_fd_sc_hd__nor2_1 _15944_ (.A(_08910_),
    .B(_08951_),
    .Y(_09040_));
 sky130_fd_sc_hd__xnor2_1 _15945_ (.A(_08911_),
    .B(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__a22o_2 _15946_ (.A1(_08911_),
    .A2(_08951_),
    .B1(_09039_),
    .B2(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__nor2_1 _15947_ (.A(_08849_),
    .B(_08912_),
    .Y(_09043_));
 sky130_fd_sc_hd__xnor2_2 _15948_ (.A(_08853_),
    .B(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__a22o_2 _15949_ (.A1(_08853_),
    .A2(_08912_),
    .B1(_09042_),
    .B2(_09044_),
    .X(_09045_));
 sky130_fd_sc_hd__nor2_1 _15950_ (.A(_08850_),
    .B(_08852_),
    .Y(_09046_));
 sky130_fd_sc_hd__inv_2 _15951_ (.A(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_1 _15952_ (.A(_09047_),
    .B(_08854_),
    .Y(_09048_));
 sky130_fd_sc_hd__xnor2_2 _15953_ (.A(_08760_),
    .B(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__a2bb2o_2 _15954_ (.A1_N(_08760_),
    .A2_N(_08854_),
    .B1(_09045_),
    .B2(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__or2_1 _15955_ (.A(_08640_),
    .B(_08691_),
    .X(_09051_));
 sky130_fd_sc_hd__nand2_1 _15956_ (.A(_08692_),
    .B(_08697_),
    .Y(_09052_));
 sky130_fd_sc_hd__nand2_1 _15957_ (.A(_08494_),
    .B(_08497_),
    .Y(_09053_));
 sky130_fd_sc_hd__nand2_1 _15958_ (.A(_08306_),
    .B(_08329_),
    .Y(_09054_));
 sky130_fd_sc_hd__o31a_1 _15959_ (.A1(_08344_),
    .A2(_08330_),
    .A3(_08351_),
    .B1(_09054_),
    .X(_09055_));
 sky130_fd_sc_hd__or4_1 _15960_ (.A(_08423_),
    .B(_08452_),
    .C(_08465_),
    .D(_08350_),
    .X(_09056_));
 sky130_fd_sc_hd__o22ai_1 _15961_ (.A1(_08424_),
    .A2(_08465_),
    .B1(_08351_),
    .B2(_08452_),
    .Y(_09057_));
 sky130_fd_sc_hd__nand2_1 _15962_ (.A(_09056_),
    .B(_09057_),
    .Y(_09058_));
 sky130_fd_sc_hd__or2_1 _15963_ (.A(_08486_),
    .B(_08485_),
    .X(_09059_));
 sky130_fd_sc_hd__xnor2_1 _15964_ (.A(_09058_),
    .B(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__xnor2_1 _15965_ (.A(_09055_),
    .B(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__xnor2_1 _15966_ (.A(_09053_),
    .B(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__or4_1 _15967_ (.A(_08318_),
    .B(_08290_),
    .C(_08305_),
    .D(_08362_),
    .X(_09063_));
 sky130_fd_sc_hd__buf_2 _15968_ (.A(_08362_),
    .X(_09064_));
 sky130_fd_sc_hd__o22ai_1 _15969_ (.A1(_08318_),
    .A2(_08387_),
    .B1(_09064_),
    .B2(_08290_),
    .Y(_09065_));
 sky130_fd_sc_hd__nand2_1 _15970_ (.A(_09063_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__nor2_1 _15971_ (.A(_08344_),
    .B(_08407_),
    .Y(_09067_));
 sky130_fd_sc_hd__xnor2_1 _15972_ (.A(_09066_),
    .B(_09067_),
    .Y(_09068_));
 sky130_fd_sc_hd__buf_4 _15973_ (.A(_08294_),
    .X(_09069_));
 sky130_fd_sc_hd__a22oi_4 _15974_ (.A1(\rbzero.wall_tracer.stepDistX[2] ),
    .A2(_06100_),
    .B1(_09069_),
    .B2(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_09070_));
 sky130_fd_sc_hd__and2_1 _15975_ (.A(_08395_),
    .B(_09070_),
    .X(_09071_));
 sky130_fd_sc_hd__a21oi_2 _15976_ (.A1(_08269_),
    .A2(_08370_),
    .B1(_09069_),
    .Y(_09072_));
 sky130_fd_sc_hd__inv_2 _15977_ (.A(_08140_),
    .Y(_09073_));
 sky130_fd_sc_hd__nor4_2 _15978_ (.A(_08121_),
    .B(_08126_),
    .C(_08134_),
    .D(_08295_),
    .Y(_09074_));
 sky130_fd_sc_hd__o41a_1 _15979_ (.A1(_08121_),
    .A2(_08126_),
    .A3(_08134_),
    .A4(_08295_),
    .B1(_08140_),
    .X(_09075_));
 sky130_fd_sc_hd__a211o_1 _15980_ (.A1(_09073_),
    .A2(_09074_),
    .B1(_09075_),
    .C1(_08269_),
    .X(_09076_));
 sky130_fd_sc_hd__a22o_2 _15981_ (.A1(\rbzero.wall_tracer.stepDistY[4] ),
    .A2(_09069_),
    .B1(_09072_),
    .B2(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__nand3_1 _15982_ (.A(_08375_),
    .B(_08404_),
    .C(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__nand2_1 _15983_ (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .B(_08354_),
    .Y(_09079_));
 sky130_fd_sc_hd__a21o_1 _15984_ (.A1(_08372_),
    .A2(_09079_),
    .B1(_06100_),
    .X(_09080_));
 sky130_fd_sc_hd__nand2_2 _15985_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_08554_),
    .Y(_09081_));
 sky130_fd_sc_hd__a2bb2o_1 _15986_ (.A1_N(_09080_),
    .A2_N(_09081_),
    .B1(_09077_),
    .B2(_08403_),
    .X(_09082_));
 sky130_fd_sc_hd__or4bb_1 _15987_ (.A(_08366_),
    .B(_09071_),
    .C_N(_09078_),
    .D_N(_09082_),
    .X(_09083_));
 sky130_fd_sc_hd__a2bb2o_1 _15988_ (.A1_N(_08366_),
    .A2_N(_09071_),
    .B1(_09078_),
    .B2(_09082_),
    .X(_09084_));
 sky130_fd_sc_hd__or2_1 _15989_ (.A(_08375_),
    .B(_08384_),
    .X(_09085_));
 sky130_fd_sc_hd__nand2_1 _15990_ (.A(_08375_),
    .B(_08384_),
    .Y(_09086_));
 sky130_fd_sc_hd__a21bo_1 _15991_ (.A1(_08367_),
    .A2(_09085_),
    .B1_N(_09086_),
    .X(_09087_));
 sky130_fd_sc_hd__nand3_2 _15992_ (.A(_09083_),
    .B(_09084_),
    .C(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__a21o_1 _15993_ (.A1(_09083_),
    .A2(_09084_),
    .B1(_09087_),
    .X(_09089_));
 sky130_fd_sc_hd__nand3_1 _15994_ (.A(_09068_),
    .B(_09088_),
    .C(_09089_),
    .Y(_09090_));
 sky130_fd_sc_hd__a21o_1 _15995_ (.A1(_09088_),
    .A2(_09089_),
    .B1(_09068_),
    .X(_09091_));
 sky130_fd_sc_hd__and2b_1 _15996_ (.A_N(_08398_),
    .B(_08386_),
    .X(_09092_));
 sky130_fd_sc_hd__a21o_1 _15997_ (.A1(_08353_),
    .A2(_08399_),
    .B1(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__nand3_1 _15998_ (.A(_09090_),
    .B(_09091_),
    .C(_09093_),
    .Y(_09094_));
 sky130_fd_sc_hd__a21o_1 _15999_ (.A1(_09090_),
    .A2(_09091_),
    .B1(_09093_),
    .X(_09095_));
 sky130_fd_sc_hd__and3_1 _16000_ (.A(_09062_),
    .B(_09094_),
    .C(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__a21oi_1 _16001_ (.A1(_09094_),
    .A2(_09095_),
    .B1(_09062_),
    .Y(_09097_));
 sky130_fd_sc_hd__or2_1 _16002_ (.A(_09096_),
    .B(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__a21oi_1 _16003_ (.A1(_08431_),
    .A2(_08501_),
    .B1(_08429_),
    .Y(_09099_));
 sky130_fd_sc_hd__nor2_1 _16004_ (.A(_09098_),
    .B(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__and2_1 _16005_ (.A(_09098_),
    .B(_09099_),
    .X(_09101_));
 sky130_fd_sc_hd__nor2_1 _16006_ (.A(_09100_),
    .B(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__o21ai_1 _16007_ (.A1(_08630_),
    .A2(_08631_),
    .B1(_08633_),
    .Y(_09103_));
 sky130_fd_sc_hd__or2_1 _16008_ (.A(_08493_),
    .B(_08499_),
    .X(_09104_));
 sky130_fd_sc_hd__or2b_1 _16009_ (.A(_08500_),
    .B_N(_08491_),
    .X(_09105_));
 sky130_fd_sc_hd__nand2_2 _16010_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08319_),
    .Y(_09106_));
 sky130_fd_sc_hd__nor2_1 _16011_ (.A(_09106_),
    .B(_08616_),
    .Y(_09107_));
 sky130_fd_sc_hd__nor2_1 _16012_ (.A(_08544_),
    .B(_08967_),
    .Y(_09108_));
 sky130_fd_sc_hd__xnor2_1 _16013_ (.A(_09107_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__or3_1 _16014_ (.A(_08561_),
    .B(_08620_),
    .C(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__o21ai_1 _16015_ (.A1(_08561_),
    .A2(_08620_),
    .B1(_09109_),
    .Y(_09111_));
 sky130_fd_sc_hd__and2_1 _16016_ (.A(_09110_),
    .B(_09111_),
    .X(_09112_));
 sky130_fd_sc_hd__nor2_1 _16017_ (.A(_08473_),
    .B(_08580_),
    .Y(_09113_));
 sky130_fd_sc_hd__nor2_1 _16018_ (.A(_08444_),
    .B(_08587_),
    .Y(_09114_));
 sky130_fd_sc_hd__xnor2_1 _16019_ (.A(_09113_),
    .B(_09114_),
    .Y(_09115_));
 sky130_fd_sc_hd__or2_1 _16020_ (.A(_08528_),
    .B(_08601_),
    .X(_09116_));
 sky130_fd_sc_hd__xnor2_1 _16021_ (.A(_09115_),
    .B(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__and2_1 _16022_ (.A(_08627_),
    .B(_08628_),
    .X(_09118_));
 sky130_fd_sc_hd__nor2_1 _16023_ (.A(_09117_),
    .B(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__and2_1 _16024_ (.A(_09117_),
    .B(_09118_),
    .X(_09120_));
 sky130_fd_sc_hd__nor2_1 _16025_ (.A(_09119_),
    .B(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__xnor2_1 _16026_ (.A(_09112_),
    .B(_09121_),
    .Y(_09122_));
 sky130_fd_sc_hd__a21o_1 _16027_ (.A1(_09104_),
    .A2(_09105_),
    .B1(_09122_),
    .X(_09123_));
 sky130_fd_sc_hd__nand3_1 _16028_ (.A(_09104_),
    .B(_09105_),
    .C(_09122_),
    .Y(_09124_));
 sky130_fd_sc_hd__nand2_1 _16029_ (.A(_09123_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__xnor2_1 _16030_ (.A(_09103_),
    .B(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__xnor2_1 _16031_ (.A(_09102_),
    .B(_09126_),
    .Y(_09127_));
 sky130_fd_sc_hd__nor2_1 _16032_ (.A(_08502_),
    .B(_08541_),
    .Y(_09128_));
 sky130_fd_sc_hd__a21oi_1 _16033_ (.A1(_08542_),
    .A2(_08639_),
    .B1(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__xor2_1 _16034_ (.A(_09127_),
    .B(_09129_),
    .X(_09130_));
 sky130_fd_sc_hd__or2b_1 _16035_ (.A(_08638_),
    .B_N(_08614_),
    .X(_09131_));
 sky130_fd_sc_hd__nand2_4 _16036_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08543_),
    .Y(_09132_));
 sky130_fd_sc_hd__buf_2 _16037_ (.A(_09132_),
    .X(_09133_));
 sky130_fd_sc_hd__or2_1 _16038_ (.A(_08550_),
    .B(_09133_),
    .X(_09134_));
 sky130_fd_sc_hd__clkbuf_4 _16039_ (.A(_08616_),
    .X(_09135_));
 sky130_fd_sc_hd__o31a_1 _16040_ (.A1(_08545_),
    .A2(_08557_),
    .A3(_09135_),
    .B1(_08622_),
    .X(_09136_));
 sky130_fd_sc_hd__nor2_1 _16041_ (.A(_09134_),
    .B(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__and2_1 _16042_ (.A(_09134_),
    .B(_09136_),
    .X(_09138_));
 sky130_fd_sc_hd__or2_1 _16043_ (.A(_09137_),
    .B(_09138_),
    .X(_09139_));
 sky130_fd_sc_hd__a21oi_2 _16044_ (.A1(_08636_),
    .A2(_09131_),
    .B1(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__and3_1 _16045_ (.A(_08636_),
    .B(_09131_),
    .C(_09139_),
    .X(_09141_));
 sky130_fd_sc_hd__nor2_1 _16046_ (.A(_09140_),
    .B(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__xnor2_1 _16047_ (.A(_09130_),
    .B(_09142_),
    .Y(_09143_));
 sky130_fd_sc_hd__a21o_1 _16048_ (.A1(_09051_),
    .A2(_09052_),
    .B1(_09143_),
    .X(_09144_));
 sky130_fd_sc_hd__nand3_1 _16049_ (.A(_09143_),
    .B(_09051_),
    .C(_09052_),
    .Y(_09145_));
 sky130_fd_sc_hd__and2_1 _16050_ (.A(_09144_),
    .B(_09145_),
    .X(_09146_));
 sky130_fd_sc_hd__xnor2_2 _16051_ (.A(_08695_),
    .B(_09146_),
    .Y(_09147_));
 sky130_fd_sc_hd__nor2_1 _16052_ (.A(_09047_),
    .B(_08760_),
    .Y(_09148_));
 sky130_fd_sc_hd__or2_1 _16053_ (.A(_08758_),
    .B(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__xnor2_2 _16054_ (.A(_09147_),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__and2b_1 _16055_ (.A_N(_09147_),
    .B(_09148_),
    .X(_09151_));
 sky130_fd_sc_hd__a21o_2 _16056_ (.A1(_09050_),
    .A2(_09150_),
    .B1(_09151_),
    .X(_09152_));
 sky130_fd_sc_hd__a21o_1 _16057_ (.A1(_09112_),
    .A2(_09121_),
    .B1(_09119_),
    .X(_09153_));
 sky130_fd_sc_hd__or2_1 _16058_ (.A(_09055_),
    .B(_09060_),
    .X(_09154_));
 sky130_fd_sc_hd__or2b_1 _16059_ (.A(_09061_),
    .B_N(_09053_),
    .X(_09155_));
 sky130_fd_sc_hd__or4_2 _16060_ (.A(_06461_),
    .B(_09106_),
    .C(_08922_),
    .D(_08967_),
    .X(_09156_));
 sky130_fd_sc_hd__buf_2 _16061_ (.A(_08967_),
    .X(_09157_));
 sky130_fd_sc_hd__buf_2 _16062_ (.A(_09106_),
    .X(_09158_));
 sky130_fd_sc_hd__o22ai_1 _16063_ (.A1(_08544_),
    .A2(_08922_),
    .B1(_09157_),
    .B2(_09158_),
    .Y(_09159_));
 sky130_fd_sc_hd__nand2_1 _16064_ (.A(_09156_),
    .B(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__or3_1 _16065_ (.A(_08616_),
    .B(_08620_),
    .C(_09160_),
    .X(_09161_));
 sky130_fd_sc_hd__clkbuf_4 _16066_ (.A(_08620_),
    .X(_09162_));
 sky130_fd_sc_hd__o21ai_1 _16067_ (.A1(_09135_),
    .A2(_09162_),
    .B1(_09160_),
    .Y(_09163_));
 sky130_fd_sc_hd__and2_1 _16068_ (.A(_09161_),
    .B(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__nor2_1 _16069_ (.A(_08486_),
    .B(_08580_),
    .Y(_09165_));
 sky130_fd_sc_hd__o22a_1 _16070_ (.A1(_08486_),
    .A2(_08587_),
    .B1(_08580_),
    .B2(_08444_),
    .X(_09166_));
 sky130_fd_sc_hd__a21o_1 _16071_ (.A1(_09114_),
    .A2(_09165_),
    .B1(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__or2_1 _16072_ (.A(_08473_),
    .B(_08601_),
    .X(_09168_));
 sky130_fd_sc_hd__xnor2_1 _16073_ (.A(_09167_),
    .B(_09168_),
    .Y(_09169_));
 sky130_fd_sc_hd__nand2_1 _16074_ (.A(_09113_),
    .B(_09114_),
    .Y(_09170_));
 sky130_fd_sc_hd__o31a_1 _16075_ (.A1(_08528_),
    .A2(_08602_),
    .A3(_09115_),
    .B1(_09170_),
    .X(_09171_));
 sky130_fd_sc_hd__nor2_1 _16076_ (.A(_09169_),
    .B(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__and2_1 _16077_ (.A(_09169_),
    .B(_09171_),
    .X(_09173_));
 sky130_fd_sc_hd__nor2_1 _16078_ (.A(_09172_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__xnor2_1 _16079_ (.A(_09164_),
    .B(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__a21o_1 _16080_ (.A1(_09154_),
    .A2(_09155_),
    .B1(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__nand3_1 _16081_ (.A(_09154_),
    .B(_09155_),
    .C(_09175_),
    .Y(_09177_));
 sky130_fd_sc_hd__nand2_1 _16082_ (.A(_09176_),
    .B(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__xnor2_1 _16083_ (.A(_09153_),
    .B(_09178_),
    .Y(_09179_));
 sky130_fd_sc_hd__o21ai_2 _16084_ (.A1(_09058_),
    .A2(_09059_),
    .B1(_09056_),
    .Y(_09180_));
 sky130_fd_sc_hd__o31a_1 _16085_ (.A1(_08492_),
    .A2(_08407_),
    .A3(_09066_),
    .B1(_09063_),
    .X(_09181_));
 sky130_fd_sc_hd__or2_1 _16086_ (.A(_08465_),
    .B(_08328_),
    .X(_09182_));
 sky130_fd_sc_hd__or3_1 _16087_ (.A(_08495_),
    .B(_08351_),
    .C(_09182_),
    .X(_09183_));
 sky130_fd_sc_hd__o22ai_1 _16088_ (.A1(_08495_),
    .A2(_08407_),
    .B1(_08351_),
    .B2(_08487_),
    .Y(_09184_));
 sky130_fd_sc_hd__nand2_1 _16089_ (.A(_09183_),
    .B(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__nor2_1 _16090_ (.A(_08424_),
    .B(_08533_),
    .Y(_09186_));
 sky130_fd_sc_hd__xor2_1 _16091_ (.A(_09185_),
    .B(_09186_),
    .X(_09187_));
 sky130_fd_sc_hd__xnor2_1 _16092_ (.A(_09181_),
    .B(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__xnor2_2 _16093_ (.A(_09180_),
    .B(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__or2_1 _16094_ (.A(_08317_),
    .B(_08362_),
    .X(_09190_));
 sky130_fd_sc_hd__or3_1 _16095_ (.A(_08290_),
    .B(_09190_),
    .C(_09071_),
    .X(_09191_));
 sky130_fd_sc_hd__buf_2 _16096_ (.A(_09071_),
    .X(_09192_));
 sky130_fd_sc_hd__o21ai_1 _16097_ (.A1(_08413_),
    .A2(_09192_),
    .B1(_09190_),
    .Y(_09193_));
 sky130_fd_sc_hd__nand2_1 _16098_ (.A(_09191_),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__nor2_1 _16099_ (.A(_08492_),
    .B(_08387_),
    .Y(_09195_));
 sky130_fd_sc_hd__xnor2_1 _16100_ (.A(_09194_),
    .B(_09195_),
    .Y(_09196_));
 sky130_fd_sc_hd__a21boi_2 _16101_ (.A1(\rbzero.wall_tracer.stepDistX[3] ),
    .A2(_06101_),
    .B1_N(_09080_),
    .Y(_09197_));
 sky130_fd_sc_hd__clkbuf_4 _16102_ (.A(_09197_),
    .X(_09198_));
 sky130_fd_sc_hd__nor2_1 _16103_ (.A(_08965_),
    .B(_09198_),
    .Y(_09199_));
 sky130_fd_sc_hd__nand2_1 _16104_ (.A(_08404_),
    .B(_09077_),
    .Y(_09200_));
 sky130_fd_sc_hd__or3_1 _16105_ (.A(_08140_),
    .B(_08142_),
    .C(_08368_),
    .X(_09201_));
 sky130_fd_sc_hd__o21ai_1 _16106_ (.A1(_08140_),
    .A2(_08368_),
    .B1(_08142_),
    .Y(_09202_));
 sky130_fd_sc_hd__a31o_1 _16107_ (.A1(_08355_),
    .A2(_09201_),
    .A3(_09202_),
    .B1(_08371_),
    .X(_09203_));
 sky130_fd_sc_hd__or3b_4 _16108_ (.A(_08390_),
    .B(_09203_),
    .C_N(_08164_),
    .X(_09204_));
 sky130_fd_sc_hd__xor2_2 _16109_ (.A(_09200_),
    .B(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__xnor2_2 _16110_ (.A(_09199_),
    .B(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__nand2_1 _16111_ (.A(_09078_),
    .B(_09083_),
    .Y(_09207_));
 sky130_fd_sc_hd__xnor2_2 _16112_ (.A(_09206_),
    .B(_09207_),
    .Y(_09208_));
 sky130_fd_sc_hd__xnor2_2 _16113_ (.A(_09196_),
    .B(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__and2_1 _16114_ (.A(_09088_),
    .B(_09090_),
    .X(_09210_));
 sky130_fd_sc_hd__xor2_2 _16115_ (.A(_09209_),
    .B(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__xor2_2 _16116_ (.A(_09189_),
    .B(_09211_),
    .X(_09212_));
 sky130_fd_sc_hd__a21boi_2 _16117_ (.A1(_09062_),
    .A2(_09095_),
    .B1_N(_09094_),
    .Y(_09213_));
 sky130_fd_sc_hd__xnor2_1 _16118_ (.A(_09212_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__xnor2_1 _16119_ (.A(_09179_),
    .B(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__a21oi_1 _16120_ (.A1(_09102_),
    .A2(_09126_),
    .B1(_09100_),
    .Y(_09216_));
 sky130_fd_sc_hd__nor2_1 _16121_ (.A(_09215_),
    .B(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__nand2_1 _16122_ (.A(_09215_),
    .B(_09216_),
    .Y(_09218_));
 sky130_fd_sc_hd__and2b_1 _16123_ (.A_N(_09217_),
    .B(_09218_),
    .X(_09219_));
 sky130_fd_sc_hd__or2b_1 _16124_ (.A(_09125_),
    .B_N(_09103_),
    .X(_09220_));
 sky130_fd_sc_hd__nand2_1 _16125_ (.A(_09107_),
    .B(_09108_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand2_4 _16126_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08319_),
    .Y(_09222_));
 sky130_fd_sc_hd__or2_1 _16127_ (.A(_08560_),
    .B(_09222_),
    .X(_09223_));
 sky130_fd_sc_hd__nor2_1 _16128_ (.A(_09134_),
    .B(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__clkbuf_4 _16129_ (.A(_09222_),
    .X(_09225_));
 sky130_fd_sc_hd__o22a_1 _16130_ (.A1(_08561_),
    .A2(_09133_),
    .B1(_09225_),
    .B2(_08550_),
    .X(_09226_));
 sky130_fd_sc_hd__or2_1 _16131_ (.A(_09224_),
    .B(_09226_),
    .X(_09227_));
 sky130_fd_sc_hd__a21oi_1 _16132_ (.A1(_09221_),
    .A2(_09110_),
    .B1(_09227_),
    .Y(_09228_));
 sky130_fd_sc_hd__and3_1 _16133_ (.A(_09221_),
    .B(_09110_),
    .C(_09227_),
    .X(_09229_));
 sky130_fd_sc_hd__nor2_1 _16134_ (.A(_09228_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__nand2_1 _16135_ (.A(_09137_),
    .B(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__or2_1 _16136_ (.A(_09137_),
    .B(_09230_),
    .X(_09232_));
 sky130_fd_sc_hd__nand2_1 _16137_ (.A(_09231_),
    .B(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__a21oi_4 _16138_ (.A1(_09123_),
    .A2(_09220_),
    .B1(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__and3_1 _16139_ (.A(_09123_),
    .B(_09220_),
    .C(_09233_),
    .X(_09235_));
 sky130_fd_sc_hd__nor2_1 _16140_ (.A(_09234_),
    .B(_09235_),
    .Y(_09236_));
 sky130_fd_sc_hd__xnor2_2 _16141_ (.A(_09219_),
    .B(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__or2_1 _16142_ (.A(_09127_),
    .B(_09129_),
    .X(_09238_));
 sky130_fd_sc_hd__nand2_1 _16143_ (.A(_09130_),
    .B(_09142_),
    .Y(_09239_));
 sky130_fd_sc_hd__nand2_1 _16144_ (.A(_09238_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__xnor2_2 _16145_ (.A(_09237_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__xnor2_1 _16146_ (.A(_09140_),
    .B(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__a21boi_1 _16147_ (.A1(_08695_),
    .A2(_09146_),
    .B1_N(_09144_),
    .Y(_09243_));
 sky130_fd_sc_hd__xor2_1 _16148_ (.A(_09242_),
    .B(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__and2b_1 _16149_ (.A_N(_09147_),
    .B(_08758_),
    .X(_09245_));
 sky130_fd_sc_hd__nand2_1 _16150_ (.A(_09244_),
    .B(_09245_),
    .Y(_09246_));
 sky130_fd_sc_hd__or2_1 _16151_ (.A(_09244_),
    .B(_09245_),
    .X(_09247_));
 sky130_fd_sc_hd__and2_2 _16152_ (.A(_09246_),
    .B(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__xor2_4 _16153_ (.A(_09152_),
    .B(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__and2b_1 _16154_ (.A_N(_08272_),
    .B(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__and2b_1 _16155_ (.A_N(_09249_),
    .B(_08272_),
    .X(_09251_));
 sky130_fd_sc_hd__nor2_1 _16156_ (.A(_09250_),
    .B(_09251_),
    .Y(_09252_));
 sky130_fd_sc_hd__xor2_4 _16157_ (.A(_09050_),
    .B(_09150_),
    .X(_09253_));
 sky130_fd_sc_hd__mux2_1 _16158_ (.A0(\rbzero.debug_overlay.playerY[-7] ),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_04618_),
    .X(_09254_));
 sky130_fd_sc_hd__or2_1 _16159_ (.A(_09253_),
    .B(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__mux2_1 _16160_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_04618_),
    .X(_09256_));
 sky130_fd_sc_hd__xor2_4 _16161_ (.A(_09045_),
    .B(_09049_),
    .X(_09257_));
 sky130_fd_sc_hd__xor2_4 _16162_ (.A(_09042_),
    .B(_09044_),
    .X(_09258_));
 sky130_fd_sc_hd__mux2_1 _16163_ (.A0(\rbzero.debug_overlay.playerY[-9] ),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_04618_),
    .X(_09259_));
 sky130_fd_sc_hd__o211a_1 _16164_ (.A1(_09256_),
    .A2(_09257_),
    .B1(_09258_),
    .C1(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__a21o_1 _16165_ (.A1(_09256_),
    .A2(_09257_),
    .B1(_09260_),
    .X(_09261_));
 sky130_fd_sc_hd__and2_1 _16166_ (.A(_09253_),
    .B(_09254_),
    .X(_09262_));
 sky130_fd_sc_hd__a21o_1 _16167_ (.A1(_09255_),
    .A2(_09261_),
    .B1(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__xnor2_1 _16168_ (.A(_09252_),
    .B(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__clkbuf_4 _16169_ (.A(_08334_),
    .X(_09265_));
 sky130_fd_sc_hd__buf_2 _16170_ (.A(_09265_),
    .X(_09266_));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(_09266_),
    .A1(_06377_),
    .S(_08263_),
    .X(_09267_));
 sky130_fd_sc_hd__clkbuf_4 _16172_ (.A(_09267_),
    .X(_09268_));
 sky130_fd_sc_hd__o21ai_1 _16173_ (.A1(_09264_),
    .A2(_09268_),
    .B1(_08270_),
    .Y(_09269_));
 sky130_fd_sc_hd__a21o_1 _16174_ (.A1(_09264_),
    .A2(_09268_),
    .B1(_09269_),
    .X(_09270_));
 sky130_fd_sc_hd__o211a_1 _16175_ (.A1(\rbzero.texu_hot[0] ),
    .A2(_08270_),
    .B1(_09270_),
    .C1(_08211_),
    .X(_00466_));
 sky130_fd_sc_hd__a21boi_2 _16176_ (.A1(_09152_),
    .A2(_09248_),
    .B1_N(_09246_),
    .Y(_09271_));
 sky130_fd_sc_hd__or2_2 _16177_ (.A(_09242_),
    .B(_09243_),
    .X(_09272_));
 sky130_fd_sc_hd__or2b_1 _16178_ (.A(_09178_),
    .B_N(_09153_),
    .X(_09273_));
 sky130_fd_sc_hd__nor2_1 _16179_ (.A(_08616_),
    .B(_09132_),
    .Y(_09274_));
 sky130_fd_sc_hd__xnor2_1 _16180_ (.A(_09223_),
    .B(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__nand2_4 _16181_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08543_),
    .Y(_09276_));
 sky130_fd_sc_hd__nor2_1 _16182_ (.A(_08549_),
    .B(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__xnor2_1 _16183_ (.A(_09275_),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__and3_1 _16184_ (.A(_09156_),
    .B(_09161_),
    .C(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__a21oi_2 _16185_ (.A1(_09156_),
    .A2(_09161_),
    .B1(_09278_),
    .Y(_09280_));
 sky130_fd_sc_hd__nor4_1 _16186_ (.A(_09224_),
    .B(_09228_),
    .C(_09279_),
    .D(_09280_),
    .Y(_09281_));
 sky130_fd_sc_hd__o22a_1 _16187_ (.A1(_09224_),
    .A2(_09228_),
    .B1(_09279_),
    .B2(_09280_),
    .X(_09282_));
 sky130_fd_sc_hd__nor2_1 _16188_ (.A(_09281_),
    .B(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__a21oi_1 _16189_ (.A1(_09176_),
    .A2(_09273_),
    .B1(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__and3_1 _16190_ (.A(_09176_),
    .B(_09273_),
    .C(_09283_),
    .X(_09285_));
 sky130_fd_sc_hd__nor2_1 _16191_ (.A(_09284_),
    .B(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__xnor2_1 _16192_ (.A(_09231_),
    .B(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__a21o_1 _16193_ (.A1(_09164_),
    .A2(_09174_),
    .B1(_09172_),
    .X(_09288_));
 sky130_fd_sc_hd__or2_1 _16194_ (.A(_09181_),
    .B(_09187_),
    .X(_09289_));
 sky130_fd_sc_hd__or2b_1 _16195_ (.A(_09188_),
    .B_N(_09180_),
    .X(_09290_));
 sky130_fd_sc_hd__nor4_1 _16196_ (.A(_06461_),
    .B(_09158_),
    .C(_08888_),
    .D(_08922_),
    .Y(_09291_));
 sky130_fd_sc_hd__o22a_1 _16197_ (.A1(_08544_),
    .A2(_08888_),
    .B1(_08922_),
    .B2(_09158_),
    .X(_09292_));
 sky130_fd_sc_hd__nor2_1 _16198_ (.A(_09291_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__nor2_1 _16199_ (.A(_09157_),
    .B(_08619_),
    .Y(_09294_));
 sky130_fd_sc_hd__xor2_1 _16200_ (.A(_09293_),
    .B(_09294_),
    .X(_09295_));
 sky130_fd_sc_hd__nor2_1 _16201_ (.A(_08424_),
    .B(_08587_),
    .Y(_09296_));
 sky130_fd_sc_hd__xnor2_1 _16202_ (.A(_09165_),
    .B(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__or2_1 _16203_ (.A(_08444_),
    .B(_08602_),
    .X(_09298_));
 sky130_fd_sc_hd__xnor2_1 _16204_ (.A(_09297_),
    .B(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__nand2_1 _16205_ (.A(_09114_),
    .B(_09165_),
    .Y(_09300_));
 sky130_fd_sc_hd__o31a_1 _16206_ (.A1(_08473_),
    .A2(_08602_),
    .A3(_09166_),
    .B1(_09300_),
    .X(_09301_));
 sky130_fd_sc_hd__nor2_1 _16207_ (.A(_09299_),
    .B(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__and2_1 _16208_ (.A(_09299_),
    .B(_09301_),
    .X(_09303_));
 sky130_fd_sc_hd__nor2_1 _16209_ (.A(_09302_),
    .B(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__xnor2_1 _16210_ (.A(_09295_),
    .B(_09304_),
    .Y(_09305_));
 sky130_fd_sc_hd__a21o_1 _16211_ (.A1(_09289_),
    .A2(_09290_),
    .B1(_09305_),
    .X(_09306_));
 sky130_fd_sc_hd__nand3_1 _16212_ (.A(_09289_),
    .B(_09290_),
    .C(_09305_),
    .Y(_09307_));
 sky130_fd_sc_hd__nand2_1 _16213_ (.A(_09306_),
    .B(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__xnor2_1 _16214_ (.A(_09288_),
    .B(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__a21bo_1 _16215_ (.A1(_09184_),
    .A2(_09186_),
    .B1_N(_09183_),
    .X(_09310_));
 sky130_fd_sc_hd__o31ai_2 _16216_ (.A1(_08492_),
    .A2(_08387_),
    .A3(_09194_),
    .B1(_09191_),
    .Y(_09311_));
 sky130_fd_sc_hd__nor2_2 _16217_ (.A(_08452_),
    .B(_08387_),
    .Y(_09312_));
 sky130_fd_sc_hd__xnor2_1 _16218_ (.A(_09182_),
    .B(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__nor2_1 _16219_ (.A(_08485_),
    .B(_08351_),
    .Y(_09314_));
 sky130_fd_sc_hd__xor2_1 _16220_ (.A(_09313_),
    .B(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__xnor2_1 _16221_ (.A(_09311_),
    .B(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__xnor2_2 _16222_ (.A(_09310_),
    .B(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__nor2_1 _16223_ (.A(_08344_),
    .B(_09064_),
    .Y(_09318_));
 sky130_fd_sc_hd__nor2_1 _16224_ (.A(_08977_),
    .B(_09192_),
    .Y(_09319_));
 sky130_fd_sc_hd__nor2_2 _16225_ (.A(_08318_),
    .B(_09197_),
    .Y(_09320_));
 sky130_fd_sc_hd__o22a_1 _16226_ (.A1(_09002_),
    .A2(_09192_),
    .B1(_09197_),
    .B2(_08413_),
    .X(_09321_));
 sky130_fd_sc_hd__a21oi_2 _16227_ (.A1(_09319_),
    .A2(_09320_),
    .B1(_09321_),
    .Y(_09322_));
 sky130_fd_sc_hd__xor2_2 _16228_ (.A(_09318_),
    .B(_09322_),
    .X(_09323_));
 sky130_fd_sc_hd__and2_1 _16229_ (.A(\rbzero.wall_tracer.stepDistX[4] ),
    .B(_06100_),
    .X(_09324_));
 sky130_fd_sc_hd__a21oi_2 _16230_ (.A1(_08292_),
    .A2(_09077_),
    .B1(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__clkbuf_4 _16231_ (.A(_09325_),
    .X(_09326_));
 sky130_fd_sc_hd__nor2_1 _16232_ (.A(_08965_),
    .B(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__o31a_1 _16233_ (.A1(_08140_),
    .A2(_08142_),
    .A3(_08368_),
    .B1(_08145_),
    .X(_09328_));
 sky130_fd_sc_hd__nor2_1 _16234_ (.A(_08142_),
    .B(_08145_),
    .Y(_09329_));
 sky130_fd_sc_hd__a31o_1 _16235_ (.A1(_09073_),
    .A2(_09074_),
    .A3(_09329_),
    .B1(_08269_),
    .X(_09330_));
 sky130_fd_sc_hd__o21ai_4 _16236_ (.A1(_09328_),
    .A2(_09330_),
    .B1(_09072_),
    .Y(_09331_));
 sky130_fd_sc_hd__or3b_1 _16237_ (.A(_08390_),
    .B(_09331_),
    .C_N(_08164_),
    .X(_09332_));
 sky130_fd_sc_hd__or2_1 _16238_ (.A(_08383_),
    .B(_09203_),
    .X(_09333_));
 sky130_fd_sc_hd__or3_2 _16239_ (.A(_08169_),
    .B(_08390_),
    .C(_09331_),
    .X(_09334_));
 sky130_fd_sc_hd__o2bb2a_1 _16240_ (.A1_N(_09332_),
    .A2_N(_09333_),
    .B1(_09204_),
    .B2(_09334_),
    .X(_09335_));
 sky130_fd_sc_hd__xor2_2 _16241_ (.A(_09327_),
    .B(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(_09200_),
    .B(_09204_),
    .Y(_09337_));
 sky130_fd_sc_hd__a21oi_1 _16243_ (.A1(_09199_),
    .A2(_09205_),
    .B1(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__xnor2_2 _16244_ (.A(_09336_),
    .B(_09338_),
    .Y(_09339_));
 sky130_fd_sc_hd__xnor2_2 _16245_ (.A(_09323_),
    .B(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__and2b_1 _16246_ (.A_N(_09206_),
    .B(_09207_),
    .X(_09341_));
 sky130_fd_sc_hd__a21o_1 _16247_ (.A1(_09196_),
    .A2(_09208_),
    .B1(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__xnor2_1 _16248_ (.A(_09340_),
    .B(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__xnor2_2 _16249_ (.A(_09317_),
    .B(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__nor2_1 _16250_ (.A(_09209_),
    .B(_09210_),
    .Y(_09345_));
 sky130_fd_sc_hd__a21oi_2 _16251_ (.A1(_09189_),
    .A2(_09211_),
    .B1(_09345_),
    .Y(_09346_));
 sky130_fd_sc_hd__nor2_1 _16252_ (.A(_09344_),
    .B(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__and2_1 _16253_ (.A(_09344_),
    .B(_09346_),
    .X(_09348_));
 sky130_fd_sc_hd__nor2_1 _16254_ (.A(_09347_),
    .B(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__xnor2_1 _16255_ (.A(_09309_),
    .B(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__or2b_1 _16256_ (.A(_09213_),
    .B_N(_09212_),
    .X(_09351_));
 sky130_fd_sc_hd__a21boi_1 _16257_ (.A1(_09179_),
    .A2(_09214_),
    .B1_N(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__nor2_1 _16258_ (.A(_09350_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__and2_1 _16259_ (.A(_09350_),
    .B(_09352_),
    .X(_09354_));
 sky130_fd_sc_hd__nor2_1 _16260_ (.A(_09353_),
    .B(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__xnor2_1 _16261_ (.A(_09287_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__a21oi_1 _16262_ (.A1(_09218_),
    .A2(_09236_),
    .B1(_09217_),
    .Y(_09357_));
 sky130_fd_sc_hd__nor2_1 _16263_ (.A(_09356_),
    .B(_09357_),
    .Y(_09358_));
 sky130_fd_sc_hd__nand2_1 _16264_ (.A(_09356_),
    .B(_09357_),
    .Y(_09359_));
 sky130_fd_sc_hd__and2b_1 _16265_ (.A_N(_09358_),
    .B(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__xnor2_4 _16266_ (.A(_09234_),
    .B(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__a21o_1 _16267_ (.A1(_09238_),
    .A2(_09239_),
    .B1(_09237_),
    .X(_09362_));
 sky130_fd_sc_hd__a21boi_4 _16268_ (.A1(_09140_),
    .A2(_09241_),
    .B1_N(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__xnor2_4 _16269_ (.A(_09361_),
    .B(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__xor2_4 _16270_ (.A(_09272_),
    .B(_09364_),
    .X(_09365_));
 sky130_fd_sc_hd__xnor2_4 _16271_ (.A(_09271_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__mux2_1 _16272_ (.A0(\rbzero.debug_overlay.playerY[-5] ),
    .A1(\rbzero.debug_overlay.playerX[-5] ),
    .S(_08263_),
    .X(_09367_));
 sky130_fd_sc_hd__xnor2_1 _16273_ (.A(_09366_),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__a21oi_1 _16274_ (.A1(_09252_),
    .A2(_09263_),
    .B1(_09250_),
    .Y(_09369_));
 sky130_fd_sc_hd__xnor2_1 _16275_ (.A(_09368_),
    .B(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__o21ai_1 _16276_ (.A1(_09268_),
    .A2(_09370_),
    .B1(_08270_),
    .Y(_09371_));
 sky130_fd_sc_hd__a21o_1 _16277_ (.A1(_09268_),
    .A2(_09370_),
    .B1(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__o211a_1 _16278_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_08270_),
    .B1(_09372_),
    .C1(_08211_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _16279_ (.A0(_08461_),
    .A1(_08456_),
    .S(_08263_),
    .X(_09373_));
 sky130_fd_sc_hd__a31o_1 _16280_ (.A1(_09137_),
    .A2(_09230_),
    .A3(_09286_),
    .B1(_09284_),
    .X(_09374_));
 sky130_fd_sc_hd__or2b_1 _16281_ (.A(_09308_),
    .B_N(_09288_),
    .X(_09375_));
 sky130_fd_sc_hd__nand2_1 _16282_ (.A(_09306_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand2_2 _16283_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08543_),
    .Y(_09377_));
 sky130_fd_sc_hd__clkbuf_4 _16284_ (.A(_09377_),
    .X(_09378_));
 sky130_fd_sc_hd__nor2_1 _16285_ (.A(_08550_),
    .B(_09378_),
    .Y(_09379_));
 sky130_fd_sc_hd__or3_1 _16286_ (.A(_09135_),
    .B(_09133_),
    .C(_09223_),
    .X(_09380_));
 sky130_fd_sc_hd__a21bo_1 _16287_ (.A1(_09275_),
    .A2(_09277_),
    .B1_N(_09380_),
    .X(_09381_));
 sky130_fd_sc_hd__nor2_1 _16288_ (.A(_08616_),
    .B(_09222_),
    .Y(_09382_));
 sky130_fd_sc_hd__nor2_1 _16289_ (.A(_08967_),
    .B(_09132_),
    .Y(_09383_));
 sky130_fd_sc_hd__xnor2_1 _16290_ (.A(_09382_),
    .B(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__or3_1 _16291_ (.A(_08560_),
    .B(_09276_),
    .C(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__o21ai_1 _16292_ (.A1(_08561_),
    .A2(_09276_),
    .B1(_09384_),
    .Y(_09386_));
 sky130_fd_sc_hd__nand2_1 _16293_ (.A(_09385_),
    .B(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__a21o_1 _16294_ (.A1(_09293_),
    .A2(_09294_),
    .B1(_09291_),
    .X(_09388_));
 sky130_fd_sc_hd__or2b_1 _16295_ (.A(_09387_),
    .B_N(_09388_),
    .X(_09389_));
 sky130_fd_sc_hd__or2b_1 _16296_ (.A(_09388_),
    .B_N(_09387_),
    .X(_09390_));
 sky130_fd_sc_hd__nand2_1 _16297_ (.A(_09389_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__xnor2_1 _16298_ (.A(_09381_),
    .B(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__o21ba_1 _16299_ (.A1(_09224_),
    .A2(_09280_),
    .B1_N(_09279_),
    .X(_09393_));
 sky130_fd_sc_hd__xor2_1 _16300_ (.A(_09392_),
    .B(_09393_),
    .X(_09394_));
 sky130_fd_sc_hd__and2_1 _16301_ (.A(_09379_),
    .B(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__nor2_1 _16302_ (.A(_09379_),
    .B(_09394_),
    .Y(_09396_));
 sky130_fd_sc_hd__or2_1 _16303_ (.A(_09395_),
    .B(_09396_),
    .X(_09397_));
 sky130_fd_sc_hd__xor2_1 _16304_ (.A(_09376_),
    .B(_09397_),
    .X(_09398_));
 sky130_fd_sc_hd__or3b_1 _16305_ (.A(_09279_),
    .B(_09280_),
    .C_N(_09228_),
    .X(_09399_));
 sky130_fd_sc_hd__xor2_1 _16306_ (.A(_09398_),
    .B(_09399_),
    .X(_09400_));
 sky130_fd_sc_hd__a21o_1 _16307_ (.A1(_09295_),
    .A2(_09304_),
    .B1(_09302_),
    .X(_09401_));
 sky130_fd_sc_hd__or2b_1 _16308_ (.A(_09316_),
    .B_N(_09310_),
    .X(_09402_));
 sky130_fd_sc_hd__a21bo_1 _16309_ (.A1(_09311_),
    .A2(_09315_),
    .B1_N(_09402_),
    .X(_09403_));
 sky130_fd_sc_hd__buf_2 _16310_ (.A(_08888_),
    .X(_09404_));
 sky130_fd_sc_hd__or3_1 _16311_ (.A(_06461_),
    .B(_09106_),
    .C(_08829_),
    .X(_09405_));
 sky130_fd_sc_hd__clkbuf_4 _16312_ (.A(_08829_),
    .X(_09406_));
 sky130_fd_sc_hd__o22ai_1 _16313_ (.A1(_08545_),
    .A2(_09406_),
    .B1(_08888_),
    .B2(_09158_),
    .Y(_09407_));
 sky130_fd_sc_hd__o21ai_1 _16314_ (.A1(_09404_),
    .A2(_09405_),
    .B1(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__buf_2 _16315_ (.A(_08922_),
    .X(_09409_));
 sky130_fd_sc_hd__nor2_1 _16316_ (.A(_09409_),
    .B(_08620_),
    .Y(_09410_));
 sky130_fd_sc_hd__xnor2_2 _16317_ (.A(_09408_),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__nor2_1 _16318_ (.A(_08590_),
    .B(_08351_),
    .Y(_09412_));
 sky130_fd_sc_hd__o22a_1 _16319_ (.A1(_08424_),
    .A2(_08590_),
    .B1(_08351_),
    .B2(_08674_),
    .X(_09413_));
 sky130_fd_sc_hd__a21o_1 _16320_ (.A1(_09296_),
    .A2(_09412_),
    .B1(_09413_),
    .X(_09414_));
 sky130_fd_sc_hd__or2_1 _16321_ (.A(_08486_),
    .B(_08602_),
    .X(_09415_));
 sky130_fd_sc_hd__xnor2_1 _16322_ (.A(_09414_),
    .B(_09415_),
    .Y(_09416_));
 sky130_fd_sc_hd__clkbuf_4 _16323_ (.A(_08602_),
    .X(_09417_));
 sky130_fd_sc_hd__nand2_1 _16324_ (.A(_09165_),
    .B(_09296_),
    .Y(_09418_));
 sky130_fd_sc_hd__o31a_1 _16325_ (.A1(_08444_),
    .A2(_09417_),
    .A3(_09297_),
    .B1(_09418_),
    .X(_09419_));
 sky130_fd_sc_hd__nor2_1 _16326_ (.A(_09416_),
    .B(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__and2_1 _16327_ (.A(_09416_),
    .B(_09419_),
    .X(_09421_));
 sky130_fd_sc_hd__nor2_1 _16328_ (.A(_09420_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__xor2_2 _16329_ (.A(_09411_),
    .B(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__xnor2_1 _16330_ (.A(_09403_),
    .B(_09423_),
    .Y(_09424_));
 sky130_fd_sc_hd__xnor2_1 _16331_ (.A(_09401_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__clkinv_2 _16332_ (.A(_09312_),
    .Y(_09426_));
 sky130_fd_sc_hd__a2bb2o_1 _16333_ (.A1_N(_09182_),
    .A2_N(_09426_),
    .B1(_09313_),
    .B2(_09314_),
    .X(_09427_));
 sky130_fd_sc_hd__a22o_1 _16334_ (.A1(_09319_),
    .A2(_09320_),
    .B1(_09322_),
    .B2(_09318_),
    .X(_09428_));
 sky130_fd_sc_hd__nor2_1 _16335_ (.A(_08465_),
    .B(_08362_),
    .Y(_09429_));
 sky130_fd_sc_hd__o22a_1 _16336_ (.A1(_08487_),
    .A2(_08387_),
    .B1(_09064_),
    .B2(_08452_),
    .X(_09430_));
 sky130_fd_sc_hd__a21o_1 _16337_ (.A1(_09312_),
    .A2(_09429_),
    .B1(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__or2_1 _16338_ (.A(_08485_),
    .B(_08407_),
    .X(_09432_));
 sky130_fd_sc_hd__xor2_1 _16339_ (.A(_09431_),
    .B(_09432_),
    .X(_09433_));
 sky130_fd_sc_hd__and2_1 _16340_ (.A(_09428_),
    .B(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__or2_1 _16341_ (.A(_09428_),
    .B(_09433_),
    .X(_09435_));
 sky130_fd_sc_hd__or2b_1 _16342_ (.A(_09434_),
    .B_N(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__xnor2_1 _16343_ (.A(_09427_),
    .B(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__or2b_1 _16344_ (.A(_09338_),
    .B_N(_09336_),
    .X(_09438_));
 sky130_fd_sc_hd__nand2_1 _16345_ (.A(_09323_),
    .B(_09339_),
    .Y(_09439_));
 sky130_fd_sc_hd__nor2_1 _16346_ (.A(_08492_),
    .B(_09192_),
    .Y(_09440_));
 sky130_fd_sc_hd__nor2_1 _16347_ (.A(_08413_),
    .B(_09325_),
    .Y(_09441_));
 sky130_fd_sc_hd__xnor2_1 _16348_ (.A(_09320_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__xnor2_1 _16349_ (.A(_09440_),
    .B(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__nand2_1 _16350_ (.A(\rbzero.wall_tracer.stepDistY[5] ),
    .B(_08390_),
    .Y(_09444_));
 sky130_fd_sc_hd__a21o_1 _16351_ (.A1(_09203_),
    .A2(_09444_),
    .B1(_06100_),
    .X(_09445_));
 sky130_fd_sc_hd__clkbuf_4 _16352_ (.A(_09445_),
    .X(_09446_));
 sky130_fd_sc_hd__nand2_1 _16353_ (.A(\rbzero.wall_tracer.stepDistX[5] ),
    .B(_06101_),
    .Y(_09447_));
 sky130_fd_sc_hd__a21oi_1 _16354_ (.A1(_09446_),
    .A2(_09447_),
    .B1(_08366_),
    .Y(_09448_));
 sky130_fd_sc_hd__or2_1 _16355_ (.A(_08142_),
    .B(_08145_),
    .X(_09449_));
 sky130_fd_sc_hd__or4_1 _16356_ (.A(_08140_),
    .B(_08149_),
    .C(_08368_),
    .D(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__inv_2 _16357_ (.A(_08149_),
    .Y(_09451_));
 sky130_fd_sc_hd__a31o_1 _16358_ (.A1(_09073_),
    .A2(_09074_),
    .A3(_09329_),
    .B1(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__a31o_1 _16359_ (.A1(_08355_),
    .A2(_09450_),
    .A3(_09452_),
    .B1(_08371_),
    .X(_09453_));
 sky130_fd_sc_hd__or3b_2 _16360_ (.A(_08390_),
    .B(_09453_),
    .C_N(_08164_),
    .X(_09454_));
 sky130_fd_sc_hd__xor2_1 _16361_ (.A(_09334_),
    .B(_09454_),
    .X(_09455_));
 sky130_fd_sc_hd__xor2_1 _16362_ (.A(_09448_),
    .B(_09455_),
    .X(_09456_));
 sky130_fd_sc_hd__nor2_1 _16363_ (.A(_09204_),
    .B(_09334_),
    .Y(_09457_));
 sky130_fd_sc_hd__a21o_1 _16364_ (.A1(_09327_),
    .A2(_09335_),
    .B1(_09457_),
    .X(_09458_));
 sky130_fd_sc_hd__xor2_1 _16365_ (.A(_09456_),
    .B(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__xnor2_1 _16366_ (.A(_09443_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__a21oi_1 _16367_ (.A1(_09438_),
    .A2(_09439_),
    .B1(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__and3_1 _16368_ (.A(_09438_),
    .B(_09439_),
    .C(_09460_),
    .X(_09462_));
 sky130_fd_sc_hd__nor2_1 _16369_ (.A(_09461_),
    .B(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__xnor2_1 _16370_ (.A(_09437_),
    .B(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__and2b_1 _16371_ (.A_N(_09340_),
    .B(_09342_),
    .X(_09465_));
 sky130_fd_sc_hd__a21oi_1 _16372_ (.A1(_09317_),
    .A2(_09343_),
    .B1(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__nor2_1 _16373_ (.A(_09464_),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__and2_1 _16374_ (.A(_09464_),
    .B(_09466_),
    .X(_09468_));
 sky130_fd_sc_hd__nor2_1 _16375_ (.A(_09467_),
    .B(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__xnor2_1 _16376_ (.A(_09425_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__a21oi_1 _16377_ (.A1(_09309_),
    .A2(_09349_),
    .B1(_09347_),
    .Y(_09471_));
 sky130_fd_sc_hd__xor2_1 _16378_ (.A(_09470_),
    .B(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__xnor2_1 _16379_ (.A(_09400_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__a21oi_1 _16380_ (.A1(_09287_),
    .A2(_09355_),
    .B1(_09353_),
    .Y(_09474_));
 sky130_fd_sc_hd__nor2_1 _16381_ (.A(_09473_),
    .B(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__and2_1 _16382_ (.A(_09473_),
    .B(_09474_),
    .X(_09476_));
 sky130_fd_sc_hd__nor2_1 _16383_ (.A(_09475_),
    .B(_09476_),
    .Y(_09477_));
 sky130_fd_sc_hd__xnor2_1 _16384_ (.A(_09374_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__a21oi_1 _16385_ (.A1(_09234_),
    .A2(_09359_),
    .B1(_09358_),
    .Y(_09479_));
 sky130_fd_sc_hd__or2_2 _16386_ (.A(_09478_),
    .B(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__nand2_1 _16387_ (.A(_09478_),
    .B(_09479_),
    .Y(_09481_));
 sky130_fd_sc_hd__or4bb_1 _16388_ (.A(_09361_),
    .B(_09363_),
    .C_N(_09480_),
    .D_N(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__a2bb2o_1 _16389_ (.A1_N(_09361_),
    .A2_N(_09363_),
    .B1(_09480_),
    .B2(_09481_),
    .X(_09483_));
 sky130_fd_sc_hd__and2_2 _16390_ (.A(_09482_),
    .B(_09483_),
    .X(_09484_));
 sky130_fd_sc_hd__a21oi_1 _16391_ (.A1(_09272_),
    .A2(_09246_),
    .B1(_09364_),
    .Y(_09485_));
 sky130_fd_sc_hd__a31o_4 _16392_ (.A1(_09152_),
    .A2(_09248_),
    .A3(_09365_),
    .B1(_09485_),
    .X(_09486_));
 sky130_fd_sc_hd__xor2_4 _16393_ (.A(_09484_),
    .B(_09486_),
    .X(_09487_));
 sky130_fd_sc_hd__or2b_1 _16394_ (.A(_09373_),
    .B_N(_09487_),
    .X(_09488_));
 sky130_fd_sc_hd__or2b_1 _16395_ (.A(_09487_),
    .B_N(_09373_),
    .X(_09489_));
 sky130_fd_sc_hd__nand2_1 _16396_ (.A(_09488_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__nand2_1 _16397_ (.A(_09366_),
    .B(_09367_),
    .Y(_09491_));
 sky130_fd_sc_hd__o21a_1 _16398_ (.A1(_09368_),
    .A2(_09369_),
    .B1(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__xnor2_1 _16399_ (.A(_09490_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__xnor2_2 _16400_ (.A(_09268_),
    .B(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__or2_1 _16401_ (.A(\rbzero.texu_hot[2] ),
    .B(_08270_),
    .X(_09495_));
 sky130_fd_sc_hd__o211a_1 _16402_ (.A1(_08355_),
    .A2(_09494_),
    .B1(_09495_),
    .C1(_08211_),
    .X(_00468_));
 sky130_fd_sc_hd__a21boi_4 _16403_ (.A1(_09484_),
    .A2(_09486_),
    .B1_N(_09482_),
    .Y(_09496_));
 sky130_fd_sc_hd__a21o_1 _16404_ (.A1(_09306_),
    .A2(_09375_),
    .B1(_09397_),
    .X(_09497_));
 sky130_fd_sc_hd__o21ai_1 _16405_ (.A1(_09398_),
    .A2(_09399_),
    .B1(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__a21o_1 _16406_ (.A1(_09392_),
    .A2(_09393_),
    .B1(_09395_),
    .X(_09499_));
 sky130_fd_sc_hd__or2b_1 _16407_ (.A(_09424_),
    .B_N(_09401_),
    .X(_09500_));
 sky130_fd_sc_hd__a21bo_1 _16408_ (.A1(_09403_),
    .A2(_09423_),
    .B1_N(_09500_),
    .X(_09501_));
 sky130_fd_sc_hd__nand2_2 _16409_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08543_),
    .Y(_09502_));
 sky130_fd_sc_hd__clkbuf_4 _16410_ (.A(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__nor2_1 _16411_ (.A(_08561_),
    .B(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__o22a_1 _16412_ (.A1(_08561_),
    .A2(_09378_),
    .B1(_09503_),
    .B2(_08550_),
    .X(_09505_));
 sky130_fd_sc_hd__a21oi_1 _16413_ (.A1(_09379_),
    .A2(_09504_),
    .B1(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__a21bo_1 _16414_ (.A1(_09382_),
    .A2(_09383_),
    .B1_N(_09385_),
    .X(_09507_));
 sky130_fd_sc_hd__o22ai_1 _16415_ (.A1(_09409_),
    .A2(_09133_),
    .B1(_09225_),
    .B2(_09157_),
    .Y(_09508_));
 sky130_fd_sc_hd__or4_1 _16416_ (.A(_09409_),
    .B(_09157_),
    .C(_09133_),
    .D(_09225_),
    .X(_09509_));
 sky130_fd_sc_hd__nand2_1 _16417_ (.A(_09508_),
    .B(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__buf_4 _16418_ (.A(_09276_),
    .X(_09511_));
 sky130_fd_sc_hd__nor2_1 _16419_ (.A(_09135_),
    .B(_09511_),
    .Y(_09512_));
 sky130_fd_sc_hd__xor2_1 _16420_ (.A(_09510_),
    .B(_09512_),
    .X(_09513_));
 sky130_fd_sc_hd__a2bb2o_1 _16421_ (.A1_N(_09404_),
    .A2_N(_09405_),
    .B1(_09407_),
    .B2(_09410_),
    .X(_09514_));
 sky130_fd_sc_hd__and2b_1 _16422_ (.A_N(_09513_),
    .B(_09514_),
    .X(_09515_));
 sky130_fd_sc_hd__and2b_1 _16423_ (.A_N(_09514_),
    .B(_09513_),
    .X(_09516_));
 sky130_fd_sc_hd__nor2_1 _16424_ (.A(_09515_),
    .B(_09516_),
    .Y(_09517_));
 sky130_fd_sc_hd__xnor2_1 _16425_ (.A(_09507_),
    .B(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__inv_2 _16426_ (.A(_09381_),
    .Y(_09519_));
 sky130_fd_sc_hd__o21a_1 _16427_ (.A1(_09519_),
    .A2(_09391_),
    .B1(_09389_),
    .X(_09520_));
 sky130_fd_sc_hd__xor2_1 _16428_ (.A(_09518_),
    .B(_09520_),
    .X(_09521_));
 sky130_fd_sc_hd__xor2_1 _16429_ (.A(_09506_),
    .B(_09521_),
    .X(_09522_));
 sky130_fd_sc_hd__xnor2_1 _16430_ (.A(_09501_),
    .B(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__xnor2_1 _16431_ (.A(_09499_),
    .B(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__a21o_1 _16432_ (.A1(_09411_),
    .A2(_09422_),
    .B1(_09420_),
    .X(_09525_));
 sky130_fd_sc_hd__clkbuf_4 _16433_ (.A(_08783_),
    .X(_09526_));
 sky130_fd_sc_hd__o22ai_1 _16434_ (.A1(_08545_),
    .A2(_09526_),
    .B1(_08829_),
    .B2(_09158_),
    .Y(_09527_));
 sky130_fd_sc_hd__or2_1 _16435_ (.A(_08783_),
    .B(_09405_),
    .X(_09528_));
 sky130_fd_sc_hd__nand2_1 _16436_ (.A(_09527_),
    .B(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__or3_1 _16437_ (.A(_08888_),
    .B(_08620_),
    .C(_09529_),
    .X(_09530_));
 sky130_fd_sc_hd__o21ai_1 _16438_ (.A1(_09404_),
    .A2(_09162_),
    .B1(_09529_),
    .Y(_09531_));
 sky130_fd_sc_hd__and2_1 _16439_ (.A(_09530_),
    .B(_09531_),
    .X(_09532_));
 sky130_fd_sc_hd__nor2_1 _16440_ (.A(_08674_),
    .B(_08407_),
    .Y(_09533_));
 sky130_fd_sc_hd__xnor2_1 _16441_ (.A(_09412_),
    .B(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__or2_1 _16442_ (.A(_08424_),
    .B(_08602_),
    .X(_09535_));
 sky130_fd_sc_hd__xnor2_1 _16443_ (.A(_09534_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__nand2_1 _16444_ (.A(_09296_),
    .B(_09412_),
    .Y(_09537_));
 sky130_fd_sc_hd__o31a_1 _16445_ (.A1(_08486_),
    .A2(_08602_),
    .A3(_09413_),
    .B1(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__nor2_1 _16446_ (.A(_09536_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__and2_1 _16447_ (.A(_09536_),
    .B(_09538_),
    .X(_09540_));
 sky130_fd_sc_hd__nor2_1 _16448_ (.A(_09539_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__xnor2_1 _16449_ (.A(_09532_),
    .B(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__a21o_1 _16450_ (.A1(_09427_),
    .A2(_09435_),
    .B1(_09434_),
    .X(_09543_));
 sky130_fd_sc_hd__or2b_1 _16451_ (.A(_09542_),
    .B_N(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__or2b_1 _16452_ (.A(_09543_),
    .B_N(_09542_),
    .X(_09545_));
 sky130_fd_sc_hd__nand2_1 _16453_ (.A(_09544_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__xnor2_1 _16454_ (.A(_09525_),
    .B(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__a2bb2o_1 _16455_ (.A1_N(_09430_),
    .A2_N(_09432_),
    .B1(_09312_),
    .B2(_09429_),
    .X(_09548_));
 sky130_fd_sc_hd__nand2_1 _16456_ (.A(_09320_),
    .B(_09441_),
    .Y(_09549_));
 sky130_fd_sc_hd__o31a_1 _16457_ (.A1(_08492_),
    .A2(_09192_),
    .A3(_09442_),
    .B1(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__nor2_1 _16458_ (.A(_08495_),
    .B(_09064_),
    .Y(_09551_));
 sky130_fd_sc_hd__nor2_1 _16459_ (.A(_08487_),
    .B(_09192_),
    .Y(_09552_));
 sky130_fd_sc_hd__o21ba_1 _16460_ (.A1(_08495_),
    .A2(_09071_),
    .B1_N(_09429_),
    .X(_09553_));
 sky130_fd_sc_hd__a21o_1 _16461_ (.A1(_09551_),
    .A2(_09552_),
    .B1(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__or2_1 _16462_ (.A(_08485_),
    .B(_08387_),
    .X(_09555_));
 sky130_fd_sc_hd__xnor2_1 _16463_ (.A(_09554_),
    .B(_09555_),
    .Y(_09556_));
 sky130_fd_sc_hd__xnor2_1 _16464_ (.A(_09550_),
    .B(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__xnor2_1 _16465_ (.A(_09548_),
    .B(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__nor2_1 _16466_ (.A(_08492_),
    .B(_09198_),
    .Y(_09559_));
 sky130_fd_sc_hd__nor2_1 _16467_ (.A(_09002_),
    .B(_09326_),
    .Y(_09560_));
 sky130_fd_sc_hd__a21oi_2 _16468_ (.A1(_09446_),
    .A2(_09447_),
    .B1(_08977_),
    .Y(_09561_));
 sky130_fd_sc_hd__xor2_1 _16469_ (.A(_09560_),
    .B(_09561_),
    .X(_09562_));
 sky130_fd_sc_hd__xor2_1 _16470_ (.A(_09559_),
    .B(_09562_),
    .X(_09563_));
 sky130_fd_sc_hd__nand2_1 _16471_ (.A(\rbzero.wall_tracer.stepDistY[6] ),
    .B(_09069_),
    .Y(_09564_));
 sky130_fd_sc_hd__a21o_2 _16472_ (.A1(_09564_),
    .A2(_09331_),
    .B1(_06100_),
    .X(_09565_));
 sky130_fd_sc_hd__nand2_1 _16473_ (.A(\rbzero.wall_tracer.stepDistX[6] ),
    .B(_06101_),
    .Y(_09566_));
 sky130_fd_sc_hd__and2_1 _16474_ (.A(_09565_),
    .B(_09566_),
    .X(_09567_));
 sky130_fd_sc_hd__inv_2 _16475_ (.A(_08152_),
    .Y(_09568_));
 sky130_fd_sc_hd__and4_1 _16476_ (.A(_09073_),
    .B(_09451_),
    .C(_09074_),
    .D(_09329_),
    .X(_09569_));
 sky130_fd_sc_hd__o41a_1 _16477_ (.A1(_08140_),
    .A2(_08149_),
    .A3(_08368_),
    .A4(_09449_),
    .B1(_08153_),
    .X(_09570_));
 sky130_fd_sc_hd__a211o_1 _16478_ (.A1(_09568_),
    .A2(_09569_),
    .B1(_09570_),
    .C1(_08270_),
    .X(_09571_));
 sky130_fd_sc_hd__a22o_4 _16479_ (.A1(\rbzero.wall_tracer.stepDistY[8] ),
    .A2(_09069_),
    .B1(_09072_),
    .B2(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__or3b_1 _16480_ (.A(_08383_),
    .B(_09454_),
    .C_N(_09572_),
    .X(_09573_));
 sky130_fd_sc_hd__nand2_1 _16481_ (.A(\rbzero.wall_tracer.stepDistY[7] ),
    .B(_09069_),
    .Y(_09574_));
 sky130_fd_sc_hd__nand2_1 _16482_ (.A(_09574_),
    .B(_09453_),
    .Y(_09575_));
 sky130_fd_sc_hd__a22o_1 _16483_ (.A1(_08404_),
    .A2(_09575_),
    .B1(_09572_),
    .B2(_08403_),
    .X(_09576_));
 sky130_fd_sc_hd__or4bb_1 _16484_ (.A(_08965_),
    .B(_09567_),
    .C_N(_09573_),
    .D_N(_09576_),
    .X(_09577_));
 sky130_fd_sc_hd__a2bb2o_1 _16485_ (.A1_N(_08965_),
    .A2_N(_09567_),
    .B1(_09573_),
    .B2(_09576_),
    .X(_09578_));
 sky130_fd_sc_hd__nor2_1 _16486_ (.A(_09334_),
    .B(_09454_),
    .Y(_09579_));
 sky130_fd_sc_hd__a21o_1 _16487_ (.A1(_09448_),
    .A2(_09455_),
    .B1(_09579_),
    .X(_09580_));
 sky130_fd_sc_hd__nand3_1 _16488_ (.A(_09577_),
    .B(_09578_),
    .C(_09580_),
    .Y(_09581_));
 sky130_fd_sc_hd__a21o_1 _16489_ (.A1(_09577_),
    .A2(_09578_),
    .B1(_09580_),
    .X(_09582_));
 sky130_fd_sc_hd__nand3_1 _16490_ (.A(_09563_),
    .B(_09581_),
    .C(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__a21o_1 _16491_ (.A1(_09581_),
    .A2(_09582_),
    .B1(_09563_),
    .X(_09584_));
 sky130_fd_sc_hd__and2_1 _16492_ (.A(_09456_),
    .B(_09458_),
    .X(_09585_));
 sky130_fd_sc_hd__a21o_1 _16493_ (.A1(_09443_),
    .A2(_09459_),
    .B1(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__nand3_1 _16494_ (.A(_09583_),
    .B(_09584_),
    .C(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__a21o_1 _16495_ (.A1(_09583_),
    .A2(_09584_),
    .B1(_09586_),
    .X(_09588_));
 sky130_fd_sc_hd__and3_1 _16496_ (.A(_09558_),
    .B(_09587_),
    .C(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__a21oi_1 _16497_ (.A1(_09587_),
    .A2(_09588_),
    .B1(_09558_),
    .Y(_09590_));
 sky130_fd_sc_hd__or2_1 _16498_ (.A(_09589_),
    .B(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__a21oi_1 _16499_ (.A1(_09437_),
    .A2(_09463_),
    .B1(_09461_),
    .Y(_09592_));
 sky130_fd_sc_hd__xor2_1 _16500_ (.A(_09591_),
    .B(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__nand2_1 _16501_ (.A(_09547_),
    .B(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__or2_1 _16502_ (.A(_09547_),
    .B(_09593_),
    .X(_09595_));
 sky130_fd_sc_hd__nand2_1 _16503_ (.A(_09594_),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__a21oi_1 _16504_ (.A1(_09425_),
    .A2(_09469_),
    .B1(_09467_),
    .Y(_09597_));
 sky130_fd_sc_hd__xor2_1 _16505_ (.A(_09596_),
    .B(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__nand2_1 _16506_ (.A(_09524_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__or2_1 _16507_ (.A(_09524_),
    .B(_09598_),
    .X(_09600_));
 sky130_fd_sc_hd__nand2_1 _16508_ (.A(_09599_),
    .B(_09600_),
    .Y(_09601_));
 sky130_fd_sc_hd__nor2_1 _16509_ (.A(_09470_),
    .B(_09471_),
    .Y(_09602_));
 sky130_fd_sc_hd__a21oi_1 _16510_ (.A1(_09400_),
    .A2(_09472_),
    .B1(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__xnor2_1 _16511_ (.A(_09601_),
    .B(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__xor2_1 _16512_ (.A(_09498_),
    .B(_09604_),
    .X(_09605_));
 sky130_fd_sc_hd__a21oi_1 _16513_ (.A1(_09374_),
    .A2(_09477_),
    .B1(_09475_),
    .Y(_09606_));
 sky130_fd_sc_hd__nor2_1 _16514_ (.A(_09605_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__and2_1 _16515_ (.A(_09605_),
    .B(_09606_),
    .X(_09608_));
 sky130_fd_sc_hd__or2_2 _16516_ (.A(_09607_),
    .B(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__xor2_4 _16517_ (.A(_09480_),
    .B(_09609_),
    .X(_09610_));
 sky130_fd_sc_hd__xor2_4 _16518_ (.A(_09496_),
    .B(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__clkinv_2 _16519_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .Y(_09612_));
 sky130_fd_sc_hd__mux2_1 _16520_ (.A0(_04856_),
    .A1(_09612_),
    .S(_08263_),
    .X(_09613_));
 sky130_fd_sc_hd__nor2_1 _16521_ (.A(_09611_),
    .B(_09613_),
    .Y(_09614_));
 sky130_fd_sc_hd__and2_1 _16522_ (.A(_09611_),
    .B(_09613_),
    .X(_09615_));
 sky130_fd_sc_hd__or2_1 _16523_ (.A(_09614_),
    .B(_09615_),
    .X(_09616_));
 sky130_fd_sc_hd__o21a_1 _16524_ (.A1(_09490_),
    .A2(_09492_),
    .B1(_09488_),
    .X(_09617_));
 sky130_fd_sc_hd__xnor2_1 _16525_ (.A(_09616_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__o21ai_1 _16526_ (.A1(_09268_),
    .A2(_09618_),
    .B1(_08270_),
    .Y(_09619_));
 sky130_fd_sc_hd__a21o_1 _16527_ (.A1(_09268_),
    .A2(_09618_),
    .B1(_09619_),
    .X(_09620_));
 sky130_fd_sc_hd__o211a_1 _16528_ (.A1(\rbzero.texu_hot[3] ),
    .A2(_08270_),
    .B1(_09620_),
    .C1(_08211_),
    .X(_00469_));
 sky130_fd_sc_hd__o21ba_1 _16529_ (.A1(_09616_),
    .A2(_09617_),
    .B1_N(_09614_),
    .X(_09621_));
 sky130_fd_sc_hd__a21oi_1 _16530_ (.A1(_09480_),
    .A2(_09482_),
    .B1(_09609_),
    .Y(_09622_));
 sky130_fd_sc_hd__a31oi_4 _16531_ (.A1(_09484_),
    .A2(_09486_),
    .A3(_09610_),
    .B1(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__or2b_1 _16532_ (.A(_09604_),
    .B_N(_09498_),
    .X(_09624_));
 sky130_fd_sc_hd__o21ai_1 _16533_ (.A1(_09601_),
    .A2(_09603_),
    .B1(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__or2b_1 _16534_ (.A(_09523_),
    .B_N(_09499_),
    .X(_09626_));
 sky130_fd_sc_hd__a21bo_1 _16535_ (.A1(_09501_),
    .A2(_09522_),
    .B1_N(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__or2_1 _16536_ (.A(_09596_),
    .B(_09597_),
    .X(_09628_));
 sky130_fd_sc_hd__a2bb2o_1 _16537_ (.A1_N(_09518_),
    .A2_N(_09520_),
    .B1(_09521_),
    .B2(_09506_),
    .X(_09629_));
 sky130_fd_sc_hd__or2b_1 _16538_ (.A(_09546_),
    .B_N(_09525_),
    .X(_09630_));
 sky130_fd_sc_hd__nand2_1 _16539_ (.A(_09379_),
    .B(_09504_),
    .Y(_09631_));
 sky130_fd_sc_hd__nor2_1 _16540_ (.A(_08561_),
    .B(_09378_),
    .Y(_09632_));
 sky130_fd_sc_hd__nor2_1 _16541_ (.A(_09135_),
    .B(_09503_),
    .Y(_09633_));
 sky130_fd_sc_hd__o22a_1 _16542_ (.A1(_09135_),
    .A2(_09378_),
    .B1(_09503_),
    .B2(_08561_),
    .X(_09634_));
 sky130_fd_sc_hd__a21o_1 _16543_ (.A1(_09632_),
    .A2(_09633_),
    .B1(_09634_),
    .X(_09635_));
 sky130_fd_sc_hd__nand2_2 _16544_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_08543_),
    .Y(_09636_));
 sky130_fd_sc_hd__clkbuf_4 _16545_ (.A(_09636_),
    .X(_09637_));
 sky130_fd_sc_hd__nor2_1 _16546_ (.A(_08550_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__xnor2_1 _16547_ (.A(_09635_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__xnor2_1 _16548_ (.A(_09631_),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__a21bo_1 _16549_ (.A1(_09508_),
    .A2(_09512_),
    .B1_N(_09509_),
    .X(_09641_));
 sky130_fd_sc_hd__nor2_1 _16550_ (.A(_09157_),
    .B(_09276_),
    .Y(_09642_));
 sky130_fd_sc_hd__o22a_1 _16551_ (.A1(_08888_),
    .A2(_09133_),
    .B1(_09225_),
    .B2(_09409_),
    .X(_09643_));
 sky130_fd_sc_hd__or2_1 _16552_ (.A(_08888_),
    .B(_09222_),
    .X(_09644_));
 sky130_fd_sc_hd__or3_1 _16553_ (.A(_08922_),
    .B(_09132_),
    .C(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__and2b_1 _16554_ (.A_N(_09643_),
    .B(_09645_),
    .X(_09646_));
 sky130_fd_sc_hd__xnor2_1 _16555_ (.A(_09642_),
    .B(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__a21oi_1 _16556_ (.A1(_09528_),
    .A2(_09530_),
    .B1(_09647_),
    .Y(_09648_));
 sky130_fd_sc_hd__and3_1 _16557_ (.A(_09528_),
    .B(_09530_),
    .C(_09647_),
    .X(_09649_));
 sky130_fd_sc_hd__nor2_1 _16558_ (.A(_09648_),
    .B(_09649_),
    .Y(_09650_));
 sky130_fd_sc_hd__xnor2_1 _16559_ (.A(_09641_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__a21oi_1 _16560_ (.A1(_09507_),
    .A2(_09517_),
    .B1(_09515_),
    .Y(_09652_));
 sky130_fd_sc_hd__nor2_1 _16561_ (.A(_09651_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__and2_1 _16562_ (.A(_09651_),
    .B(_09652_),
    .X(_09654_));
 sky130_fd_sc_hd__nor2_1 _16563_ (.A(_09653_),
    .B(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__xnor2_1 _16564_ (.A(_09640_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__a21o_1 _16565_ (.A1(_09544_),
    .A2(_09630_),
    .B1(_09656_),
    .X(_09657_));
 sky130_fd_sc_hd__nand3_1 _16566_ (.A(_09544_),
    .B(_09630_),
    .C(_09656_),
    .Y(_09658_));
 sky130_fd_sc_hd__nand2_1 _16567_ (.A(_09657_),
    .B(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__xnor2_1 _16568_ (.A(_09629_),
    .B(_09659_),
    .Y(_09660_));
 sky130_fd_sc_hd__or2_1 _16569_ (.A(_09591_),
    .B(_09592_),
    .X(_09661_));
 sky130_fd_sc_hd__a21o_1 _16570_ (.A1(_09532_),
    .A2(_09541_),
    .B1(_09539_),
    .X(_09662_));
 sky130_fd_sc_hd__or2b_1 _16571_ (.A(_09557_),
    .B_N(_09548_),
    .X(_09663_));
 sky130_fd_sc_hd__o21ai_2 _16572_ (.A1(_09550_),
    .A2(_09556_),
    .B1(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__nor2_1 _16573_ (.A(_08544_),
    .B(_08422_),
    .Y(_09665_));
 sky130_fd_sc_hd__nor2_1 _16574_ (.A(_09158_),
    .B(_08783_),
    .Y(_09666_));
 sky130_fd_sc_hd__xnor2_1 _16575_ (.A(_09665_),
    .B(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__or3_1 _16576_ (.A(_08829_),
    .B(_08620_),
    .C(_09667_),
    .X(_09668_));
 sky130_fd_sc_hd__o21ai_1 _16577_ (.A1(_09406_),
    .A2(_09162_),
    .B1(_09667_),
    .Y(_09669_));
 sky130_fd_sc_hd__and2_1 _16578_ (.A(_09668_),
    .B(_09669_),
    .X(_09670_));
 sky130_fd_sc_hd__clkbuf_4 _16579_ (.A(_08590_),
    .X(_09671_));
 sky130_fd_sc_hd__nor2_1 _16580_ (.A(_09671_),
    .B(_08387_),
    .Y(_09672_));
 sky130_fd_sc_hd__o22a_1 _16581_ (.A1(_08674_),
    .A2(_08387_),
    .B1(_08407_),
    .B2(_09671_),
    .X(_09673_));
 sky130_fd_sc_hd__a21oi_1 _16582_ (.A1(_09533_),
    .A2(_09672_),
    .B1(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__nor2_1 _16583_ (.A(_09417_),
    .B(_08351_),
    .Y(_09675_));
 sky130_fd_sc_hd__xnor2_1 _16584_ (.A(_09674_),
    .B(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__nand2_1 _16585_ (.A(_09412_),
    .B(_09533_),
    .Y(_09677_));
 sky130_fd_sc_hd__o31a_1 _16586_ (.A1(_08424_),
    .A2(_09417_),
    .A3(_09534_),
    .B1(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__nor2_1 _16587_ (.A(_09676_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__and2_1 _16588_ (.A(_09676_),
    .B(_09678_),
    .X(_09680_));
 sky130_fd_sc_hd__nor2_1 _16589_ (.A(_09679_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__xor2_1 _16590_ (.A(_09670_),
    .B(_09681_),
    .X(_09682_));
 sky130_fd_sc_hd__xnor2_1 _16591_ (.A(_09664_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__xnor2_1 _16592_ (.A(_09662_),
    .B(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__a2bb2o_1 _16593_ (.A1_N(_09553_),
    .A2_N(_09555_),
    .B1(_09551_),
    .B2(_09552_),
    .X(_09685_));
 sky130_fd_sc_hd__a22o_1 _16594_ (.A1(_09560_),
    .A2(_09561_),
    .B1(_09562_),
    .B2(_09559_),
    .X(_09686_));
 sky130_fd_sc_hd__nor2_1 _16595_ (.A(_08495_),
    .B(_09198_),
    .Y(_09687_));
 sky130_fd_sc_hd__xnor2_1 _16596_ (.A(_09552_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__or3_1 _16597_ (.A(_08533_),
    .B(_09064_),
    .C(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__o21ai_1 _16598_ (.A1(_08533_),
    .A2(_09064_),
    .B1(_09688_),
    .Y(_09690_));
 sky130_fd_sc_hd__and2_1 _16599_ (.A(_09689_),
    .B(_09690_),
    .X(_09691_));
 sky130_fd_sc_hd__xor2_2 _16600_ (.A(_09686_),
    .B(_09691_),
    .X(_09692_));
 sky130_fd_sc_hd__xor2_2 _16601_ (.A(_09685_),
    .B(_09692_),
    .X(_09693_));
 sky130_fd_sc_hd__or3b_1 _16602_ (.A(_09002_),
    .B(_09567_),
    .C_N(_09561_),
    .X(_09694_));
 sky130_fd_sc_hd__and2_1 _16603_ (.A(_09445_),
    .B(_09447_),
    .X(_09695_));
 sky130_fd_sc_hd__buf_2 _16604_ (.A(_09695_),
    .X(_09696_));
 sky130_fd_sc_hd__buf_2 _16605_ (.A(_09567_),
    .X(_09697_));
 sky130_fd_sc_hd__o22ai_1 _16606_ (.A1(_09002_),
    .A2(_09696_),
    .B1(_09697_),
    .B2(_08977_),
    .Y(_09698_));
 sky130_fd_sc_hd__nand2_1 _16607_ (.A(_09694_),
    .B(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__clkbuf_4 _16608_ (.A(_08344_),
    .X(_09700_));
 sky130_fd_sc_hd__nor2_1 _16609_ (.A(_09700_),
    .B(_09326_),
    .Y(_09701_));
 sky130_fd_sc_hd__xnor2_2 _16610_ (.A(_09699_),
    .B(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__a21o_1 _16611_ (.A1(_09574_),
    .A2(_09453_),
    .B1(_06101_),
    .X(_09703_));
 sky130_fd_sc_hd__nand2_1 _16612_ (.A(\rbzero.wall_tracer.stepDistX[7] ),
    .B(_06101_),
    .Y(_09704_));
 sky130_fd_sc_hd__and2_1 _16613_ (.A(_09703_),
    .B(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__buf_2 _16614_ (.A(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__nor2_1 _16615_ (.A(_08965_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand2_1 _16616_ (.A(_08404_),
    .B(_09572_),
    .Y(_09708_));
 sky130_fd_sc_hd__or3_1 _16617_ (.A(_08153_),
    .B(_08155_),
    .C(_09450_),
    .X(_09709_));
 sky130_fd_sc_hd__o21ai_1 _16618_ (.A1(_08153_),
    .A2(_09450_),
    .B1(_08155_),
    .Y(_09710_));
 sky130_fd_sc_hd__a31o_1 _16619_ (.A1(_08355_),
    .A2(_09709_),
    .A3(_09710_),
    .B1(_08371_),
    .X(_09711_));
 sky130_fd_sc_hd__or3b_1 _16620_ (.A(_08390_),
    .B(_09711_),
    .C_N(_08164_),
    .X(_09712_));
 sky130_fd_sc_hd__xor2_1 _16621_ (.A(_09708_),
    .B(_09712_),
    .X(_09713_));
 sky130_fd_sc_hd__xnor2_1 _16622_ (.A(_09707_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__nand2_1 _16623_ (.A(_09573_),
    .B(_09577_),
    .Y(_09715_));
 sky130_fd_sc_hd__xnor2_1 _16624_ (.A(_09714_),
    .B(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__xnor2_2 _16625_ (.A(_09702_),
    .B(_09716_),
    .Y(_09717_));
 sky130_fd_sc_hd__and2_1 _16626_ (.A(_09581_),
    .B(_09583_),
    .X(_09718_));
 sky130_fd_sc_hd__xor2_2 _16627_ (.A(_09717_),
    .B(_09718_),
    .X(_09719_));
 sky130_fd_sc_hd__xnor2_2 _16628_ (.A(_09693_),
    .B(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__a21boi_2 _16629_ (.A1(_09558_),
    .A2(_09588_),
    .B1_N(_09587_),
    .Y(_09721_));
 sky130_fd_sc_hd__nor2_1 _16630_ (.A(_09720_),
    .B(_09721_),
    .Y(_09722_));
 sky130_fd_sc_hd__nand2_1 _16631_ (.A(_09720_),
    .B(_09721_),
    .Y(_09723_));
 sky130_fd_sc_hd__and2b_1 _16632_ (.A_N(_09722_),
    .B(_09723_),
    .X(_09724_));
 sky130_fd_sc_hd__xnor2_1 _16633_ (.A(_09684_),
    .B(_09724_),
    .Y(_09725_));
 sky130_fd_sc_hd__a21oi_1 _16634_ (.A1(_09661_),
    .A2(_09594_),
    .B1(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__and3_1 _16635_ (.A(_09661_),
    .B(_09594_),
    .C(_09725_),
    .X(_09727_));
 sky130_fd_sc_hd__nor2_1 _16636_ (.A(_09726_),
    .B(_09727_),
    .Y(_09728_));
 sky130_fd_sc_hd__xnor2_1 _16637_ (.A(_09660_),
    .B(_09728_),
    .Y(_09729_));
 sky130_fd_sc_hd__a21oi_2 _16638_ (.A1(_09628_),
    .A2(_09599_),
    .B1(_09729_),
    .Y(_09730_));
 sky130_fd_sc_hd__and3_1 _16639_ (.A(_09628_),
    .B(_09599_),
    .C(_09729_),
    .X(_09731_));
 sky130_fd_sc_hd__nor2_1 _16640_ (.A(_09730_),
    .B(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__xnor2_1 _16641_ (.A(_09627_),
    .B(_09732_),
    .Y(_09733_));
 sky130_fd_sc_hd__xnor2_1 _16642_ (.A(_09625_),
    .B(_09733_),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_1 _16643_ (.A(_09607_),
    .B(_09734_),
    .Y(_09735_));
 sky130_fd_sc_hd__or2_1 _16644_ (.A(_09607_),
    .B(_09734_),
    .X(_09736_));
 sky130_fd_sc_hd__nand2_2 _16645_ (.A(_09735_),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__xor2_4 _16646_ (.A(_09623_),
    .B(_09737_),
    .X(_09738_));
 sky130_fd_sc_hd__mux2_1 _16647_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_08263_),
    .X(_09739_));
 sky130_fd_sc_hd__nor2_1 _16648_ (.A(_09738_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__and2_1 _16649_ (.A(_09738_),
    .B(_09739_),
    .X(_09741_));
 sky130_fd_sc_hd__nor2_1 _16650_ (.A(_09740_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__xnor2_1 _16651_ (.A(_09268_),
    .B(_09742_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand2_1 _16652_ (.A(_09621_),
    .B(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__or2_1 _16653_ (.A(_09621_),
    .B(_09743_),
    .X(_09745_));
 sky130_fd_sc_hd__a21o_1 _16654_ (.A1(_09744_),
    .A2(_09745_),
    .B1(_08355_),
    .X(_09746_));
 sky130_fd_sc_hd__o211a_1 _16655_ (.A1(\rbzero.texu_hot[4] ),
    .A2(_08270_),
    .B1(_09746_),
    .C1(_08211_),
    .X(_00470_));
 sky130_fd_sc_hd__o21ba_1 _16656_ (.A1(_09621_),
    .A2(_09740_),
    .B1_N(_09741_),
    .X(_09747_));
 sky130_fd_sc_hd__o21a_1 _16657_ (.A1(_09623_),
    .A2(_09737_),
    .B1(_09735_),
    .X(_09748_));
 sky130_fd_sc_hd__or2b_2 _16658_ (.A(_09733_),
    .B_N(_09625_),
    .X(_09749_));
 sky130_fd_sc_hd__or2b_1 _16659_ (.A(_09659_),
    .B_N(_09629_),
    .X(_09750_));
 sky130_fd_sc_hd__or2b_1 _16660_ (.A(_09631_),
    .B_N(_09639_),
    .X(_09751_));
 sky130_fd_sc_hd__a21oi_1 _16661_ (.A1(_09657_),
    .A2(_09750_),
    .B1(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__and3_1 _16662_ (.A(_09751_),
    .B(_09657_),
    .C(_09750_),
    .X(_09753_));
 sky130_fd_sc_hd__nor2_1 _16663_ (.A(_09752_),
    .B(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_4 _16664_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_08543_),
    .Y(_09755_));
 sky130_fd_sc_hd__or2_1 _16665_ (.A(_08548_),
    .B(_09755_),
    .X(_09756_));
 sky130_fd_sc_hd__xnor2_2 _16666_ (.A(_09754_),
    .B(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__a21o_1 _16667_ (.A1(_09640_),
    .A2(_09655_),
    .B1(_09653_),
    .X(_09758_));
 sky130_fd_sc_hd__nand2_1 _16668_ (.A(_09664_),
    .B(_09682_),
    .Y(_09759_));
 sky130_fd_sc_hd__or2b_1 _16669_ (.A(_09683_),
    .B_N(_09662_),
    .X(_09760_));
 sky130_fd_sc_hd__nor2_1 _16670_ (.A(_09409_),
    .B(_09377_),
    .Y(_09761_));
 sky130_fd_sc_hd__o22a_1 _16671_ (.A1(_09409_),
    .A2(_09511_),
    .B1(_09378_),
    .B2(_09157_),
    .X(_09762_));
 sky130_fd_sc_hd__a21oi_1 _16672_ (.A1(_09642_),
    .A2(_09761_),
    .B1(_09762_),
    .Y(_09763_));
 sky130_fd_sc_hd__xnor2_1 _16673_ (.A(_09633_),
    .B(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__nand2_1 _16674_ (.A(_09632_),
    .B(_09633_),
    .Y(_09765_));
 sky130_fd_sc_hd__o31a_1 _16675_ (.A1(_08550_),
    .A2(_09635_),
    .A3(_09637_),
    .B1(_09765_),
    .X(_09766_));
 sky130_fd_sc_hd__xor2_1 _16676_ (.A(_09764_),
    .B(_09766_),
    .X(_09767_));
 sky130_fd_sc_hd__clkbuf_4 _16677_ (.A(_09637_),
    .X(_09768_));
 sky130_fd_sc_hd__nor2_1 _16678_ (.A(_08561_),
    .B(_09768_),
    .Y(_09769_));
 sky130_fd_sc_hd__xor2_1 _16679_ (.A(_09767_),
    .B(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__a21bo_1 _16680_ (.A1(_09642_),
    .A2(_09646_),
    .B1_N(_09645_),
    .X(_09771_));
 sky130_fd_sc_hd__a21bo_1 _16681_ (.A1(_09665_),
    .A2(_09666_),
    .B1_N(_09668_),
    .X(_09772_));
 sky130_fd_sc_hd__or2_1 _16682_ (.A(_08783_),
    .B(_09132_),
    .X(_09773_));
 sky130_fd_sc_hd__o22ai_1 _16683_ (.A1(_09526_),
    .A2(_08620_),
    .B1(_09133_),
    .B2(_08829_),
    .Y(_09774_));
 sky130_fd_sc_hd__o31a_1 _16684_ (.A1(_09406_),
    .A2(_08620_),
    .A3(_09773_),
    .B1(_09774_),
    .X(_09775_));
 sky130_fd_sc_hd__xnor2_1 _16685_ (.A(_09644_),
    .B(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__and2_1 _16686_ (.A(_09772_),
    .B(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__or2_1 _16687_ (.A(_09772_),
    .B(_09776_),
    .X(_09778_));
 sky130_fd_sc_hd__and2b_1 _16688_ (.A_N(_09777_),
    .B(_09778_),
    .X(_09779_));
 sky130_fd_sc_hd__xnor2_1 _16689_ (.A(_09771_),
    .B(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__a21oi_1 _16690_ (.A1(_09641_),
    .A2(_09650_),
    .B1(_09648_),
    .Y(_09781_));
 sky130_fd_sc_hd__nor2_1 _16691_ (.A(_09780_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__nand2_1 _16692_ (.A(_09780_),
    .B(_09781_),
    .Y(_09783_));
 sky130_fd_sc_hd__and2b_1 _16693_ (.A_N(_09782_),
    .B(_09783_),
    .X(_09784_));
 sky130_fd_sc_hd__xnor2_1 _16694_ (.A(_09770_),
    .B(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__a21o_1 _16695_ (.A1(_09759_),
    .A2(_09760_),
    .B1(_09785_),
    .X(_09786_));
 sky130_fd_sc_hd__nand3_1 _16696_ (.A(_09759_),
    .B(_09760_),
    .C(_09785_),
    .Y(_09787_));
 sky130_fd_sc_hd__nand2_1 _16697_ (.A(_09786_),
    .B(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__xnor2_2 _16698_ (.A(_09758_),
    .B(_09788_),
    .Y(_09789_));
 sky130_fd_sc_hd__a21o_1 _16699_ (.A1(_09670_),
    .A2(_09681_),
    .B1(_09679_),
    .X(_09790_));
 sky130_fd_sc_hd__nand2_1 _16700_ (.A(_09686_),
    .B(_09691_),
    .Y(_09791_));
 sky130_fd_sc_hd__a21bo_1 _16701_ (.A1(_09685_),
    .A2(_09692_),
    .B1_N(_09791_),
    .X(_09792_));
 sky130_fd_sc_hd__clkbuf_4 _16702_ (.A(_08422_),
    .X(_09793_));
 sky130_fd_sc_hd__or2_1 _16703_ (.A(_09158_),
    .B(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__or4_1 _16704_ (.A(_08545_),
    .B(_08602_),
    .C(_08407_),
    .D(_08349_),
    .X(_09795_));
 sky130_fd_sc_hd__inv_2 _16705_ (.A(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__o22a_1 _16706_ (.A1(_09417_),
    .A2(_08407_),
    .B1(_08349_),
    .B2(_08545_),
    .X(_09797_));
 sky130_fd_sc_hd__nor2_1 _16707_ (.A(_09796_),
    .B(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__xnor2_1 _16708_ (.A(_09794_),
    .B(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__a21o_1 _16709_ (.A1(_08395_),
    .A2(_09070_),
    .B1(_08587_),
    .X(_09800_));
 sky130_fd_sc_hd__nor3_1 _16710_ (.A(_08533_),
    .B(_09064_),
    .C(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__or2_1 _16711_ (.A(_08674_),
    .B(_09064_),
    .X(_09802_));
 sky130_fd_sc_hd__o21ai_1 _16712_ (.A1(_08533_),
    .A2(_09192_),
    .B1(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__and2b_1 _16713_ (.A_N(_09801_),
    .B(_09803_),
    .X(_09804_));
 sky130_fd_sc_hd__xnor2_1 _16714_ (.A(_09672_),
    .B(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__a22oi_1 _16715_ (.A1(_09533_),
    .A2(_09672_),
    .B1(_09674_),
    .B2(_09675_),
    .Y(_09806_));
 sky130_fd_sc_hd__nor2_1 _16716_ (.A(_09805_),
    .B(_09806_),
    .Y(_09807_));
 sky130_fd_sc_hd__and2_1 _16717_ (.A(_09805_),
    .B(_09806_),
    .X(_09808_));
 sky130_fd_sc_hd__nor2_1 _16718_ (.A(_09807_),
    .B(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__xnor2_1 _16719_ (.A(_09799_),
    .B(_09809_),
    .Y(_09810_));
 sky130_fd_sc_hd__xor2_1 _16720_ (.A(_09792_),
    .B(_09810_),
    .X(_09811_));
 sky130_fd_sc_hd__xnor2_2 _16721_ (.A(_09790_),
    .B(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__a21bo_1 _16722_ (.A1(_09552_),
    .A2(_09687_),
    .B1_N(_09689_),
    .X(_09813_));
 sky130_fd_sc_hd__o31a_1 _16723_ (.A1(_09700_),
    .A2(_09326_),
    .A3(_09699_),
    .B1(_09694_),
    .X(_09814_));
 sky130_fd_sc_hd__or2_1 _16724_ (.A(_08858_),
    .B(_09198_),
    .X(_09815_));
 sky130_fd_sc_hd__nor2_1 _16725_ (.A(_08868_),
    .B(_09696_),
    .Y(_09816_));
 sky130_fd_sc_hd__or2_1 _16726_ (.A(_08495_),
    .B(_09325_),
    .X(_09817_));
 sky130_fd_sc_hd__o21a_1 _16727_ (.A1(_08492_),
    .A2(_09695_),
    .B1(_09817_),
    .X(_09818_));
 sky130_fd_sc_hd__a21oi_1 _16728_ (.A1(_09701_),
    .A2(_09816_),
    .B1(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__xnor2_1 _16729_ (.A(_09815_),
    .B(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__xnor2_1 _16730_ (.A(_09814_),
    .B(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__xor2_2 _16731_ (.A(_09813_),
    .B(_09821_),
    .X(_09822_));
 sky130_fd_sc_hd__or2_1 _16732_ (.A(_09002_),
    .B(_09697_),
    .X(_09823_));
 sky130_fd_sc_hd__and2_1 _16733_ (.A(\rbzero.wall_tracer.stepDistX[8] ),
    .B(_06101_),
    .X(_09824_));
 sky130_fd_sc_hd__a21o_1 _16734_ (.A1(_08292_),
    .A2(_09572_),
    .B1(_09824_),
    .X(_09825_));
 sky130_fd_sc_hd__a21oi_2 _16735_ (.A1(_09703_),
    .A2(_09704_),
    .B1(_08977_),
    .Y(_09826_));
 sky130_fd_sc_hd__and3_1 _16736_ (.A(_08782_),
    .B(_09825_),
    .C(_09826_),
    .X(_09827_));
 sky130_fd_sc_hd__a21oi_1 _16737_ (.A1(_08782_),
    .A2(_09825_),
    .B1(_09826_),
    .Y(_09828_));
 sky130_fd_sc_hd__nor2_1 _16738_ (.A(_09827_),
    .B(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__xnor2_1 _16739_ (.A(_09823_),
    .B(_09829_),
    .Y(_09830_));
 sky130_fd_sc_hd__or4_1 _16740_ (.A(_08153_),
    .B(_08155_),
    .C(_08157_),
    .D(_09450_),
    .X(_09831_));
 sky130_fd_sc_hd__a21o_1 _16741_ (.A1(_08355_),
    .A2(_09831_),
    .B1(_08371_),
    .X(_09832_));
 sky130_fd_sc_hd__or3b_4 _16742_ (.A(_08390_),
    .B(_09832_),
    .C_N(_08164_),
    .X(_09833_));
 sky130_fd_sc_hd__mux2_1 _16743_ (.A0(\rbzero.wall_tracer.visualWallDist[10] ),
    .A1(_09755_),
    .S(_09833_),
    .X(_09834_));
 sky130_fd_sc_hd__nand2_1 _16744_ (.A(\rbzero.wall_tracer.stepDistY[9] ),
    .B(_09069_),
    .Y(_09835_));
 sky130_fd_sc_hd__a21oi_1 _16745_ (.A1(_09835_),
    .A2(_09711_),
    .B1(_08383_),
    .Y(_09836_));
 sky130_fd_sc_hd__xor2_1 _16746_ (.A(_09834_),
    .B(_09836_),
    .X(_09837_));
 sky130_fd_sc_hd__or2_1 _16747_ (.A(_09708_),
    .B(_09712_),
    .X(_09838_));
 sky130_fd_sc_hd__a21boi_1 _16748_ (.A1(_09707_),
    .A2(_09713_),
    .B1_N(_09838_),
    .Y(_09839_));
 sky130_fd_sc_hd__xor2_1 _16749_ (.A(_09837_),
    .B(_09839_),
    .X(_09840_));
 sky130_fd_sc_hd__xnor2_1 _16750_ (.A(_09830_),
    .B(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__and2b_1 _16751_ (.A_N(_09714_),
    .B(_09715_),
    .X(_09842_));
 sky130_fd_sc_hd__a21o_1 _16752_ (.A1(_09702_),
    .A2(_09716_),
    .B1(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__xnor2_1 _16753_ (.A(_09841_),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__xnor2_2 _16754_ (.A(_09822_),
    .B(_09844_),
    .Y(_09845_));
 sky130_fd_sc_hd__nor2_1 _16755_ (.A(_09717_),
    .B(_09718_),
    .Y(_09846_));
 sky130_fd_sc_hd__a21o_1 _16756_ (.A1(_09693_),
    .A2(_09719_),
    .B1(_09846_),
    .X(_09847_));
 sky130_fd_sc_hd__xnor2_1 _16757_ (.A(_09845_),
    .B(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__xnor2_2 _16758_ (.A(_09812_),
    .B(_09848_),
    .Y(_09849_));
 sky130_fd_sc_hd__a21o_1 _16759_ (.A1(_09684_),
    .A2(_09723_),
    .B1(_09722_),
    .X(_09850_));
 sky130_fd_sc_hd__xnor2_2 _16760_ (.A(_09849_),
    .B(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__xnor2_2 _16761_ (.A(_09789_),
    .B(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__a21oi_1 _16762_ (.A1(_09660_),
    .A2(_09728_),
    .B1(_09726_),
    .Y(_09853_));
 sky130_fd_sc_hd__xor2_2 _16763_ (.A(_09852_),
    .B(_09853_),
    .X(_09854_));
 sky130_fd_sc_hd__xnor2_4 _16764_ (.A(_09757_),
    .B(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__a21oi_4 _16765_ (.A1(_09627_),
    .A2(_09732_),
    .B1(_09730_),
    .Y(_09856_));
 sky130_fd_sc_hd__xnor2_4 _16766_ (.A(_09855_),
    .B(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__xor2_4 _16767_ (.A(_09749_),
    .B(_09857_),
    .X(_09858_));
 sky130_fd_sc_hd__xnor2_4 _16768_ (.A(_09748_),
    .B(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__mux2_1 _16769_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_08263_),
    .X(_09860_));
 sky130_fd_sc_hd__xnor2_1 _16770_ (.A(_09268_),
    .B(_09860_),
    .Y(_09861_));
 sky130_fd_sc_hd__xnor2_1 _16771_ (.A(_09859_),
    .B(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__xnor2_2 _16772_ (.A(_09747_),
    .B(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__or2_1 _16773_ (.A(\rbzero.texu_hot[5] ),
    .B(_08270_),
    .X(_09864_));
 sky130_fd_sc_hd__o211a_1 _16774_ (.A1(_08355_),
    .A2(_09863_),
    .B1(_09864_),
    .C1(_08211_),
    .X(_00471_));
 sky130_fd_sc_hd__nor2_1 _16775_ (.A(_04549_),
    .B(_04869_),
    .Y(_09865_));
 sky130_fd_sc_hd__and4_1 _16776_ (.A(_04186_),
    .B(_04770_),
    .C(_05200_),
    .D(_09865_),
    .X(_09866_));
 sky130_fd_sc_hd__buf_4 _16777_ (.A(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__or2_1 _16778_ (.A(_04544_),
    .B(_09867_),
    .X(_09868_));
 sky130_fd_sc_hd__clkbuf_2 _16779_ (.A(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__nor2_1 _16780_ (.A(_04105_),
    .B(_09869_),
    .Y(_00472_));
 sky130_fd_sc_hd__nor2_8 _16781_ (.A(_04544_),
    .B(_09867_),
    .Y(_09870_));
 sky130_fd_sc_hd__and3_1 _16782_ (.A(_04580_),
    .B(_04581_),
    .C(_09870_),
    .X(_09871_));
 sky130_fd_sc_hd__clkbuf_1 _16783_ (.A(_09871_),
    .X(_00473_));
 sky130_fd_sc_hd__or2_1 _16784_ (.A(_04544_),
    .B(_04769_),
    .X(_09872_));
 sky130_fd_sc_hd__a21oi_1 _16785_ (.A1(_04579_),
    .A2(_04580_),
    .B1(_09872_),
    .Y(_00474_));
 sky130_fd_sc_hd__nor2_1 _16786_ (.A(net64),
    .B(_05188_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _16787_ (.A(_05207_),
    .B(_09869_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _16788_ (.A(_05212_),
    .B(_09869_),
    .Y(_00477_));
 sky130_fd_sc_hd__and2_1 _16789_ (.A(_05186_),
    .B(_09870_),
    .X(_09873_));
 sky130_fd_sc_hd__clkbuf_1 _16790_ (.A(_09873_),
    .X(_00478_));
 sky130_fd_sc_hd__nor2_1 _16791_ (.A(_05223_),
    .B(_09869_),
    .Y(_00479_));
 sky130_fd_sc_hd__and4_1 _16792_ (.A(_04110_),
    .B(_04550_),
    .C(_04769_),
    .D(_05392_),
    .X(_09874_));
 sky130_fd_sc_hd__a31o_1 _16793_ (.A1(_04550_),
    .A2(_04769_),
    .A3(_05392_),
    .B1(_04110_),
    .X(_09875_));
 sky130_fd_sc_hd__and3b_1 _16794_ (.A_N(_09874_),
    .B(_09875_),
    .C(_09870_),
    .X(_09876_));
 sky130_fd_sc_hd__clkbuf_1 _16795_ (.A(_09876_),
    .X(_00480_));
 sky130_fd_sc_hd__a21oi_1 _16796_ (.A1(_04111_),
    .A2(_09874_),
    .B1(_09869_),
    .Y(_09877_));
 sky130_fd_sc_hd__o21a_1 _16797_ (.A1(_04111_),
    .A2(_09874_),
    .B1(_09877_),
    .X(_00481_));
 sky130_fd_sc_hd__and3_1 _16798_ (.A(\rbzero.trace_state[0] ),
    .B(_05173_),
    .C(_09867_),
    .X(_09878_));
 sky130_fd_sc_hd__nor2_1 _16799_ (.A(_04566_),
    .B(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__clkbuf_4 _16800_ (.A(_09879_),
    .X(_09880_));
 sky130_fd_sc_hd__buf_4 _16801_ (.A(_09880_),
    .X(_09881_));
 sky130_fd_sc_hd__buf_4 _16802_ (.A(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__and4_1 _16803_ (.A(_04571_),
    .B(_04567_),
    .C(_05173_),
    .D(_09867_),
    .X(_09883_));
 sky130_fd_sc_hd__buf_6 _16804_ (.A(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__buf_4 _16805_ (.A(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__a22o_1 _16806_ (.A1(\rbzero.row_render.side ),
    .A2(_09882_),
    .B1(_09885_),
    .B2(_08263_),
    .X(_00482_));
 sky130_fd_sc_hd__a22o_1 _16807_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_09882_),
    .B1(_09885_),
    .B2(_08050_),
    .X(_00483_));
 sky130_fd_sc_hd__a22o_1 _16808_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_09882_),
    .B1(_09885_),
    .B2(_08064_),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _16809_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_09882_),
    .B1(_09885_),
    .B2(_08074_),
    .X(_00485_));
 sky130_fd_sc_hd__a22o_1 _16810_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_09882_),
    .B1(_09885_),
    .B2(_08085_),
    .X(_00486_));
 sky130_fd_sc_hd__a22o_1 _16811_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_09882_),
    .B1(_09885_),
    .B2(_08094_),
    .X(_00487_));
 sky130_fd_sc_hd__a22o_1 _16812_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_09882_),
    .B1(_09885_),
    .B2(_08100_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_4 _16813_ (.A(_09880_),
    .X(_09886_));
 sky130_fd_sc_hd__buf_4 _16814_ (.A(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__a22o_1 _16815_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_09887_),
    .B1(_09885_),
    .B2(_08104_),
    .X(_00489_));
 sky130_fd_sc_hd__buf_4 _16816_ (.A(_09884_),
    .X(_09888_));
 sky130_fd_sc_hd__buf_4 _16817_ (.A(_09888_),
    .X(_09889_));
 sky130_fd_sc_hd__a22o_1 _16818_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(_08111_),
    .X(_00490_));
 sky130_fd_sc_hd__a22o_1 _16819_ (.A1(\rbzero.row_render.size[8] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(_08117_),
    .X(_00491_));
 sky130_fd_sc_hd__a22o_1 _16820_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(_08121_),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _16821_ (.A1(\rbzero.row_render.size[10] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(_08126_),
    .X(_00493_));
 sky130_fd_sc_hd__a22o_1 _16822_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(\rbzero.texu_hot[0] ),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _16823_ (.A1(\rbzero.row_render.texu[1] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(\rbzero.texu_hot[1] ),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _16824_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(\rbzero.texu_hot[2] ),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_1 _16825_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(\rbzero.texu_hot[3] ),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _16826_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_09887_),
    .B1(_09889_),
    .B2(\rbzero.texu_hot[4] ),
    .X(_00498_));
 sky130_fd_sc_hd__clkbuf_4 _16827_ (.A(_09886_),
    .X(_09890_));
 sky130_fd_sc_hd__a22o_1 _16828_ (.A1(\rbzero.traced_texa[-11] ),
    .A2(_09890_),
    .B1(_09889_),
    .B2(_08164_),
    .X(_00499_));
 sky130_fd_sc_hd__clkbuf_4 _16829_ (.A(_09888_),
    .X(_09891_));
 sky130_fd_sc_hd__a22o_1 _16830_ (.A1(\rbzero.traced_texa[-10] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _16831_ (.A1(\rbzero.traced_texa[-9] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_1 _16832_ (.A1(\rbzero.traced_texa[-8] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(net518),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _16833_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _16834_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _16835_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _16836_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(_00506_));
 sky130_fd_sc_hd__a22o_1 _16837_ (.A1(\rbzero.traced_texa[-3] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _16838_ (.A1(\rbzero.traced_texa[-2] ),
    .A2(_09890_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_00508_));
 sky130_fd_sc_hd__clkbuf_4 _16839_ (.A(_09881_),
    .X(_09892_));
 sky130_fd_sc_hd__a22o_1 _16840_ (.A1(\rbzero.traced_texa[-1] ),
    .A2(_09892_),
    .B1(_09891_),
    .B2(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_00509_));
 sky130_fd_sc_hd__buf_2 _16841_ (.A(_09884_),
    .X(_09893_));
 sky130_fd_sc_hd__a22o_1 _16842_ (.A1(\rbzero.traced_texa[0] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_00510_));
 sky130_fd_sc_hd__a22o_1 _16843_ (.A1(\rbzero.traced_texa[1] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_00511_));
 sky130_fd_sc_hd__a22o_1 _16844_ (.A1(\rbzero.traced_texa[2] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _16845_ (.A1(\rbzero.traced_texa[3] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(_00513_));
 sky130_fd_sc_hd__a22o_1 _16846_ (.A1(\rbzero.traced_texa[4] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_1 _16847_ (.A1(\rbzero.traced_texa[5] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _16848_ (.A1(\rbzero.traced_texa[6] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_00516_));
 sky130_fd_sc_hd__a22o_1 _16849_ (.A1(\rbzero.traced_texa[7] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _16850_ (.A1(\rbzero.traced_texa[8] ),
    .A2(_09892_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_00518_));
 sky130_fd_sc_hd__buf_4 _16851_ (.A(_09881_),
    .X(_09894_));
 sky130_fd_sc_hd__a22o_1 _16852_ (.A1(\rbzero.traced_texa[9] ),
    .A2(_09894_),
    .B1(_09893_),
    .B2(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_00519_));
 sky130_fd_sc_hd__buf_2 _16853_ (.A(_09884_),
    .X(_09895_));
 sky130_fd_sc_hd__a22o_1 _16854_ (.A1(\rbzero.traced_texa[10] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _16855_ (.A0(\rbzero.row_render.wall[0] ),
    .A1(_04592_),
    .S(_09884_),
    .X(_09896_));
 sky130_fd_sc_hd__clkbuf_1 _16856_ (.A(_09896_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _16857_ (.A0(\rbzero.row_render.wall[1] ),
    .A1(\rbzero.wall_hot[1] ),
    .S(_09884_),
    .X(_09897_));
 sky130_fd_sc_hd__clkbuf_1 _16858_ (.A(_09897_),
    .X(_00522_));
 sky130_fd_sc_hd__o21a_1 _16859_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(\rbzero.wall_tracer.mapX[5] ),
    .B1(_09265_),
    .X(_09898_));
 sky130_fd_sc_hd__xor2_1 _16860_ (.A(\rbzero.wall_tracer.mapX[5] ),
    .B(_09265_),
    .X(_09899_));
 sky130_fd_sc_hd__xnor2_1 _16861_ (.A(_06186_),
    .B(_09265_),
    .Y(_09900_));
 sky130_fd_sc_hd__or2_1 _16862_ (.A(_06223_),
    .B(_09265_),
    .X(_09901_));
 sky130_fd_sc_hd__and2_1 _16863_ (.A(\rbzero.map_rom.f3 ),
    .B(_08334_),
    .X(_09902_));
 sky130_fd_sc_hd__nor2_1 _16864_ (.A(\rbzero.map_rom.f3 ),
    .B(_08334_),
    .Y(_09903_));
 sky130_fd_sc_hd__nor2_1 _16865_ (.A(_09902_),
    .B(_09903_),
    .Y(_09904_));
 sky130_fd_sc_hd__and2_1 _16866_ (.A(\rbzero.map_rom.f4 ),
    .B(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__xnor2_1 _16867_ (.A(_06200_),
    .B(_08334_),
    .Y(_09906_));
 sky130_fd_sc_hd__o21ai_1 _16868_ (.A1(_09902_),
    .A2(_09905_),
    .B1(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__a21bo_1 _16869_ (.A1(_06184_),
    .A2(_09265_),
    .B1_N(_09907_),
    .X(_09908_));
 sky130_fd_sc_hd__nand2_1 _16870_ (.A(_06223_),
    .B(_09265_),
    .Y(_09909_));
 sky130_fd_sc_hd__or2b_1 _16871_ (.A(_09908_),
    .B_N(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__and3_1 _16872_ (.A(_09900_),
    .B(_09901_),
    .C(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__and2_1 _16873_ (.A(_09899_),
    .B(_09911_),
    .X(_09912_));
 sky130_fd_sc_hd__xor2_1 _16874_ (.A(\rbzero.wall_tracer.mapX[6] ),
    .B(_09265_),
    .X(_09913_));
 sky130_fd_sc_hd__o21a_1 _16875_ (.A1(_09898_),
    .A2(_09912_),
    .B1(_09913_),
    .X(_09914_));
 sky130_fd_sc_hd__buf_6 _16876_ (.A(_06180_),
    .X(_09915_));
 sky130_fd_sc_hd__a211o_4 _16877_ (.A1(_06180_),
    .A2(_08292_),
    .B1(_06283_),
    .C1(_08264_),
    .X(_09916_));
 sky130_fd_sc_hd__nor2_2 _16878_ (.A(_09915_),
    .B(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__o31ai_1 _16879_ (.A1(_09913_),
    .A2(_09898_),
    .A3(_09912_),
    .B1(_09917_),
    .Y(_09918_));
 sky130_fd_sc_hd__buf_6 _16880_ (.A(_09916_),
    .X(_09919_));
 sky130_fd_sc_hd__buf_4 _16881_ (.A(_09919_),
    .X(_09920_));
 sky130_fd_sc_hd__a2bb2o_1 _16882_ (.A1_N(_09914_),
    .A2_N(_09918_),
    .B1(\rbzero.wall_tracer.mapX[6] ),
    .B2(_09920_),
    .X(_00523_));
 sky130_fd_sc_hd__xor2_1 _16883_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(_09265_),
    .X(_09921_));
 sky130_fd_sc_hd__a21o_1 _16884_ (.A1(\rbzero.wall_tracer.mapX[6] ),
    .A2(_09266_),
    .B1(_09914_),
    .X(_09922_));
 sky130_fd_sc_hd__xor2_1 _16885_ (.A(_09921_),
    .B(_09922_),
    .X(_09923_));
 sky130_fd_sc_hd__a22o_1 _16886_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(_09920_),
    .B1(_09917_),
    .B2(_09923_),
    .X(_00524_));
 sky130_fd_sc_hd__xor2_1 _16887_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(_09266_),
    .X(_09924_));
 sky130_fd_sc_hd__and3_1 _16888_ (.A(_09913_),
    .B(_09912_),
    .C(_09921_),
    .X(_09925_));
 sky130_fd_sc_hd__o21a_1 _16889_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(\rbzero.wall_tracer.mapX[6] ),
    .B1(_09265_),
    .X(_09926_));
 sky130_fd_sc_hd__or3_1 _16890_ (.A(_09898_),
    .B(_09925_),
    .C(_09926_),
    .X(_09927_));
 sky130_fd_sc_hd__xor2_1 _16891_ (.A(_09924_),
    .B(_09927_),
    .X(_09928_));
 sky130_fd_sc_hd__a22o_1 _16892_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09920_),
    .B1(_09917_),
    .B2(_09928_),
    .X(_00525_));
 sky130_fd_sc_hd__a22o_1 _16893_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09266_),
    .B1(_09924_),
    .B2(_09927_),
    .X(_09929_));
 sky130_fd_sc_hd__xnor2_1 _16894_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(_09266_),
    .Y(_09930_));
 sky130_fd_sc_hd__xnor2_1 _16895_ (.A(_09929_),
    .B(_09930_),
    .Y(_09931_));
 sky130_fd_sc_hd__a22o_1 _16896_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09920_),
    .B1(_09917_),
    .B2(_09931_),
    .X(_00526_));
 sky130_fd_sc_hd__o21a_1 _16897_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09266_),
    .B1(_09929_),
    .X(_09932_));
 sky130_fd_sc_hd__a21oi_1 _16898_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09266_),
    .B1(_09932_),
    .Y(_09933_));
 sky130_fd_sc_hd__xnor2_1 _16899_ (.A(\rbzero.wall_tracer.mapX[10] ),
    .B(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__nand2_1 _16900_ (.A(_09266_),
    .B(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__or2_1 _16901_ (.A(_09266_),
    .B(_09934_),
    .X(_09936_));
 sky130_fd_sc_hd__a32o_1 _16902_ (.A1(_09917_),
    .A2(_09935_),
    .A3(_09936_),
    .B1(_09919_),
    .B2(\rbzero.wall_tracer.mapX[10] ),
    .X(_00527_));
 sky130_fd_sc_hd__buf_12 _16903_ (.A(_06095_),
    .X(_09937_));
 sky130_fd_sc_hd__clkbuf_16 _16904_ (.A(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__a21oi_1 _16905_ (.A1(_08989_),
    .A2(_09037_),
    .B1(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__o21ai_1 _16906_ (.A1(_08989_),
    .A2(_09037_),
    .B1(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__o21ai_1 _16907_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09937_),
    .Y(_09941_));
 sky130_fd_sc_hd__a21oi_1 _16908_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09941_),
    .Y(_09942_));
 sky130_fd_sc_hd__nor2_1 _16909_ (.A(_09919_),
    .B(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__inv_2 _16910_ (.A(_09916_),
    .Y(_09944_));
 sky130_fd_sc_hd__buf_4 _16911_ (.A(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__buf_4 _16912_ (.A(_09945_),
    .X(_09946_));
 sky130_fd_sc_hd__o2bb2a_1 _16913_ (.A1_N(_09940_),
    .A2_N(_09943_),
    .B1(\rbzero.wall_tracer.trackDistX[-11] ),
    .B2(_09946_),
    .X(_00528_));
 sky130_fd_sc_hd__xnor2_1 _16914_ (.A(_09039_),
    .B(_09041_),
    .Y(_09947_));
 sky130_fd_sc_hd__or2_1 _16915_ (.A(_09938_),
    .B(_09947_),
    .X(_09948_));
 sky130_fd_sc_hd__or2_1 _16916_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_09949_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_09950_));
 sky130_fd_sc_hd__and4_1 _16918_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .C(_09949_),
    .D(_09950_),
    .X(_09951_));
 sky130_fd_sc_hd__a22oi_1 _16919_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09949_),
    .B2(_09950_),
    .Y(_09952_));
 sky130_fd_sc_hd__o31a_1 _16920_ (.A1(_06288_),
    .A2(_09951_),
    .A3(_09952_),
    .B1(_09945_),
    .X(_09953_));
 sky130_fd_sc_hd__o2bb2a_1 _16921_ (.A1_N(_09948_),
    .A2_N(_09953_),
    .B1(\rbzero.wall_tracer.trackDistX[-10] ),
    .B2(_09946_),
    .X(_00529_));
 sky130_fd_sc_hd__buf_4 _16922_ (.A(_06287_),
    .X(_09954_));
 sky130_fd_sc_hd__a21oi_1 _16923_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(\rbzero.wall_tracer.stepDistX[-10] ),
    .B1(_09951_),
    .Y(_09955_));
 sky130_fd_sc_hd__nor2_1 _16924_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .Y(_09956_));
 sky130_fd_sc_hd__and2_1 _16925_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_09957_));
 sky130_fd_sc_hd__nor3_1 _16926_ (.A(_09955_),
    .B(_09956_),
    .C(_09957_),
    .Y(_09958_));
 sky130_fd_sc_hd__o21a_1 _16927_ (.A1(_09956_),
    .A2(_09957_),
    .B1(_09955_),
    .X(_09959_));
 sky130_fd_sc_hd__nand2_1 _16928_ (.A(_09915_),
    .B(_09258_),
    .Y(_09960_));
 sky130_fd_sc_hd__o311a_1 _16929_ (.A1(_09954_),
    .A2(_09958_),
    .A3(_09959_),
    .B1(_09945_),
    .C1(_09960_),
    .X(_09961_));
 sky130_fd_sc_hd__a21oi_1 _16930_ (.A1(_06138_),
    .A2(_09920_),
    .B1(_09961_),
    .Y(_00530_));
 sky130_fd_sc_hd__or2_1 _16931_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_09962_));
 sky130_fd_sc_hd__nand2_1 _16932_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_09963_));
 sky130_fd_sc_hd__o21bai_1 _16933_ (.A1(_09955_),
    .A2(_09956_),
    .B1_N(_09957_),
    .Y(_09964_));
 sky130_fd_sc_hd__and3_1 _16934_ (.A(_09962_),
    .B(_09963_),
    .C(_09964_),
    .X(_09965_));
 sky130_fd_sc_hd__a21oi_1 _16935_ (.A1(_09962_),
    .A2(_09963_),
    .B1(_09964_),
    .Y(_09966_));
 sky130_fd_sc_hd__nand2_1 _16936_ (.A(_09915_),
    .B(_09257_),
    .Y(_09967_));
 sky130_fd_sc_hd__o311a_1 _16937_ (.A1(_09954_),
    .A2(_09965_),
    .A3(_09966_),
    .B1(_09945_),
    .C1(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__a21oi_1 _16938_ (.A1(_06153_),
    .A2(_09920_),
    .B1(_09968_),
    .Y(_00531_));
 sky130_fd_sc_hd__nor2_1 _16939_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09969_));
 sky130_fd_sc_hd__nand2_1 _16940_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09970_));
 sky130_fd_sc_hd__or2b_1 _16941_ (.A(_09969_),
    .B_N(_09970_),
    .X(_09971_));
 sky130_fd_sc_hd__a21boi_1 _16942_ (.A1(_09962_),
    .A2(_09964_),
    .B1_N(_09963_),
    .Y(_09972_));
 sky130_fd_sc_hd__nor2_1 _16943_ (.A(_09971_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__buf_4 _16944_ (.A(_06180_),
    .X(_09974_));
 sky130_fd_sc_hd__a21o_1 _16945_ (.A1(_09971_),
    .A2(_09972_),
    .B1(_09974_),
    .X(_09975_));
 sky130_fd_sc_hd__nand2_1 _16946_ (.A(_06287_),
    .B(_09253_),
    .Y(_09976_));
 sky130_fd_sc_hd__o21ai_1 _16947_ (.A1(_09973_),
    .A2(_09975_),
    .B1(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__buf_6 _16948_ (.A(_09944_),
    .X(_09978_));
 sky130_fd_sc_hd__mux2_1 _16949_ (.A0(\rbzero.wall_tracer.trackDistX[-7] ),
    .A1(_09977_),
    .S(_09978_),
    .X(_09979_));
 sky130_fd_sc_hd__clkbuf_1 _16950_ (.A(_09979_),
    .X(_00532_));
 sky130_fd_sc_hd__or2_1 _16951_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_09980_));
 sky130_fd_sc_hd__nand2_1 _16952_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_09981_));
 sky130_fd_sc_hd__o21ai_1 _16953_ (.A1(_09969_),
    .A2(_09972_),
    .B1(_09970_),
    .Y(_09982_));
 sky130_fd_sc_hd__and3_1 _16954_ (.A(_09980_),
    .B(_09981_),
    .C(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__a21oi_1 _16955_ (.A1(_09980_),
    .A2(_09981_),
    .B1(_09982_),
    .Y(_09984_));
 sky130_fd_sc_hd__nand2_1 _16956_ (.A(_09915_),
    .B(_09249_),
    .Y(_09985_));
 sky130_fd_sc_hd__o311a_1 _16957_ (.A1(_09954_),
    .A2(_09983_),
    .A3(_09984_),
    .B1(_09945_),
    .C1(_09985_),
    .X(_09986_));
 sky130_fd_sc_hd__a21oi_1 _16958_ (.A1(_06124_),
    .A2(_09920_),
    .B1(_09986_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_1 _16959_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_1 _16960_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09988_));
 sky130_fd_sc_hd__or2b_1 _16961_ (.A(_09987_),
    .B_N(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__a21boi_1 _16962_ (.A1(_09980_),
    .A2(_09982_),
    .B1_N(_09981_),
    .Y(_09990_));
 sky130_fd_sc_hd__nor2_1 _16963_ (.A(_09989_),
    .B(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__a21o_1 _16964_ (.A1(_09989_),
    .A2(_09990_),
    .B1(_09974_),
    .X(_09992_));
 sky130_fd_sc_hd__nand2_1 _16965_ (.A(_06287_),
    .B(_09366_),
    .Y(_09993_));
 sky130_fd_sc_hd__o21ai_1 _16966_ (.A1(_09991_),
    .A2(_09992_),
    .B1(_09993_),
    .Y(_09994_));
 sky130_fd_sc_hd__mux2_1 _16967_ (.A0(\rbzero.wall_tracer.trackDistX[-5] ),
    .A1(_09994_),
    .S(_09978_),
    .X(_09995_));
 sky130_fd_sc_hd__clkbuf_1 _16968_ (.A(_09995_),
    .X(_00534_));
 sky130_fd_sc_hd__or2_1 _16969_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(_09996_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09997_));
 sky130_fd_sc_hd__o21ai_1 _16971_ (.A1(_09987_),
    .A2(_09990_),
    .B1(_09988_),
    .Y(_09998_));
 sky130_fd_sc_hd__and3_1 _16972_ (.A(_09996_),
    .B(_09997_),
    .C(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__a21oi_1 _16973_ (.A1(_09996_),
    .A2(_09997_),
    .B1(_09998_),
    .Y(_10000_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(_09915_),
    .B(_09487_),
    .Y(_10001_));
 sky130_fd_sc_hd__o311a_1 _16975_ (.A1(_09954_),
    .A2(_09999_),
    .A3(_10000_),
    .B1(_09945_),
    .C1(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__a21oi_1 _16976_ (.A1(_06129_),
    .A2(_09920_),
    .B1(_10002_),
    .Y(_00535_));
 sky130_fd_sc_hd__nor2_1 _16977_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_10003_));
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_10004_));
 sky130_fd_sc_hd__or2b_1 _16979_ (.A(_10003_),
    .B_N(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__a21boi_1 _16980_ (.A1(_09996_),
    .A2(_09998_),
    .B1_N(_09997_),
    .Y(_10006_));
 sky130_fd_sc_hd__nor2_1 _16981_ (.A(_10005_),
    .B(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__a21o_1 _16982_ (.A1(_10005_),
    .A2(_10006_),
    .B1(_09974_),
    .X(_10008_));
 sky130_fd_sc_hd__xnor2_4 _16983_ (.A(_09496_),
    .B(_09610_),
    .Y(_10009_));
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(_06287_),
    .B(_10009_),
    .Y(_10010_));
 sky130_fd_sc_hd__o21ai_1 _16985_ (.A1(_10007_),
    .A2(_10008_),
    .B1(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__mux2_1 _16986_ (.A0(\rbzero.wall_tracer.trackDistX[-3] ),
    .A1(_10011_),
    .S(_09978_),
    .X(_10012_));
 sky130_fd_sc_hd__clkbuf_1 _16987_ (.A(_10012_),
    .X(_00536_));
 sky130_fd_sc_hd__or2_1 _16988_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_10013_));
 sky130_fd_sc_hd__nand2_1 _16989_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_10014_));
 sky130_fd_sc_hd__o21ai_1 _16990_ (.A1(_10003_),
    .A2(_10006_),
    .B1(_10004_),
    .Y(_10015_));
 sky130_fd_sc_hd__and3_1 _16991_ (.A(_10013_),
    .B(_10014_),
    .C(_10015_),
    .X(_10016_));
 sky130_fd_sc_hd__a21oi_1 _16992_ (.A1(_10013_),
    .A2(_10014_),
    .B1(_10015_),
    .Y(_10017_));
 sky130_fd_sc_hd__nand2_1 _16993_ (.A(_09915_),
    .B(_09738_),
    .Y(_10018_));
 sky130_fd_sc_hd__o311a_1 _16994_ (.A1(_09954_),
    .A2(_10016_),
    .A3(_10017_),
    .B1(_09978_),
    .C1(_10018_),
    .X(_10019_));
 sky130_fd_sc_hd__a21oi_1 _16995_ (.A1(_06113_),
    .A2(_09920_),
    .B1(_10019_),
    .Y(_00537_));
 sky130_fd_sc_hd__nor2_1 _16996_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_10020_));
 sky130_fd_sc_hd__and2_1 _16997_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(_10021_));
 sky130_fd_sc_hd__or2_1 _16998_ (.A(_10020_),
    .B(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__a21boi_1 _16999_ (.A1(_10013_),
    .A2(_10015_),
    .B1_N(_10014_),
    .Y(_10023_));
 sky130_fd_sc_hd__nor2_1 _17000_ (.A(_10022_),
    .B(_10023_),
    .Y(_10024_));
 sky130_fd_sc_hd__a21o_1 _17001_ (.A1(_10022_),
    .A2(_10023_),
    .B1(_09974_),
    .X(_10025_));
 sky130_fd_sc_hd__nand2_1 _17002_ (.A(_06287_),
    .B(_09859_),
    .Y(_10026_));
 sky130_fd_sc_hd__o21ai_1 _17003_ (.A1(_10024_),
    .A2(_10025_),
    .B1(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__mux2_1 _17004_ (.A0(\rbzero.wall_tracer.trackDistX[-1] ),
    .A1(_10027_),
    .S(_09978_),
    .X(_10028_));
 sky130_fd_sc_hd__clkbuf_1 _17005_ (.A(_10028_),
    .X(_00538_));
 sky130_fd_sc_hd__nor2_4 _17006_ (.A(_09855_),
    .B(_09856_),
    .Y(_10029_));
 sky130_fd_sc_hd__nor2_4 _17007_ (.A(_08217_),
    .B(_08390_),
    .Y(_10030_));
 sky130_fd_sc_hd__a31o_1 _17008_ (.A1(_08550_),
    .A2(_09754_),
    .A3(_10030_),
    .B1(_09752_),
    .X(_10031_));
 sky130_fd_sc_hd__or2b_1 _17009_ (.A(_09788_),
    .B_N(_09758_),
    .X(_10032_));
 sky130_fd_sc_hd__o2bb2a_1 _17010_ (.A1_N(_09767_),
    .A2_N(_09769_),
    .B1(_09764_),
    .B2(_09766_),
    .X(_10033_));
 sky130_fd_sc_hd__a21oi_4 _17011_ (.A1(_09786_),
    .A2(_10032_),
    .B1(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__and3_1 _17012_ (.A(_09786_),
    .B(_10032_),
    .C(_10033_),
    .X(_10035_));
 sky130_fd_sc_hd__nor2_1 _17013_ (.A(_10034_),
    .B(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__a21o_1 _17014_ (.A1(_09770_),
    .A2(_09783_),
    .B1(_09782_),
    .X(_10037_));
 sky130_fd_sc_hd__or2b_1 _17015_ (.A(_09810_),
    .B_N(_09792_),
    .X(_10038_));
 sky130_fd_sc_hd__or2b_1 _17016_ (.A(_09811_),
    .B_N(_09790_),
    .X(_10039_));
 sky130_fd_sc_hd__nor2_1 _17017_ (.A(_09157_),
    .B(_09502_),
    .Y(_10040_));
 sky130_fd_sc_hd__xnor2_1 _17018_ (.A(_09761_),
    .B(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__or2_1 _17019_ (.A(_09135_),
    .B(_09636_),
    .X(_10042_));
 sky130_fd_sc_hd__xnor2_1 _17020_ (.A(_10041_),
    .B(_10042_),
    .Y(_10043_));
 sky130_fd_sc_hd__nand2_1 _17021_ (.A(_09642_),
    .B(_09761_),
    .Y(_10044_));
 sky130_fd_sc_hd__o31a_1 _17022_ (.A1(_09135_),
    .A2(_09503_),
    .A3(_09762_),
    .B1(_10044_),
    .X(_10045_));
 sky130_fd_sc_hd__nor2_1 _17023_ (.A(_10043_),
    .B(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__and2_1 _17024_ (.A(_10043_),
    .B(_10045_),
    .X(_10047_));
 sky130_fd_sc_hd__nor2_1 _17025_ (.A(_10046_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__or2_1 _17026_ (.A(_08553_),
    .B(_09755_),
    .X(_10049_));
 sky130_fd_sc_hd__xnor2_1 _17027_ (.A(_10048_),
    .B(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__or2b_1 _17028_ (.A(_09644_),
    .B_N(_09775_),
    .X(_10051_));
 sky130_fd_sc_hd__o31ai_2 _17029_ (.A1(_09406_),
    .A2(_09162_),
    .A3(_09773_),
    .B1(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__o21ai_1 _17030_ (.A1(_09794_),
    .A2(_09797_),
    .B1(_09795_),
    .Y(_10053_));
 sky130_fd_sc_hd__o21ai_1 _17031_ (.A1(_08829_),
    .A2(_09225_),
    .B1(_09773_),
    .Y(_10054_));
 sky130_fd_sc_hd__or3_1 _17032_ (.A(_08829_),
    .B(_09222_),
    .C(_09773_),
    .X(_10055_));
 sky130_fd_sc_hd__nand2_1 _17033_ (.A(_10054_),
    .B(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__nor2_1 _17034_ (.A(_09404_),
    .B(_09276_),
    .Y(_10057_));
 sky130_fd_sc_hd__xnor2_1 _17035_ (.A(_10056_),
    .B(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__and2_1 _17036_ (.A(_10053_),
    .B(_10058_),
    .X(_10059_));
 sky130_fd_sc_hd__nor2_1 _17037_ (.A(_10053_),
    .B(_10058_),
    .Y(_10060_));
 sky130_fd_sc_hd__nor2_1 _17038_ (.A(_10059_),
    .B(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__xnor2_1 _17039_ (.A(_10052_),
    .B(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__a21oi_1 _17040_ (.A1(_09771_),
    .A2(_09779_),
    .B1(_09777_),
    .Y(_10063_));
 sky130_fd_sc_hd__nor2_1 _17041_ (.A(_10062_),
    .B(_10063_),
    .Y(_10064_));
 sky130_fd_sc_hd__and2_1 _17042_ (.A(_10062_),
    .B(_10063_),
    .X(_10065_));
 sky130_fd_sc_hd__nor2_1 _17043_ (.A(_10064_),
    .B(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__xnor2_1 _17044_ (.A(_10050_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__a21o_1 _17045_ (.A1(_10038_),
    .A2(_10039_),
    .B1(_10067_),
    .X(_10068_));
 sky130_fd_sc_hd__nand3_1 _17046_ (.A(_10038_),
    .B(_10039_),
    .C(_10067_),
    .Y(_10069_));
 sky130_fd_sc_hd__nand2_1 _17047_ (.A(_10068_),
    .B(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__xnor2_1 _17048_ (.A(_10037_),
    .B(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__a21o_1 _17049_ (.A1(_09799_),
    .A2(_09809_),
    .B1(_09807_),
    .X(_10072_));
 sky130_fd_sc_hd__and2b_1 _17050_ (.A_N(_09814_),
    .B(_09820_),
    .X(_10073_));
 sky130_fd_sc_hd__a21o_1 _17051_ (.A1(_09813_),
    .A2(_09821_),
    .B1(_10073_),
    .X(_10074_));
 sky130_fd_sc_hd__buf_2 _17052_ (.A(_08509_),
    .X(_10075_));
 sky130_fd_sc_hd__o22ai_1 _17053_ (.A1(_08545_),
    .A2(_10075_),
    .B1(_08349_),
    .B2(_09158_),
    .Y(_10076_));
 sky130_fd_sc_hd__or4_1 _17054_ (.A(_08544_),
    .B(_09158_),
    .C(_08509_),
    .D(_08349_),
    .X(_10077_));
 sky130_fd_sc_hd__nand2_1 _17055_ (.A(_10076_),
    .B(_10077_),
    .Y(_10078_));
 sky130_fd_sc_hd__or3_1 _17056_ (.A(_09793_),
    .B(_09162_),
    .C(_10078_),
    .X(_10079_));
 sky130_fd_sc_hd__o21ai_1 _17057_ (.A1(_09793_),
    .A2(_09162_),
    .B1(_10078_),
    .Y(_10080_));
 sky130_fd_sc_hd__and2_1 _17058_ (.A(_10079_),
    .B(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__or2_1 _17059_ (.A(_08590_),
    .B(_09192_),
    .X(_10082_));
 sky130_fd_sc_hd__o21a_1 _17060_ (.A1(_08590_),
    .A2(_09064_),
    .B1(_09800_),
    .X(_10083_));
 sky130_fd_sc_hd__o21ba_1 _17061_ (.A1(_09802_),
    .A2(_10082_),
    .B1_N(_10083_),
    .X(_10084_));
 sky130_fd_sc_hd__nor2_1 _17062_ (.A(_09417_),
    .B(_08387_),
    .Y(_10085_));
 sky130_fd_sc_hd__xnor2_1 _17063_ (.A(_10084_),
    .B(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__a21oi_1 _17064_ (.A1(_09672_),
    .A2(_09804_),
    .B1(_09801_),
    .Y(_10087_));
 sky130_fd_sc_hd__nor2_1 _17065_ (.A(_10086_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__and2_1 _17066_ (.A(_10086_),
    .B(_10087_),
    .X(_10089_));
 sky130_fd_sc_hd__nor2_1 _17067_ (.A(_10088_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__xnor2_1 _17068_ (.A(_10081_),
    .B(_10090_),
    .Y(_10091_));
 sky130_fd_sc_hd__xor2_1 _17069_ (.A(_10074_),
    .B(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__xnor2_1 _17070_ (.A(_10072_),
    .B(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__a2bb2o_1 _17071_ (.A1_N(_09815_),
    .A2_N(_09818_),
    .B1(_09816_),
    .B2(_09701_),
    .X(_10094_));
 sky130_fd_sc_hd__o21ba_1 _17072_ (.A1(_09823_),
    .A2(_09828_),
    .B1_N(_09827_),
    .X(_10095_));
 sky130_fd_sc_hd__or3_1 _17073_ (.A(_08858_),
    .B(_09695_),
    .C(_09817_),
    .X(_10096_));
 sky130_fd_sc_hd__o22ai_1 _17074_ (.A1(_08858_),
    .A2(_09326_),
    .B1(_09696_),
    .B2(_08868_),
    .Y(_10097_));
 sky130_fd_sc_hd__nand2_1 _17075_ (.A(_10096_),
    .B(_10097_),
    .Y(_10098_));
 sky130_fd_sc_hd__nor2_1 _17076_ (.A(_08533_),
    .B(_09198_),
    .Y(_10099_));
 sky130_fd_sc_hd__xnor2_1 _17077_ (.A(_10098_),
    .B(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__xnor2_1 _17078_ (.A(_10095_),
    .B(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__xor2_1 _17079_ (.A(_10094_),
    .B(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__nor2_1 _17080_ (.A(_09700_),
    .B(_09697_),
    .Y(_10103_));
 sky130_fd_sc_hd__a21oi_4 _17081_ (.A1(_08292_),
    .A2(_09572_),
    .B1(_09824_),
    .Y(_10104_));
 sky130_fd_sc_hd__nor2_1 _17082_ (.A(_09002_),
    .B(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__o22a_1 _17083_ (.A1(_09002_),
    .A2(_09705_),
    .B1(_10104_),
    .B2(_08977_),
    .X(_10106_));
 sky130_fd_sc_hd__a21oi_1 _17084_ (.A1(_09826_),
    .A2(_10105_),
    .B1(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__xor2_1 _17085_ (.A(_10103_),
    .B(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__nand2_1 _17086_ (.A(_09755_),
    .B(_09833_),
    .Y(_10109_));
 sky130_fd_sc_hd__a2bb2o_1 _17087_ (.A1_N(_08217_),
    .A2_N(_09833_),
    .B1(_10109_),
    .B2(_09836_),
    .X(_10110_));
 sky130_fd_sc_hd__nand2_2 _17088_ (.A(\rbzero.wall_tracer.stepDistX[10] ),
    .B(_06100_),
    .Y(_10111_));
 sky130_fd_sc_hd__nand2_1 _17089_ (.A(\rbzero.wall_tracer.stepDistY[10] ),
    .B(_09069_),
    .Y(_10112_));
 sky130_fd_sc_hd__a21o_1 _17090_ (.A1(_09832_),
    .A2(_10112_),
    .B1(_06100_),
    .X(_10113_));
 sky130_fd_sc_hd__a21o_2 _17091_ (.A1(_10111_),
    .A2(_10113_),
    .B1(_08965_),
    .X(_10114_));
 sky130_fd_sc_hd__a21o_2 _17092_ (.A1(_09835_),
    .A2(_09711_),
    .B1(_06101_),
    .X(_10115_));
 sky130_fd_sc_hd__nand2_2 _17093_ (.A(\rbzero.wall_tracer.stepDistX[9] ),
    .B(_06101_),
    .Y(_10116_));
 sky130_fd_sc_hd__a21oi_1 _17094_ (.A1(_10115_),
    .A2(_10116_),
    .B1(_08965_),
    .Y(_10117_));
 sky130_fd_sc_hd__or3_1 _17095_ (.A(_08169_),
    .B(_08390_),
    .C(_09832_),
    .X(_10118_));
 sky130_fd_sc_hd__mux2_1 _17096_ (.A0(_08646_),
    .A1(_10118_),
    .S(_09833_),
    .X(_10119_));
 sky130_fd_sc_hd__mux2_1 _17097_ (.A0(_10114_),
    .A1(_10117_),
    .S(_10119_),
    .X(_10120_));
 sky130_fd_sc_hd__xor2_2 _17098_ (.A(_10110_),
    .B(_10120_),
    .X(_10121_));
 sky130_fd_sc_hd__xnor2_1 _17099_ (.A(_10108_),
    .B(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__nor2_1 _17100_ (.A(_09837_),
    .B(_09839_),
    .Y(_10123_));
 sky130_fd_sc_hd__a21o_1 _17101_ (.A1(_09830_),
    .A2(_09840_),
    .B1(_10123_),
    .X(_10124_));
 sky130_fd_sc_hd__xnor2_1 _17102_ (.A(_10122_),
    .B(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__xnor2_1 _17103_ (.A(_10102_),
    .B(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__or2b_1 _17104_ (.A(_09841_),
    .B_N(_09843_),
    .X(_10127_));
 sky130_fd_sc_hd__a21bo_1 _17105_ (.A1(_09822_),
    .A2(_09844_),
    .B1_N(_10127_),
    .X(_10128_));
 sky130_fd_sc_hd__xnor2_1 _17106_ (.A(_10126_),
    .B(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__xnor2_1 _17107_ (.A(_10093_),
    .B(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__and2b_1 _17108_ (.A_N(_09845_),
    .B(_09847_),
    .X(_10131_));
 sky130_fd_sc_hd__a21oi_1 _17109_ (.A1(_09812_),
    .A2(_09848_),
    .B1(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__or2_1 _17110_ (.A(_10130_),
    .B(_10132_),
    .X(_10133_));
 sky130_fd_sc_hd__nand2_1 _17111_ (.A(_10130_),
    .B(_10132_),
    .Y(_10134_));
 sky130_fd_sc_hd__and2_1 _17112_ (.A(_10133_),
    .B(_10134_),
    .X(_10135_));
 sky130_fd_sc_hd__xnor2_1 _17113_ (.A(_10071_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__or2b_1 _17114_ (.A(_09849_),
    .B_N(_09850_),
    .X(_10137_));
 sky130_fd_sc_hd__a21boi_1 _17115_ (.A1(_09789_),
    .A2(_09851_),
    .B1_N(_10137_),
    .Y(_10138_));
 sky130_fd_sc_hd__xor2_1 _17116_ (.A(_10136_),
    .B(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__nand2_1 _17117_ (.A(_10036_),
    .B(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__or2_1 _17118_ (.A(_10036_),
    .B(_10139_),
    .X(_10141_));
 sky130_fd_sc_hd__nand2_1 _17119_ (.A(_10140_),
    .B(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__o2bb2a_1 _17120_ (.A1_N(_09757_),
    .A2_N(_09854_),
    .B1(_09853_),
    .B2(_09852_),
    .X(_10143_));
 sky130_fd_sc_hd__xor2_1 _17121_ (.A(_10142_),
    .B(_10143_),
    .X(_10144_));
 sky130_fd_sc_hd__nand2_1 _17122_ (.A(_10031_),
    .B(_10144_),
    .Y(_10145_));
 sky130_fd_sc_hd__or2_1 _17123_ (.A(_10031_),
    .B(_10144_),
    .X(_10146_));
 sky130_fd_sc_hd__and2_2 _17124_ (.A(_10145_),
    .B(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__xor2_4 _17125_ (.A(_10029_),
    .B(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__inv_2 _17126_ (.A(_09858_),
    .Y(_10149_));
 sky130_fd_sc_hd__a21o_1 _17127_ (.A1(_09749_),
    .A2(_09735_),
    .B1(_09857_),
    .X(_10150_));
 sky130_fd_sc_hd__o31a_4 _17128_ (.A1(_09623_),
    .A2(_09737_),
    .A3(_10149_),
    .B1(_10150_),
    .X(_10151_));
 sky130_fd_sc_hd__xnor2_4 _17129_ (.A(_10148_),
    .B(_10151_),
    .Y(_10152_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(_06288_),
    .B(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__or2_1 _17131_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .X(_10154_));
 sky130_fd_sc_hd__nand2_1 _17132_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_10155_));
 sky130_fd_sc_hd__a211oi_1 _17133_ (.A1(_10154_),
    .A2(_10155_),
    .B1(_10021_),
    .C1(_10024_),
    .Y(_10156_));
 sky130_fd_sc_hd__o211a_1 _17134_ (.A1(_10021_),
    .A2(_10024_),
    .B1(_10154_),
    .C1(_10155_),
    .X(_10157_));
 sky130_fd_sc_hd__o31a_1 _17135_ (.A1(_06288_),
    .A2(_10156_),
    .A3(_10157_),
    .B1(_09945_),
    .X(_10158_));
 sky130_fd_sc_hd__o2bb2a_1 _17136_ (.A1_N(_10153_),
    .A2_N(_10158_),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_09946_),
    .X(_00539_));
 sky130_fd_sc_hd__or2_1 _17137_ (.A(_10142_),
    .B(_10143_),
    .X(_10159_));
 sky130_fd_sc_hd__nand2_2 _17138_ (.A(_10159_),
    .B(_10145_),
    .Y(_10160_));
 sky130_fd_sc_hd__or2b_1 _17139_ (.A(_10070_),
    .B_N(_10037_),
    .X(_10161_));
 sky130_fd_sc_hd__o21ba_1 _17140_ (.A1(_10047_),
    .A2(_10049_),
    .B1_N(_10046_),
    .X(_10162_));
 sky130_fd_sc_hd__a21oi_1 _17141_ (.A1(_10068_),
    .A2(_10161_),
    .B1(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__and3_1 _17142_ (.A(_10068_),
    .B(_10161_),
    .C(_10162_),
    .X(_10164_));
 sky130_fd_sc_hd__nor2_1 _17143_ (.A(_10163_),
    .B(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__nand2_1 _17144_ (.A(_10071_),
    .B(_10135_),
    .Y(_10166_));
 sky130_fd_sc_hd__a21o_1 _17145_ (.A1(_10050_),
    .A2(_10066_),
    .B1(_10064_),
    .X(_10167_));
 sky130_fd_sc_hd__or2b_1 _17146_ (.A(_10091_),
    .B_N(_10074_),
    .X(_10168_));
 sky130_fd_sc_hd__or2b_1 _17147_ (.A(_10092_),
    .B_N(_10072_),
    .X(_10169_));
 sky130_fd_sc_hd__nand2_1 _17148_ (.A(_10168_),
    .B(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__o22a_1 _17149_ (.A1(_09404_),
    .A2(_09377_),
    .B1(_09503_),
    .B2(_09409_),
    .X(_10171_));
 sky130_fd_sc_hd__or2_1 _17150_ (.A(_08888_),
    .B(_09502_),
    .X(_10172_));
 sky130_fd_sc_hd__or3_1 _17151_ (.A(_09409_),
    .B(_09377_),
    .C(_10172_),
    .X(_10173_));
 sky130_fd_sc_hd__and2b_1 _17152_ (.A_N(_10171_),
    .B(_10173_),
    .X(_10174_));
 sky130_fd_sc_hd__nor2_1 _17153_ (.A(_09157_),
    .B(_09637_),
    .Y(_10175_));
 sky130_fd_sc_hd__xnor2_1 _17154_ (.A(_10174_),
    .B(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__nand2_1 _17155_ (.A(_09761_),
    .B(_10040_),
    .Y(_10177_));
 sky130_fd_sc_hd__o31a_1 _17156_ (.A1(_09135_),
    .A2(_09637_),
    .A3(_10041_),
    .B1(_10177_),
    .X(_10178_));
 sky130_fd_sc_hd__xor2_1 _17157_ (.A(_10176_),
    .B(_10178_),
    .X(_10179_));
 sky130_fd_sc_hd__and2_1 _17158_ (.A(_09135_),
    .B(_10030_),
    .X(_10180_));
 sky130_fd_sc_hd__xor2_1 _17159_ (.A(_10179_),
    .B(_10180_),
    .X(_10181_));
 sky130_fd_sc_hd__o31ai_2 _17160_ (.A1(_09404_),
    .A2(_09511_),
    .A3(_10056_),
    .B1(_10055_),
    .Y(_10182_));
 sky130_fd_sc_hd__o22ai_1 _17161_ (.A1(_09793_),
    .A2(_09133_),
    .B1(_09225_),
    .B2(_09526_),
    .Y(_10183_));
 sky130_fd_sc_hd__or3_1 _17162_ (.A(_08422_),
    .B(_09225_),
    .C(_09773_),
    .X(_10184_));
 sky130_fd_sc_hd__nand2_1 _17163_ (.A(_10183_),
    .B(_10184_),
    .Y(_10185_));
 sky130_fd_sc_hd__nor2_1 _17164_ (.A(_09406_),
    .B(_09511_),
    .Y(_10186_));
 sky130_fd_sc_hd__xor2_1 _17165_ (.A(_10185_),
    .B(_10186_),
    .X(_10187_));
 sky130_fd_sc_hd__a21oi_1 _17166_ (.A1(_10077_),
    .A2(_10079_),
    .B1(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__and3_1 _17167_ (.A(_10077_),
    .B(_10079_),
    .C(_10187_),
    .X(_10189_));
 sky130_fd_sc_hd__nor2_1 _17168_ (.A(_10188_),
    .B(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__xnor2_1 _17169_ (.A(_10182_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__a21oi_1 _17170_ (.A1(_10052_),
    .A2(_10061_),
    .B1(_10059_),
    .Y(_10192_));
 sky130_fd_sc_hd__nor2_1 _17171_ (.A(_10191_),
    .B(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__and2_1 _17172_ (.A(_10191_),
    .B(_10192_),
    .X(_10194_));
 sky130_fd_sc_hd__nor2_1 _17173_ (.A(_10193_),
    .B(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__xor2_1 _17174_ (.A(_10181_),
    .B(_10195_),
    .X(_10196_));
 sky130_fd_sc_hd__xnor2_1 _17175_ (.A(_10170_),
    .B(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__xnor2_1 _17176_ (.A(_10167_),
    .B(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__a21o_1 _17177_ (.A1(_10081_),
    .A2(_10090_),
    .B1(_10088_),
    .X(_10199_));
 sky130_fd_sc_hd__and2b_1 _17178_ (.A_N(_10095_),
    .B(_10100_),
    .X(_10200_));
 sky130_fd_sc_hd__a21o_1 _17179_ (.A1(_10094_),
    .A2(_10101_),
    .B1(_10200_),
    .X(_10201_));
 sky130_fd_sc_hd__nor2_1 _17180_ (.A(_09158_),
    .B(_10075_),
    .Y(_10202_));
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08554_),
    .Y(_10203_));
 sky130_fd_sc_hd__nand2_1 _17182_ (.A(_08292_),
    .B(_08303_),
    .Y(_10204_));
 sky130_fd_sc_hd__clkbuf_2 _17183_ (.A(_10204_),
    .X(_10205_));
 sky130_fd_sc_hd__nor2_1 _17184_ (.A(_10203_),
    .B(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__xnor2_1 _17185_ (.A(_10202_),
    .B(_10206_),
    .Y(_10207_));
 sky130_fd_sc_hd__clkbuf_4 _17186_ (.A(_08349_),
    .X(_10208_));
 sky130_fd_sc_hd__nor2_1 _17187_ (.A(_10208_),
    .B(_09162_),
    .Y(_10209_));
 sky130_fd_sc_hd__xnor2_1 _17188_ (.A(_10207_),
    .B(_10209_),
    .Y(_10210_));
 sky130_fd_sc_hd__or3_1 _17189_ (.A(_08590_),
    .B(_09198_),
    .C(_09800_),
    .X(_10211_));
 sky130_fd_sc_hd__o22ai_1 _17190_ (.A1(_08590_),
    .A2(_09192_),
    .B1(_09198_),
    .B2(_08674_),
    .Y(_10212_));
 sky130_fd_sc_hd__and2_1 _17191_ (.A(_10211_),
    .B(_10212_),
    .X(_10213_));
 sky130_fd_sc_hd__nor2_1 _17192_ (.A(_09417_),
    .B(_09064_),
    .Y(_10214_));
 sky130_fd_sc_hd__xnor2_1 _17193_ (.A(_10213_),
    .B(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__a2bb2oi_1 _17194_ (.A1_N(_09802_),
    .A2_N(_10082_),
    .B1(_10084_),
    .B2(_10085_),
    .Y(_10216_));
 sky130_fd_sc_hd__nor2_1 _17195_ (.A(_10215_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__nand2_1 _17196_ (.A(_10215_),
    .B(_10216_),
    .Y(_10218_));
 sky130_fd_sc_hd__and2b_1 _17197_ (.A_N(_10217_),
    .B(_10218_),
    .X(_10219_));
 sky130_fd_sc_hd__xor2_1 _17198_ (.A(_10210_),
    .B(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__xnor2_1 _17199_ (.A(_10201_),
    .B(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__xnor2_1 _17200_ (.A(_10199_),
    .B(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__a21bo_1 _17201_ (.A1(_10097_),
    .A2(_10099_),
    .B1_N(_10096_),
    .X(_10223_));
 sky130_fd_sc_hd__a22oi_2 _17202_ (.A1(_09826_),
    .A2(_10105_),
    .B1(_10107_),
    .B2(_10103_),
    .Y(_10224_));
 sky130_fd_sc_hd__nor2_1 _17203_ (.A(_08858_),
    .B(_09696_),
    .Y(_10225_));
 sky130_fd_sc_hd__a21oi_2 _17204_ (.A1(_09565_),
    .A2(_09566_),
    .B1(_08868_),
    .Y(_10226_));
 sky130_fd_sc_hd__xnor2_1 _17205_ (.A(_10225_),
    .B(_10226_),
    .Y(_10227_));
 sky130_fd_sc_hd__buf_2 _17206_ (.A(_08533_),
    .X(_10228_));
 sky130_fd_sc_hd__nor2_1 _17207_ (.A(_10228_),
    .B(_09326_),
    .Y(_10229_));
 sky130_fd_sc_hd__xnor2_1 _17208_ (.A(_10227_),
    .B(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__xnor2_1 _17209_ (.A(_10224_),
    .B(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__xor2_1 _17210_ (.A(_10223_),
    .B(_10231_),
    .X(_10232_));
 sky130_fd_sc_hd__nor2_1 _17211_ (.A(_09700_),
    .B(_09706_),
    .Y(_10233_));
 sky130_fd_sc_hd__a21o_1 _17212_ (.A1(_10115_),
    .A2(_10116_),
    .B1(_08977_),
    .X(_10234_));
 sky130_fd_sc_hd__xnor2_1 _17213_ (.A(_10105_),
    .B(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__xor2_2 _17214_ (.A(_10233_),
    .B(_10235_),
    .X(_10236_));
 sky130_fd_sc_hd__and2_1 _17215_ (.A(_09833_),
    .B(_10118_),
    .X(_10237_));
 sky130_fd_sc_hd__nor3_4 _17216_ (.A(_09081_),
    .B(_09833_),
    .C(_10114_),
    .Y(_10238_));
 sky130_fd_sc_hd__a21oi_4 _17217_ (.A1(_10237_),
    .A2(_10114_),
    .B1(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__xnor2_1 _17218_ (.A(_10236_),
    .B(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__and2_1 _17219_ (.A(_10110_),
    .B(_10120_),
    .X(_10241_));
 sky130_fd_sc_hd__a21oi_2 _17220_ (.A1(_10108_),
    .A2(_10121_),
    .B1(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__xor2_1 _17221_ (.A(_10240_),
    .B(_10242_),
    .X(_10243_));
 sky130_fd_sc_hd__xnor2_1 _17222_ (.A(_10232_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__or2b_1 _17223_ (.A(_10122_),
    .B_N(_10124_),
    .X(_10245_));
 sky130_fd_sc_hd__a21bo_1 _17224_ (.A1(_10102_),
    .A2(_10125_),
    .B1_N(_10245_),
    .X(_10246_));
 sky130_fd_sc_hd__xnor2_1 _17225_ (.A(_10244_),
    .B(_10246_),
    .Y(_10247_));
 sky130_fd_sc_hd__xnor2_1 _17226_ (.A(_10222_),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__and2b_1 _17227_ (.A_N(_10126_),
    .B(_10128_),
    .X(_10249_));
 sky130_fd_sc_hd__a21oi_1 _17228_ (.A1(_10093_),
    .A2(_10129_),
    .B1(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__nor2_1 _17229_ (.A(_10248_),
    .B(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__and2_1 _17230_ (.A(_10248_),
    .B(_10250_),
    .X(_10252_));
 sky130_fd_sc_hd__nor2_1 _17231_ (.A(_10251_),
    .B(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__xnor2_1 _17232_ (.A(_10198_),
    .B(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__a21oi_1 _17233_ (.A1(_10133_),
    .A2(_10166_),
    .B1(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__and3_1 _17234_ (.A(_10133_),
    .B(_10166_),
    .C(_10254_),
    .X(_10256_));
 sky130_fd_sc_hd__nor2_1 _17235_ (.A(_10255_),
    .B(_10256_),
    .Y(_10257_));
 sky130_fd_sc_hd__xnor2_1 _17236_ (.A(_10165_),
    .B(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__o21a_1 _17237_ (.A1(_10136_),
    .A2(_10138_),
    .B1(_10140_),
    .X(_10259_));
 sky130_fd_sc_hd__nor2_1 _17238_ (.A(_10258_),
    .B(_10259_),
    .Y(_10260_));
 sky130_fd_sc_hd__and2_1 _17239_ (.A(_10258_),
    .B(_10259_),
    .X(_10261_));
 sky130_fd_sc_hd__nor2_2 _17240_ (.A(_10260_),
    .B(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__xnor2_4 _17241_ (.A(_10034_),
    .B(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__xnor2_4 _17242_ (.A(_10160_),
    .B(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__nor2_1 _17243_ (.A(_10029_),
    .B(_10147_),
    .Y(_10265_));
 sky130_fd_sc_hd__nand2_1 _17244_ (.A(_10029_),
    .B(_10147_),
    .Y(_10266_));
 sky130_fd_sc_hd__o21ai_2 _17245_ (.A1(_10265_),
    .A2(_10151_),
    .B1(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__xor2_4 _17246_ (.A(_10264_),
    .B(_10267_),
    .X(_10268_));
 sky130_fd_sc_hd__nand2_1 _17247_ (.A(_09915_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__nand2_1 _17248_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_10270_));
 sky130_fd_sc_hd__or2_1 _17249_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_10271_));
 sky130_fd_sc_hd__a21o_1 _17250_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(\rbzero.wall_tracer.stepDistX[0] ),
    .B1(_10157_),
    .X(_10272_));
 sky130_fd_sc_hd__and3_1 _17251_ (.A(_10270_),
    .B(_10271_),
    .C(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__a21o_1 _17252_ (.A1(_10270_),
    .A2(_10271_),
    .B1(_10272_),
    .X(_10274_));
 sky130_fd_sc_hd__or3b_1 _17253_ (.A(_09974_),
    .B(_10273_),
    .C_N(_10274_),
    .X(_10275_));
 sky130_fd_sc_hd__nand2_1 _17254_ (.A(_10269_),
    .B(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__mux2_1 _17255_ (.A0(\rbzero.wall_tracer.trackDistX[1] ),
    .A1(_10276_),
    .S(_09978_),
    .X(_10277_));
 sky130_fd_sc_hd__clkbuf_1 _17256_ (.A(_10277_),
    .X(_00540_));
 sky130_fd_sc_hd__nand2_1 _17257_ (.A(_10170_),
    .B(_10196_),
    .Y(_10278_));
 sky130_fd_sc_hd__or2b_1 _17258_ (.A(_10197_),
    .B_N(_10167_),
    .X(_10279_));
 sky130_fd_sc_hd__o2bb2a_1 _17259_ (.A1_N(_10179_),
    .A2_N(_10180_),
    .B1(_10176_),
    .B2(_10178_),
    .X(_10280_));
 sky130_fd_sc_hd__a21oi_1 _17260_ (.A1(_10278_),
    .A2(_10279_),
    .B1(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__and3_1 _17261_ (.A(_10278_),
    .B(_10279_),
    .C(_10280_),
    .X(_10282_));
 sky130_fd_sc_hd__nor2_1 _17262_ (.A(_10281_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__a21o_1 _17263_ (.A1(_10181_),
    .A2(_10195_),
    .B1(_10193_),
    .X(_10284_));
 sky130_fd_sc_hd__or2b_1 _17264_ (.A(_10221_),
    .B_N(_10199_),
    .X(_10285_));
 sky130_fd_sc_hd__a21bo_1 _17265_ (.A1(_10201_),
    .A2(_10220_),
    .B1_N(_10285_),
    .X(_10286_));
 sky130_fd_sc_hd__o21ai_1 _17266_ (.A1(_09406_),
    .A2(_09378_),
    .B1(_10172_),
    .Y(_10287_));
 sky130_fd_sc_hd__or2_1 _17267_ (.A(_09406_),
    .B(_09502_),
    .X(_10288_));
 sky130_fd_sc_hd__or3_1 _17268_ (.A(_09404_),
    .B(_09377_),
    .C(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__nand2_1 _17269_ (.A(_10287_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__nor2_1 _17270_ (.A(_09409_),
    .B(_09636_),
    .Y(_10291_));
 sky130_fd_sc_hd__xor2_1 _17271_ (.A(_10290_),
    .B(_10291_),
    .X(_10292_));
 sky130_fd_sc_hd__o31a_1 _17272_ (.A1(_09157_),
    .A2(_09637_),
    .A3(_10171_),
    .B1(_10173_),
    .X(_10293_));
 sky130_fd_sc_hd__xor2_1 _17273_ (.A(_10292_),
    .B(_10293_),
    .X(_10294_));
 sky130_fd_sc_hd__and2_1 _17274_ (.A(_09157_),
    .B(_10030_),
    .X(_10295_));
 sky130_fd_sc_hd__xor2_1 _17275_ (.A(_10294_),
    .B(_10295_),
    .X(_10296_));
 sky130_fd_sc_hd__a21bo_1 _17276_ (.A1(_10183_),
    .A2(_10186_),
    .B1_N(_10184_),
    .X(_10297_));
 sky130_fd_sc_hd__or2_1 _17277_ (.A(_08422_),
    .B(_09225_),
    .X(_10298_));
 sky130_fd_sc_hd__or2_1 _17278_ (.A(_08349_),
    .B(_09133_),
    .X(_10299_));
 sky130_fd_sc_hd__xnor2_1 _17279_ (.A(_10298_),
    .B(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__nor2_1 _17280_ (.A(_09526_),
    .B(_09511_),
    .Y(_10301_));
 sky130_fd_sc_hd__xor2_1 _17281_ (.A(_10300_),
    .B(_10301_),
    .X(_10302_));
 sky130_fd_sc_hd__nand2_1 _17282_ (.A(_10202_),
    .B(_10206_),
    .Y(_10303_));
 sky130_fd_sc_hd__o31ai_1 _17283_ (.A1(_10208_),
    .A2(_09162_),
    .A3(_10207_),
    .B1(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__and2b_1 _17284_ (.A_N(_10302_),
    .B(_10304_),
    .X(_10305_));
 sky130_fd_sc_hd__and2b_1 _17285_ (.A_N(_10304_),
    .B(_10302_),
    .X(_10306_));
 sky130_fd_sc_hd__nor2_1 _17286_ (.A(_10305_),
    .B(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__xnor2_1 _17287_ (.A(_10297_),
    .B(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__a21oi_1 _17288_ (.A1(_10182_),
    .A2(_10190_),
    .B1(_10188_),
    .Y(_10309_));
 sky130_fd_sc_hd__nor2_1 _17289_ (.A(_10308_),
    .B(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__and2_1 _17290_ (.A(_10308_),
    .B(_10309_),
    .X(_10311_));
 sky130_fd_sc_hd__nor2_1 _17291_ (.A(_10310_),
    .B(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__xor2_1 _17292_ (.A(_10296_),
    .B(_10312_),
    .X(_10313_));
 sky130_fd_sc_hd__xnor2_1 _17293_ (.A(_10286_),
    .B(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__xnor2_1 _17294_ (.A(_10284_),
    .B(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__a21o_1 _17295_ (.A1(_10210_),
    .A2(_10218_),
    .B1(_10217_),
    .X(_10316_));
 sky130_fd_sc_hd__and2b_1 _17296_ (.A_N(_10224_),
    .B(_10230_),
    .X(_10317_));
 sky130_fd_sc_hd__a21oi_1 _17297_ (.A1(_10223_),
    .A2(_10231_),
    .B1(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__a2bb2o_1 _17298_ (.A1_N(_08545_),
    .A2_N(_08360_),
    .B1(_08556_),
    .B2(_08303_),
    .X(_10319_));
 sky130_fd_sc_hd__or4_2 _17299_ (.A(_10203_),
    .B(_08555_),
    .C(_10204_),
    .D(_08394_),
    .X(_10320_));
 sky130_fd_sc_hd__nand2_1 _17300_ (.A(_10319_),
    .B(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__or3_1 _17301_ (.A(_10075_),
    .B(_09162_),
    .C(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__o21ai_1 _17302_ (.A1(_10075_),
    .A2(_09162_),
    .B1(_10321_),
    .Y(_10323_));
 sky130_fd_sc_hd__and2_1 _17303_ (.A(_10322_),
    .B(_10323_),
    .X(_10324_));
 sky130_fd_sc_hd__nor2_1 _17304_ (.A(_09671_),
    .B(_09198_),
    .Y(_10325_));
 sky130_fd_sc_hd__nor2_1 _17305_ (.A(_08674_),
    .B(_09326_),
    .Y(_10326_));
 sky130_fd_sc_hd__xnor2_1 _17306_ (.A(_10325_),
    .B(_10326_),
    .Y(_10327_));
 sky130_fd_sc_hd__or2_1 _17307_ (.A(_09417_),
    .B(_09192_),
    .X(_10328_));
 sky130_fd_sc_hd__xnor2_1 _17308_ (.A(_10327_),
    .B(_10328_),
    .Y(_10329_));
 sky130_fd_sc_hd__a21boi_1 _17309_ (.A1(_10213_),
    .A2(_10214_),
    .B1_N(_10211_),
    .Y(_10330_));
 sky130_fd_sc_hd__nor2_1 _17310_ (.A(_10329_),
    .B(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(_10329_),
    .B(_10330_),
    .Y(_10332_));
 sky130_fd_sc_hd__and2b_1 _17312_ (.A_N(_10331_),
    .B(_10332_),
    .X(_10333_));
 sky130_fd_sc_hd__xor2_1 _17313_ (.A(_10324_),
    .B(_10333_),
    .X(_10334_));
 sky130_fd_sc_hd__xnor2_1 _17314_ (.A(_10318_),
    .B(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__xor2_1 _17315_ (.A(_10316_),
    .B(_10335_),
    .X(_10336_));
 sky130_fd_sc_hd__nand2_1 _17316_ (.A(_10225_),
    .B(_10226_),
    .Y(_10337_));
 sky130_fd_sc_hd__o31ai_2 _17317_ (.A1(_10228_),
    .A2(_09326_),
    .A3(_10227_),
    .B1(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__or2_1 _17318_ (.A(_08977_),
    .B(_10104_),
    .X(_10339_));
 sky130_fd_sc_hd__a21o_1 _17319_ (.A1(_10115_),
    .A2(_10116_),
    .B1(_09002_),
    .X(_10340_));
 sky130_fd_sc_hd__a2bb2o_1 _17320_ (.A1_N(_10339_),
    .A2_N(_10340_),
    .B1(_10235_),
    .B2(_10233_),
    .X(_10341_));
 sky130_fd_sc_hd__or3b_1 _17321_ (.A(_08858_),
    .B(_09706_),
    .C_N(_10226_),
    .X(_10342_));
 sky130_fd_sc_hd__o22ai_1 _17322_ (.A1(_08858_),
    .A2(_09697_),
    .B1(_09706_),
    .B2(_08868_),
    .Y(_10343_));
 sky130_fd_sc_hd__nand2_1 _17323_ (.A(_10342_),
    .B(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__nor2_1 _17324_ (.A(_08533_),
    .B(_09696_),
    .Y(_10345_));
 sky130_fd_sc_hd__xnor2_1 _17325_ (.A(_10344_),
    .B(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__xor2_1 _17326_ (.A(_10341_),
    .B(_10346_),
    .X(_10347_));
 sky130_fd_sc_hd__xor2_1 _17327_ (.A(_10338_),
    .B(_10347_),
    .X(_10348_));
 sky130_fd_sc_hd__nor2_1 _17328_ (.A(_09700_),
    .B(_10104_),
    .Y(_10349_));
 sky130_fd_sc_hd__a21oi_1 _17329_ (.A1(_10111_),
    .A2(_10113_),
    .B1(_08977_),
    .Y(_10350_));
 sky130_fd_sc_hd__xnor2_1 _17330_ (.A(_10340_),
    .B(_10350_),
    .Y(_10351_));
 sky130_fd_sc_hd__xor2_2 _17331_ (.A(_10349_),
    .B(_10351_),
    .X(_10352_));
 sky130_fd_sc_hd__xor2_1 _17332_ (.A(_10239_),
    .B(_10352_),
    .X(_10353_));
 sky130_fd_sc_hd__a21o_1 _17333_ (.A1(_10236_),
    .A2(_10239_),
    .B1(_10238_),
    .X(_10354_));
 sky130_fd_sc_hd__xor2_1 _17334_ (.A(_10353_),
    .B(_10354_),
    .X(_10355_));
 sky130_fd_sc_hd__xnor2_1 _17335_ (.A(_10348_),
    .B(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__nor2_1 _17336_ (.A(_10240_),
    .B(_10242_),
    .Y(_10357_));
 sky130_fd_sc_hd__a21o_1 _17337_ (.A1(_10232_),
    .A2(_10243_),
    .B1(_10357_),
    .X(_10358_));
 sky130_fd_sc_hd__xnor2_1 _17338_ (.A(_10356_),
    .B(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__xnor2_1 _17339_ (.A(_10336_),
    .B(_10359_),
    .Y(_10360_));
 sky130_fd_sc_hd__and2b_1 _17340_ (.A_N(_10244_),
    .B(_10246_),
    .X(_10361_));
 sky130_fd_sc_hd__a21oi_1 _17341_ (.A1(_10222_),
    .A2(_10247_),
    .B1(_10361_),
    .Y(_10362_));
 sky130_fd_sc_hd__nor2_1 _17342_ (.A(_10360_),
    .B(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__and2_1 _17343_ (.A(_10360_),
    .B(_10362_),
    .X(_10364_));
 sky130_fd_sc_hd__nor2_1 _17344_ (.A(_10363_),
    .B(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__xnor2_1 _17345_ (.A(_10315_),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__a21oi_1 _17346_ (.A1(_10198_),
    .A2(_10253_),
    .B1(_10251_),
    .Y(_10367_));
 sky130_fd_sc_hd__nor2_1 _17347_ (.A(_10366_),
    .B(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__and2_1 _17348_ (.A(_10366_),
    .B(_10367_),
    .X(_10369_));
 sky130_fd_sc_hd__nor2_1 _17349_ (.A(_10368_),
    .B(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__xnor2_1 _17350_ (.A(_10283_),
    .B(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__a21oi_1 _17351_ (.A1(_10165_),
    .A2(_10257_),
    .B1(_10255_),
    .Y(_10372_));
 sky130_fd_sc_hd__xor2_1 _17352_ (.A(_10371_),
    .B(_10372_),
    .X(_10373_));
 sky130_fd_sc_hd__nand2_1 _17353_ (.A(_10163_),
    .B(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__or2_1 _17354_ (.A(_10163_),
    .B(_10373_),
    .X(_10375_));
 sky130_fd_sc_hd__nand2_1 _17355_ (.A(_10374_),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__a21oi_1 _17356_ (.A1(_10034_),
    .A2(_10262_),
    .B1(_10260_),
    .Y(_10377_));
 sky130_fd_sc_hd__or2_1 _17357_ (.A(_10376_),
    .B(_10377_),
    .X(_10378_));
 sky130_fd_sc_hd__nand2_1 _17358_ (.A(_10376_),
    .B(_10377_),
    .Y(_10379_));
 sky130_fd_sc_hd__and2_1 _17359_ (.A(_10378_),
    .B(_10379_),
    .X(_10380_));
 sky130_fd_sc_hd__nand2_1 _17360_ (.A(_10148_),
    .B(_10264_),
    .Y(_10381_));
 sky130_fd_sc_hd__a21o_1 _17361_ (.A1(_10159_),
    .A2(_10145_),
    .B1(_10263_),
    .X(_10382_));
 sky130_fd_sc_hd__and3_1 _17362_ (.A(_10159_),
    .B(_10145_),
    .C(_10263_),
    .X(_10383_));
 sky130_fd_sc_hd__a21o_1 _17363_ (.A1(_10266_),
    .A2(_10382_),
    .B1(_10383_),
    .X(_10384_));
 sky130_fd_sc_hd__o21ai_1 _17364_ (.A1(_10151_),
    .A2(_10381_),
    .B1(_10384_),
    .Y(_10385_));
 sky130_fd_sc_hd__nand2_1 _17365_ (.A(_10380_),
    .B(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__inv_2 _17366_ (.A(_10380_),
    .Y(_10387_));
 sky130_fd_sc_hd__o21a_1 _17367_ (.A1(_10151_),
    .A2(_10381_),
    .B1(_10384_),
    .X(_10388_));
 sky130_fd_sc_hd__nand2_1 _17368_ (.A(_10387_),
    .B(_10388_),
    .Y(_10389_));
 sky130_fd_sc_hd__and2_2 _17369_ (.A(_10386_),
    .B(_10389_),
    .X(_10390_));
 sky130_fd_sc_hd__nand2_1 _17370_ (.A(_06288_),
    .B(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__inv_2 _17371_ (.A(_10270_),
    .Y(_10392_));
 sky130_fd_sc_hd__nand2_1 _17372_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .Y(_10393_));
 sky130_fd_sc_hd__or2_1 _17373_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_10394_));
 sky130_fd_sc_hd__o211ai_2 _17374_ (.A1(_10392_),
    .A2(_10273_),
    .B1(_10393_),
    .C1(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__a211o_1 _17375_ (.A1(_10393_),
    .A2(_10394_),
    .B1(_10392_),
    .C1(_10273_),
    .X(_10396_));
 sky130_fd_sc_hd__a31oi_1 _17376_ (.A1(_09938_),
    .A2(_10395_),
    .A3(_10396_),
    .B1(_09919_),
    .Y(_10397_));
 sky130_fd_sc_hd__o2bb2a_1 _17377_ (.A1_N(_10391_),
    .A2_N(_10397_),
    .B1(\rbzero.wall_tracer.trackDistX[2] ),
    .B2(_09946_),
    .X(_00541_));
 sky130_fd_sc_hd__or2_1 _17378_ (.A(_10371_),
    .B(_10372_),
    .X(_10398_));
 sky130_fd_sc_hd__nand2_1 _17379_ (.A(_10286_),
    .B(_10313_),
    .Y(_10399_));
 sky130_fd_sc_hd__or2b_1 _17380_ (.A(_10314_),
    .B_N(_10284_),
    .X(_10400_));
 sky130_fd_sc_hd__o2bb2a_1 _17381_ (.A1_N(_10294_),
    .A2_N(_10295_),
    .B1(_10292_),
    .B2(_10293_),
    .X(_10401_));
 sky130_fd_sc_hd__a21oi_1 _17382_ (.A1(_10399_),
    .A2(_10400_),
    .B1(_10401_),
    .Y(_10402_));
 sky130_fd_sc_hd__and3_1 _17383_ (.A(_10399_),
    .B(_10400_),
    .C(_10401_),
    .X(_10403_));
 sky130_fd_sc_hd__nor2_1 _17384_ (.A(_10402_),
    .B(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__a21o_1 _17385_ (.A1(_10296_),
    .A2(_10312_),
    .B1(_10310_),
    .X(_10405_));
 sky130_fd_sc_hd__or2b_1 _17386_ (.A(_10318_),
    .B_N(_10334_),
    .X(_10406_));
 sky130_fd_sc_hd__a21bo_1 _17387_ (.A1(_10316_),
    .A2(_10335_),
    .B1_N(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__or2_1 _17388_ (.A(_09526_),
    .B(_09377_),
    .X(_10408_));
 sky130_fd_sc_hd__xnor2_1 _17389_ (.A(_10288_),
    .B(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__or3_1 _17390_ (.A(_09404_),
    .B(_09636_),
    .C(_10409_),
    .X(_10410_));
 sky130_fd_sc_hd__o21ai_1 _17391_ (.A1(_09404_),
    .A2(_09637_),
    .B1(_10409_),
    .Y(_10411_));
 sky130_fd_sc_hd__nand2_1 _17392_ (.A(_10410_),
    .B(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__o31a_1 _17393_ (.A1(_09409_),
    .A2(_09637_),
    .A3(_10290_),
    .B1(_10289_),
    .X(_10413_));
 sky130_fd_sc_hd__xnor2_1 _17394_ (.A(_10412_),
    .B(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__nor2_1 _17395_ (.A(_08962_),
    .B(_09755_),
    .Y(_10415_));
 sky130_fd_sc_hd__xnor2_1 _17396_ (.A(_10414_),
    .B(_10415_),
    .Y(_10416_));
 sky130_fd_sc_hd__or3_1 _17397_ (.A(_09526_),
    .B(_09511_),
    .C(_10300_),
    .X(_10417_));
 sky130_fd_sc_hd__o21ai_1 _17398_ (.A1(_10298_),
    .A2(_10299_),
    .B1(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__o22ai_1 _17399_ (.A1(_08509_),
    .A2(_09133_),
    .B1(_09225_),
    .B2(_08349_),
    .Y(_10419_));
 sky130_fd_sc_hd__or4_1 _17400_ (.A(_08509_),
    .B(_08349_),
    .C(_09132_),
    .D(_09222_),
    .X(_10420_));
 sky130_fd_sc_hd__nand2_1 _17401_ (.A(_10419_),
    .B(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__nor2_1 _17402_ (.A(_09793_),
    .B(_09276_),
    .Y(_10422_));
 sky130_fd_sc_hd__xor2_1 _17403_ (.A(_10421_),
    .B(_10422_),
    .X(_10423_));
 sky130_fd_sc_hd__a21oi_1 _17404_ (.A1(_10320_),
    .A2(_10322_),
    .B1(_10423_),
    .Y(_10424_));
 sky130_fd_sc_hd__and3_1 _17405_ (.A(_10320_),
    .B(_10322_),
    .C(_10423_),
    .X(_10425_));
 sky130_fd_sc_hd__nor2_1 _17406_ (.A(_10424_),
    .B(_10425_),
    .Y(_10426_));
 sky130_fd_sc_hd__xnor2_1 _17407_ (.A(_10418_),
    .B(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__a21oi_1 _17408_ (.A1(_10297_),
    .A2(_10307_),
    .B1(_10305_),
    .Y(_10428_));
 sky130_fd_sc_hd__nor2_1 _17409_ (.A(_10427_),
    .B(_10428_),
    .Y(_10429_));
 sky130_fd_sc_hd__and2_1 _17410_ (.A(_10427_),
    .B(_10428_),
    .X(_10430_));
 sky130_fd_sc_hd__nor2_1 _17411_ (.A(_10429_),
    .B(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__xor2_1 _17412_ (.A(_10416_),
    .B(_10431_),
    .X(_10432_));
 sky130_fd_sc_hd__nand2_1 _17413_ (.A(_10407_),
    .B(_10432_),
    .Y(_10433_));
 sky130_fd_sc_hd__or2_1 _17414_ (.A(_10407_),
    .B(_10432_),
    .X(_10434_));
 sky130_fd_sc_hd__nand2_1 _17415_ (.A(_10433_),
    .B(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__xnor2_1 _17416_ (.A(_10405_),
    .B(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__a21o_1 _17417_ (.A1(_10324_),
    .A2(_10332_),
    .B1(_10331_),
    .X(_10437_));
 sky130_fd_sc_hd__and2_1 _17418_ (.A(_10341_),
    .B(_10346_),
    .X(_10438_));
 sky130_fd_sc_hd__a21oi_1 _17419_ (.A1(_10338_),
    .A2(_10347_),
    .B1(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__nand2_1 _17420_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08554_),
    .Y(_10440_));
 sky130_fd_sc_hd__a2bb2o_1 _17421_ (.A1_N(_08555_),
    .A2_N(_08394_),
    .B1(_08391_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_10441_));
 sky130_fd_sc_hd__or4_1 _17422_ (.A(_06461_),
    .B(_08555_),
    .C(_08394_),
    .D(_08395_),
    .X(_10442_));
 sky130_fd_sc_hd__nand2_1 _17423_ (.A(_10441_),
    .B(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__or3_1 _17424_ (.A(_10205_),
    .B(_10440_),
    .C(_10443_),
    .X(_10444_));
 sky130_fd_sc_hd__buf_2 _17425_ (.A(_10440_),
    .X(_10445_));
 sky130_fd_sc_hd__o21ai_1 _17426_ (.A1(_10205_),
    .A2(_10445_),
    .B1(_10443_),
    .Y(_10446_));
 sky130_fd_sc_hd__and2_2 _17427_ (.A(_10444_),
    .B(_10446_),
    .X(_10447_));
 sky130_fd_sc_hd__or2_1 _17428_ (.A(_08590_),
    .B(_09326_),
    .X(_10448_));
 sky130_fd_sc_hd__or3_1 _17429_ (.A(_08674_),
    .B(_09695_),
    .C(_10448_),
    .X(_10449_));
 sky130_fd_sc_hd__o21ai_1 _17430_ (.A1(_08856_),
    .A2(_09696_),
    .B1(_10448_),
    .Y(_10450_));
 sky130_fd_sc_hd__nand2_1 _17431_ (.A(_10449_),
    .B(_10450_),
    .Y(_10451_));
 sky130_fd_sc_hd__or2_1 _17432_ (.A(_09417_),
    .B(_09198_),
    .X(_10452_));
 sky130_fd_sc_hd__xnor2_1 _17433_ (.A(_10451_),
    .B(_10452_),
    .Y(_10453_));
 sky130_fd_sc_hd__o2bb2a_1 _17434_ (.A1_N(_10325_),
    .A2_N(_10326_),
    .B1(_10327_),
    .B2(_10328_),
    .X(_10454_));
 sky130_fd_sc_hd__xor2_1 _17435_ (.A(_10453_),
    .B(_10454_),
    .X(_10455_));
 sky130_fd_sc_hd__xnor2_1 _17436_ (.A(_10447_),
    .B(_10455_),
    .Y(_10456_));
 sky130_fd_sc_hd__xnor2_1 _17437_ (.A(_10439_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__xnor2_1 _17438_ (.A(_10437_),
    .B(_10457_),
    .Y(_10458_));
 sky130_fd_sc_hd__a21bo_1 _17439_ (.A1(_10343_),
    .A2(_10345_),
    .B1_N(_10342_),
    .X(_10459_));
 sky130_fd_sc_hd__and2_1 _17440_ (.A(_10115_),
    .B(_10116_),
    .X(_10460_));
 sky130_fd_sc_hd__buf_2 _17441_ (.A(_10460_),
    .X(_10461_));
 sky130_fd_sc_hd__a211o_1 _17442_ (.A1(_10111_),
    .A2(_10113_),
    .B1(_08318_),
    .C1(_08413_),
    .X(_10462_));
 sky130_fd_sc_hd__a2bb2o_1 _17443_ (.A1_N(_10461_),
    .A2_N(_10462_),
    .B1(_10351_),
    .B2(_10349_),
    .X(_10463_));
 sky130_fd_sc_hd__nor2_1 _17444_ (.A(_08487_),
    .B(_09705_),
    .Y(_10464_));
 sky130_fd_sc_hd__nor2_1 _17445_ (.A(_08868_),
    .B(_10104_),
    .Y(_10465_));
 sky130_fd_sc_hd__xnor2_1 _17446_ (.A(_10464_),
    .B(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__nor2_1 _17447_ (.A(_08533_),
    .B(_09697_),
    .Y(_10467_));
 sky130_fd_sc_hd__xnor2_1 _17448_ (.A(_10466_),
    .B(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__xnor2_1 _17449_ (.A(_10463_),
    .B(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__xnor2_1 _17450_ (.A(_10459_),
    .B(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__and2_1 _17451_ (.A(_08318_),
    .B(_08413_),
    .X(_10471_));
 sky130_fd_sc_hd__and2_1 _17452_ (.A(_10111_),
    .B(_10113_),
    .X(_10472_));
 sky130_fd_sc_hd__buf_2 _17453_ (.A(_10472_),
    .X(_10473_));
 sky130_fd_sc_hd__or3b_1 _17454_ (.A(_10471_),
    .B(_10473_),
    .C_N(_10462_),
    .X(_10474_));
 sky130_fd_sc_hd__clkbuf_2 _17455_ (.A(_10474_),
    .X(_10475_));
 sky130_fd_sc_hd__nor2_1 _17456_ (.A(_09700_),
    .B(_10461_),
    .Y(_10476_));
 sky130_fd_sc_hd__xnor2_1 _17457_ (.A(_10475_),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__xnor2_1 _17458_ (.A(_10239_),
    .B(_10477_),
    .Y(_10478_));
 sky130_fd_sc_hd__a21oi_1 _17459_ (.A1(_10239_),
    .A2(_10352_),
    .B1(_10238_),
    .Y(_10479_));
 sky130_fd_sc_hd__xor2_1 _17460_ (.A(_10478_),
    .B(_10479_),
    .X(_10480_));
 sky130_fd_sc_hd__xnor2_1 _17461_ (.A(_10470_),
    .B(_10480_),
    .Y(_10481_));
 sky130_fd_sc_hd__nand2_1 _17462_ (.A(_10353_),
    .B(_10354_),
    .Y(_10482_));
 sky130_fd_sc_hd__a21bo_1 _17463_ (.A1(_10348_),
    .A2(_10355_),
    .B1_N(_10482_),
    .X(_10483_));
 sky130_fd_sc_hd__xnor2_1 _17464_ (.A(_10481_),
    .B(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__xnor2_1 _17465_ (.A(_10458_),
    .B(_10484_),
    .Y(_10485_));
 sky130_fd_sc_hd__and2b_1 _17466_ (.A_N(_10356_),
    .B(_10358_),
    .X(_10486_));
 sky130_fd_sc_hd__a21oi_1 _17467_ (.A1(_10336_),
    .A2(_10359_),
    .B1(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__nor2_1 _17468_ (.A(_10485_),
    .B(_10487_),
    .Y(_10488_));
 sky130_fd_sc_hd__and2_1 _17469_ (.A(_10485_),
    .B(_10487_),
    .X(_10489_));
 sky130_fd_sc_hd__nor2_1 _17470_ (.A(_10488_),
    .B(_10489_),
    .Y(_10490_));
 sky130_fd_sc_hd__xnor2_1 _17471_ (.A(_10436_),
    .B(_10490_),
    .Y(_10491_));
 sky130_fd_sc_hd__a21oi_1 _17472_ (.A1(_10315_),
    .A2(_10365_),
    .B1(_10363_),
    .Y(_10492_));
 sky130_fd_sc_hd__xor2_1 _17473_ (.A(_10491_),
    .B(_10492_),
    .X(_10493_));
 sky130_fd_sc_hd__nand2_1 _17474_ (.A(_10404_),
    .B(_10493_),
    .Y(_10494_));
 sky130_fd_sc_hd__or2_1 _17475_ (.A(_10404_),
    .B(_10493_),
    .X(_10495_));
 sky130_fd_sc_hd__nand2_1 _17476_ (.A(_10494_),
    .B(_10495_),
    .Y(_10496_));
 sky130_fd_sc_hd__a21oi_1 _17477_ (.A1(_10283_),
    .A2(_10370_),
    .B1(_10368_),
    .Y(_10497_));
 sky130_fd_sc_hd__xor2_1 _17478_ (.A(_10496_),
    .B(_10497_),
    .X(_10498_));
 sky130_fd_sc_hd__nand2_1 _17479_ (.A(_10281_),
    .B(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__or2_1 _17480_ (.A(_10281_),
    .B(_10498_),
    .X(_10500_));
 sky130_fd_sc_hd__nand2_1 _17481_ (.A(_10499_),
    .B(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__a21o_1 _17482_ (.A1(_10398_),
    .A2(_10374_),
    .B1(_10501_),
    .X(_10502_));
 sky130_fd_sc_hd__and3_1 _17483_ (.A(_10398_),
    .B(_10374_),
    .C(_10501_),
    .X(_10503_));
 sky130_fd_sc_hd__inv_2 _17484_ (.A(_10503_),
    .Y(_10504_));
 sky130_fd_sc_hd__nand2_1 _17485_ (.A(_10502_),
    .B(_10504_),
    .Y(_10505_));
 sky130_fd_sc_hd__a21oi_1 _17486_ (.A1(_10378_),
    .A2(_10386_),
    .B1(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__a31o_1 _17487_ (.A1(_10378_),
    .A2(_10386_),
    .A3(_10505_),
    .B1(_09937_),
    .X(_10507_));
 sky130_fd_sc_hd__or2_2 _17488_ (.A(_10506_),
    .B(_10507_),
    .X(_10508_));
 sky130_fd_sc_hd__buf_4 _17489_ (.A(_06287_),
    .X(_10509_));
 sky130_fd_sc_hd__and2_1 _17490_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_10510_));
 sky130_fd_sc_hd__nor2_1 _17491_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_10511_));
 sky130_fd_sc_hd__o211a_1 _17492_ (.A1(_10510_),
    .A2(_10511_),
    .B1(_10393_),
    .C1(_10395_),
    .X(_10512_));
 sky130_fd_sc_hd__a211oi_2 _17493_ (.A1(_10393_),
    .A2(_10395_),
    .B1(_10510_),
    .C1(_10511_),
    .Y(_10513_));
 sky130_fd_sc_hd__o31a_1 _17494_ (.A1(_10509_),
    .A2(_10512_),
    .A3(_10513_),
    .B1(_09945_),
    .X(_10514_));
 sky130_fd_sc_hd__o2bb2a_1 _17495_ (.A1_N(_10508_),
    .A2_N(_10514_),
    .B1(\rbzero.wall_tracer.trackDistX[3] ),
    .B2(_09946_),
    .X(_00542_));
 sky130_fd_sc_hd__or2b_1 _17496_ (.A(_10435_),
    .B_N(_10405_),
    .X(_10515_));
 sky130_fd_sc_hd__o32a_1 _17497_ (.A1(_08962_),
    .A2(_09755_),
    .A3(_10414_),
    .B1(_10413_),
    .B2(_10412_),
    .X(_10516_));
 sky130_fd_sc_hd__a21oi_2 _17498_ (.A1(_10433_),
    .A2(_10515_),
    .B1(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__and3_1 _17499_ (.A(_10433_),
    .B(_10515_),
    .C(_10516_),
    .X(_10518_));
 sky130_fd_sc_hd__nor2_1 _17500_ (.A(_10517_),
    .B(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__a21o_1 _17501_ (.A1(_10416_),
    .A2(_10431_),
    .B1(_10429_),
    .X(_10520_));
 sky130_fd_sc_hd__or2_1 _17502_ (.A(_10439_),
    .B(_10456_),
    .X(_01663_));
 sky130_fd_sc_hd__or2b_1 _17503_ (.A(_10457_),
    .B_N(_10437_),
    .X(_01664_));
 sky130_fd_sc_hd__nor2_1 _17504_ (.A(_09526_),
    .B(_09502_),
    .Y(_01665_));
 sky130_fd_sc_hd__nor2_1 _17505_ (.A(_09793_),
    .B(_09377_),
    .Y(_01666_));
 sky130_fd_sc_hd__xnor2_1 _17506_ (.A(_01665_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__or2_1 _17507_ (.A(_09406_),
    .B(_09636_),
    .X(_01668_));
 sky130_fd_sc_hd__xnor2_1 _17508_ (.A(_01667_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__o21a_1 _17509_ (.A1(_10288_),
    .A2(_10408_),
    .B1(_10410_),
    .X(_01670_));
 sky130_fd_sc_hd__xor2_1 _17510_ (.A(_01669_),
    .B(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__and2_1 _17511_ (.A(_09404_),
    .B(_10030_),
    .X(_01672_));
 sky130_fd_sc_hd__xor2_1 _17512_ (.A(_01671_),
    .B(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__a21bo_1 _17513_ (.A1(_10419_),
    .A2(_10422_),
    .B1_N(_10420_),
    .X(_01674_));
 sky130_fd_sc_hd__nand2_1 _17514_ (.A(_10442_),
    .B(_10444_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_4 _17515_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08554_),
    .Y(_01676_));
 sky130_fd_sc_hd__or2b_1 _17516_ (.A(_09222_),
    .B_N(_08323_),
    .X(_01677_));
 sky130_fd_sc_hd__or3_1 _17517_ (.A(_10205_),
    .B(_01676_),
    .C(_01677_),
    .X(_01678_));
 sky130_fd_sc_hd__o21ai_1 _17518_ (.A1(_10205_),
    .A2(_01676_),
    .B1(_01677_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _17519_ (.A(_01678_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__nor2_1 _17520_ (.A(_10208_),
    .B(_09511_),
    .Y(_01681_));
 sky130_fd_sc_hd__xor2_2 _17521_ (.A(_01680_),
    .B(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__xnor2_2 _17522_ (.A(_01675_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__xnor2_1 _17523_ (.A(_01674_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__a21oi_1 _17524_ (.A1(_10418_),
    .A2(_10426_),
    .B1(_10424_),
    .Y(_01685_));
 sky130_fd_sc_hd__nor2_1 _17525_ (.A(_01684_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__and2_1 _17526_ (.A(_01684_),
    .B(_01685_),
    .X(_01687_));
 sky130_fd_sc_hd__nor2_1 _17527_ (.A(_01686_),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__xnor2_1 _17528_ (.A(_01673_),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__a21o_1 _17529_ (.A1(_01663_),
    .A2(_01664_),
    .B1(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__nand3_1 _17530_ (.A(_01663_),
    .B(_01664_),
    .C(_01689_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _17531_ (.A(_01690_),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__xnor2_1 _17532_ (.A(_10520_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__nor2_1 _17533_ (.A(_10453_),
    .B(_10454_),
    .Y(_01694_));
 sky130_fd_sc_hd__a21o_1 _17534_ (.A1(_10447_),
    .A2(_10455_),
    .B1(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__or2b_1 _17535_ (.A(_10469_),
    .B_N(_10459_),
    .X(_01696_));
 sky130_fd_sc_hd__a21bo_1 _17536_ (.A1(_10463_),
    .A2(_10468_),
    .B1_N(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__buf_2 _17537_ (.A(_08555_),
    .X(_01698_));
 sky130_fd_sc_hd__or4_1 _17538_ (.A(_10203_),
    .B(_01698_),
    .C(_08395_),
    .D(_09080_),
    .X(_01699_));
 sky130_fd_sc_hd__buf_2 _17539_ (.A(_10203_),
    .X(_01700_));
 sky130_fd_sc_hd__o22ai_1 _17540_ (.A1(_01698_),
    .A2(_08395_),
    .B1(_09080_),
    .B2(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_1 _17541_ (.A(_01699_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__or3_1 _17542_ (.A(_08201_),
    .B(_08394_),
    .C(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__o21ai_1 _17543_ (.A1(_08201_),
    .A2(_08394_),
    .B1(_01702_),
    .Y(_01704_));
 sky130_fd_sc_hd__and2_1 _17544_ (.A(_01703_),
    .B(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__nor2_1 _17545_ (.A(_08856_),
    .B(_09696_),
    .Y(_01706_));
 sky130_fd_sc_hd__nor2_1 _17546_ (.A(_09671_),
    .B(_09697_),
    .Y(_01707_));
 sky130_fd_sc_hd__o22a_1 _17547_ (.A1(_09671_),
    .A2(_09696_),
    .B1(_09697_),
    .B2(_08856_),
    .X(_01708_));
 sky130_fd_sc_hd__a21oi_1 _17548_ (.A1(_01706_),
    .A2(_01707_),
    .B1(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__buf_2 _17549_ (.A(_09417_),
    .X(_01710_));
 sky130_fd_sc_hd__nor2_1 _17550_ (.A(_01710_),
    .B(_09326_),
    .Y(_01711_));
 sky130_fd_sc_hd__xnor2_1 _17551_ (.A(_01709_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__o31a_1 _17552_ (.A1(_01710_),
    .A2(_09198_),
    .A3(_10451_),
    .B1(_10449_),
    .X(_01713_));
 sky130_fd_sc_hd__xor2_1 _17553_ (.A(_01712_),
    .B(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__xnor2_1 _17554_ (.A(_01705_),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__xor2_1 _17555_ (.A(_01697_),
    .B(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__xnor2_1 _17556_ (.A(_01695_),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__or3_1 _17557_ (.A(_10228_),
    .B(_09697_),
    .C(_10466_),
    .X(_01718_));
 sky130_fd_sc_hd__a21bo_1 _17558_ (.A1(_10464_),
    .A2(_10465_),
    .B1_N(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__o31ai_1 _17559_ (.A1(_09700_),
    .A2(_10461_),
    .A3(_10475_),
    .B1(_10462_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor2_1 _17560_ (.A(_08858_),
    .B(_10104_),
    .Y(_01721_));
 sky130_fd_sc_hd__nor2_1 _17561_ (.A(_08868_),
    .B(_10460_),
    .Y(_01722_));
 sky130_fd_sc_hd__xnor2_1 _17562_ (.A(_01721_),
    .B(_01722_),
    .Y(_01723_));
 sky130_fd_sc_hd__nor2_1 _17563_ (.A(_10228_),
    .B(_09706_),
    .Y(_01724_));
 sky130_fd_sc_hd__xor2_1 _17564_ (.A(_01723_),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__xor2_1 _17565_ (.A(_01720_),
    .B(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__xnor2_1 _17566_ (.A(_01719_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__a21o_1 _17567_ (.A1(_10239_),
    .A2(_10477_),
    .B1(_10238_),
    .X(_01728_));
 sky130_fd_sc_hd__nor2_1 _17568_ (.A(_09700_),
    .B(_10473_),
    .Y(_01729_));
 sky130_fd_sc_hd__mux2_2 _17569_ (.A0(_09700_),
    .A1(_01729_),
    .S(_10475_),
    .X(_01730_));
 sky130_fd_sc_hd__xor2_1 _17570_ (.A(_10239_),
    .B(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__and2_1 _17571_ (.A(_01728_),
    .B(_01731_),
    .X(_01732_));
 sky130_fd_sc_hd__nor2_1 _17572_ (.A(_01728_),
    .B(_01731_),
    .Y(_01733_));
 sky130_fd_sc_hd__nor2_1 _17573_ (.A(_01732_),
    .B(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__xnor2_1 _17574_ (.A(_01727_),
    .B(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__nor2_1 _17575_ (.A(_10478_),
    .B(_10479_),
    .Y(_01736_));
 sky130_fd_sc_hd__a21oi_1 _17576_ (.A1(_10470_),
    .A2(_10480_),
    .B1(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__xor2_1 _17577_ (.A(_01735_),
    .B(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__xnor2_1 _17578_ (.A(_01717_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__and2b_1 _17579_ (.A_N(_10481_),
    .B(_10483_),
    .X(_01740_));
 sky130_fd_sc_hd__a21oi_1 _17580_ (.A1(_10458_),
    .A2(_10484_),
    .B1(_01740_),
    .Y(_01741_));
 sky130_fd_sc_hd__xor2_1 _17581_ (.A(_01739_),
    .B(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__xnor2_1 _17582_ (.A(_01693_),
    .B(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__a21oi_1 _17583_ (.A1(_10436_),
    .A2(_10490_),
    .B1(_10488_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _17584_ (.A(_01743_),
    .B(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__nand2_1 _17585_ (.A(_01743_),
    .B(_01744_),
    .Y(_01746_));
 sky130_fd_sc_hd__and2b_1 _17586_ (.A_N(_01745_),
    .B(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__xnor2_1 _17587_ (.A(_10519_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__o21a_1 _17588_ (.A1(_10491_),
    .A2(_10492_),
    .B1(_10494_),
    .X(_01749_));
 sky130_fd_sc_hd__xor2_1 _17589_ (.A(_01748_),
    .B(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__nand2_1 _17590_ (.A(_10402_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__or2_1 _17591_ (.A(_10402_),
    .B(_01750_),
    .X(_01752_));
 sky130_fd_sc_hd__nand2_2 _17592_ (.A(_01751_),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__o21a_1 _17593_ (.A1(_10496_),
    .A2(_10497_),
    .B1(_10499_),
    .X(_01754_));
 sky130_fd_sc_hd__xor2_4 _17594_ (.A(_01753_),
    .B(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__a21oi_1 _17595_ (.A1(_10378_),
    .A2(_10502_),
    .B1(_10503_),
    .Y(_01756_));
 sky130_fd_sc_hd__a41o_2 _17596_ (.A1(_10380_),
    .A2(_10385_),
    .A3(_10502_),
    .A4(_10504_),
    .B1(_01756_),
    .X(_01757_));
 sky130_fd_sc_hd__a21oi_1 _17597_ (.A1(_01755_),
    .A2(_01757_),
    .B1(_09938_),
    .Y(_01758_));
 sky130_fd_sc_hd__o21ai_4 _17598_ (.A1(_01755_),
    .A2(_01757_),
    .B1(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__nand2_1 _17599_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_01760_));
 sky130_fd_sc_hd__or2_1 _17600_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_01761_));
 sky130_fd_sc_hd__o211a_1 _17601_ (.A1(_10510_),
    .A2(_10513_),
    .B1(_01760_),
    .C1(_01761_),
    .X(_01762_));
 sky130_fd_sc_hd__a211oi_1 _17602_ (.A1(_01760_),
    .A2(_01761_),
    .B1(_10510_),
    .C1(_10513_),
    .Y(_01763_));
 sky130_fd_sc_hd__o31a_1 _17603_ (.A1(_10509_),
    .A2(_01762_),
    .A3(_01763_),
    .B1(_09945_),
    .X(_01764_));
 sky130_fd_sc_hd__o2bb2a_1 _17604_ (.A1_N(_01759_),
    .A2_N(_01764_),
    .B1(\rbzero.wall_tracer.trackDistX[4] ),
    .B2(_09946_),
    .X(_00543_));
 sky130_fd_sc_hd__nor2_1 _17605_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_01765_));
 sky130_fd_sc_hd__and2_1 _17606_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_01766_));
 sky130_fd_sc_hd__a21oi_1 _17607_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(\rbzero.wall_tracer.stepDistX[4] ),
    .B1(_01762_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor3_1 _17608_ (.A(_01765_),
    .B(_01766_),
    .C(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__o21a_1 _17609_ (.A1(_01765_),
    .A2(_01766_),
    .B1(_01767_),
    .X(_01769_));
 sky130_fd_sc_hd__or2_1 _17610_ (.A(_01748_),
    .B(_01749_),
    .X(_01770_));
 sky130_fd_sc_hd__or2b_1 _17611_ (.A(_01692_),
    .B_N(_10520_),
    .X(_01771_));
 sky130_fd_sc_hd__o2bb2a_1 _17612_ (.A1_N(_01671_),
    .A2_N(_01672_),
    .B1(_01669_),
    .B2(_01670_),
    .X(_01772_));
 sky130_fd_sc_hd__a21oi_1 _17613_ (.A1(_01690_),
    .A2(_01771_),
    .B1(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__and3_1 _17614_ (.A(_01690_),
    .B(_01771_),
    .C(_01772_),
    .X(_01774_));
 sky130_fd_sc_hd__nor2_1 _17615_ (.A(_01773_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21o_1 _17616_ (.A1(_01673_),
    .A2(_01688_),
    .B1(_01686_),
    .X(_01776_));
 sky130_fd_sc_hd__or2b_1 _17617_ (.A(_01715_),
    .B_N(_01697_),
    .X(_01777_));
 sky130_fd_sc_hd__or2b_1 _17618_ (.A(_01716_),
    .B_N(_01695_),
    .X(_01778_));
 sky130_fd_sc_hd__nor2_1 _17619_ (.A(_09793_),
    .B(_09503_),
    .Y(_01779_));
 sky130_fd_sc_hd__nor2_1 _17620_ (.A(_10208_),
    .B(_09378_),
    .Y(_01780_));
 sky130_fd_sc_hd__xnor2_1 _17621_ (.A(_01779_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__or2_1 _17622_ (.A(_09526_),
    .B(_09636_),
    .X(_01782_));
 sky130_fd_sc_hd__xnor2_1 _17623_ (.A(_01781_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__nand2_1 _17624_ (.A(_01665_),
    .B(_01666_),
    .Y(_01784_));
 sky130_fd_sc_hd__o31a_1 _17625_ (.A1(_09406_),
    .A2(_09637_),
    .A3(_01667_),
    .B1(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__xnor2_1 _17626_ (.A(_01783_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _17627_ (.A(_09406_),
    .B(_10030_),
    .Y(_01787_));
 sky130_fd_sc_hd__xor2_1 _17628_ (.A(_01786_),
    .B(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__o31ai_2 _17629_ (.A1(_10208_),
    .A2(_09511_),
    .A3(_01680_),
    .B1(_01678_),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_2 _17630_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08554_),
    .Y(_01790_));
 sky130_fd_sc_hd__or2_1 _17631_ (.A(_08360_),
    .B(_09132_),
    .X(_01791_));
 sky130_fd_sc_hd__or3_1 _17632_ (.A(_10205_),
    .B(_01790_),
    .C(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__o21ai_1 _17633_ (.A1(_10205_),
    .A2(_01790_),
    .B1(_01791_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _17634_ (.A(_01792_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _17635_ (.A(_10075_),
    .B(_09511_),
    .Y(_01795_));
 sky130_fd_sc_hd__xor2_1 _17636_ (.A(_01794_),
    .B(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__a21oi_1 _17637_ (.A1(_01699_),
    .A2(_01703_),
    .B1(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__and3_1 _17638_ (.A(_01699_),
    .B(_01703_),
    .C(_01796_),
    .X(_01798_));
 sky130_fd_sc_hd__nor2_1 _17639_ (.A(_01797_),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__xnor2_1 _17640_ (.A(_01789_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__a21oi_1 _17641_ (.A1(_10442_),
    .A2(_10444_),
    .B1(_01682_),
    .Y(_01801_));
 sky130_fd_sc_hd__a21oi_1 _17642_ (.A1(_01674_),
    .A2(_01683_),
    .B1(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _17643_ (.A(_01800_),
    .B(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__and2_1 _17644_ (.A(_01800_),
    .B(_01802_),
    .X(_01804_));
 sky130_fd_sc_hd__nor2_1 _17645_ (.A(_01803_),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__xnor2_1 _17646_ (.A(_01788_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__a21o_1 _17647_ (.A1(_01777_),
    .A2(_01778_),
    .B1(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__nand3_1 _17648_ (.A(_01777_),
    .B(_01778_),
    .C(_01806_),
    .Y(_01808_));
 sky130_fd_sc_hd__nand2_1 _17649_ (.A(_01807_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__xnor2_1 _17650_ (.A(_01776_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _17651_ (.A(_01712_),
    .B(_01713_),
    .Y(_01811_));
 sky130_fd_sc_hd__a21o_1 _17652_ (.A1(_01705_),
    .A2(_01714_),
    .B1(_01811_),
    .X(_01812_));
 sky130_fd_sc_hd__or2b_1 _17653_ (.A(_01725_),
    .B_N(_01720_),
    .X(_01813_));
 sky130_fd_sc_hd__or2b_1 _17654_ (.A(_01726_),
    .B_N(_01719_),
    .X(_01814_));
 sky130_fd_sc_hd__buf_2 _17655_ (.A(_09080_),
    .X(_01815_));
 sky130_fd_sc_hd__nand2_2 _17656_ (.A(_08292_),
    .B(_09077_),
    .Y(_01816_));
 sky130_fd_sc_hd__or4_1 _17657_ (.A(_01700_),
    .B(_01698_),
    .C(_01815_),
    .D(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__o22ai_1 _17658_ (.A1(_01698_),
    .A2(_01815_),
    .B1(_01816_),
    .B2(_01700_),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_1 _17659_ (.A(_01817_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__or3_1 _17660_ (.A(_08201_),
    .B(_08395_),
    .C(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__o21ai_1 _17661_ (.A1(_08201_),
    .A2(_08395_),
    .B1(_01819_),
    .Y(_01821_));
 sky130_fd_sc_hd__and2_1 _17662_ (.A(_01820_),
    .B(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__nor2_1 _17663_ (.A(_08856_),
    .B(_09706_),
    .Y(_01823_));
 sky130_fd_sc_hd__xnor2_1 _17664_ (.A(_01707_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _17665_ (.A(_09417_),
    .B(_09696_),
    .Y(_01825_));
 sky130_fd_sc_hd__xor2_1 _17666_ (.A(_01824_),
    .B(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__a22oi_1 _17667_ (.A1(_01706_),
    .A2(_01707_),
    .B1(_01709_),
    .B2(_01711_),
    .Y(_01827_));
 sky130_fd_sc_hd__nor2_1 _17668_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__and2_1 _17669_ (.A(_01826_),
    .B(_01827_),
    .X(_01829_));
 sky130_fd_sc_hd__nor2_1 _17670_ (.A(_01828_),
    .B(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__xnor2_1 _17671_ (.A(_01822_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__a21o_1 _17672_ (.A1(_01813_),
    .A2(_01814_),
    .B1(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__nand3_1 _17673_ (.A(_01813_),
    .B(_01814_),
    .C(_01831_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _17674_ (.A(_01832_),
    .B(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__xnor2_1 _17675_ (.A(_01812_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__or3_1 _17676_ (.A(_10228_),
    .B(_09706_),
    .C(_01723_),
    .X(_01836_));
 sky130_fd_sc_hd__a21bo_1 _17677_ (.A1(_01721_),
    .A2(_01722_),
    .B1_N(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__o21ai_4 _17678_ (.A1(_09700_),
    .A2(_10475_),
    .B1(_10462_),
    .Y(_01838_));
 sky130_fd_sc_hd__or3_1 _17679_ (.A(_08868_),
    .B(_08487_),
    .C(_10473_),
    .X(_01839_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17680_ (.A(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__o22ai_1 _17681_ (.A1(_08868_),
    .A2(_10473_),
    .B1(_10460_),
    .B2(_08858_),
    .Y(_01841_));
 sky130_fd_sc_hd__o21ai_1 _17682_ (.A1(_10461_),
    .A2(_01840_),
    .B1(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__nor2_1 _17683_ (.A(_10228_),
    .B(_10104_),
    .Y(_01843_));
 sky130_fd_sc_hd__xnor2_1 _17684_ (.A(_01842_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__xnor2_1 _17685_ (.A(_01838_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__xnor2_1 _17686_ (.A(_01837_),
    .B(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__nand2_1 _17687_ (.A(_10238_),
    .B(_01730_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand3b_1 _17688_ (.A_N(_01730_),
    .B(_10237_),
    .C(_10114_),
    .Y(_01848_));
 sky130_fd_sc_hd__and2_1 _17689_ (.A(_01847_),
    .B(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__buf_2 _17690_ (.A(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__xnor2_1 _17691_ (.A(_01846_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__a21oi_1 _17692_ (.A1(_01727_),
    .A2(_01734_),
    .B1(_01732_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _17693_ (.A(_01851_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__and2_1 _17694_ (.A(_01851_),
    .B(_01852_),
    .X(_01854_));
 sky130_fd_sc_hd__nor2_1 _17695_ (.A(_01853_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__xnor2_1 _17696_ (.A(_01835_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _17697_ (.A(_01735_),
    .B(_01737_),
    .Y(_01857_));
 sky130_fd_sc_hd__a21oi_1 _17698_ (.A1(_01717_),
    .A2(_01738_),
    .B1(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__xor2_1 _17699_ (.A(_01856_),
    .B(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__xnor2_1 _17700_ (.A(_01810_),
    .B(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor2_1 _17701_ (.A(_01739_),
    .B(_01741_),
    .Y(_01861_));
 sky130_fd_sc_hd__a21oi_1 _17702_ (.A1(_01693_),
    .A2(_01742_),
    .B1(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__xor2_1 _17703_ (.A(_01860_),
    .B(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(_01775_),
    .B(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21oi_1 _17705_ (.A1(_10519_),
    .A2(_01746_),
    .B1(_01745_),
    .Y(_01865_));
 sky130_fd_sc_hd__nor2_1 _17706_ (.A(_01864_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand2_1 _17707_ (.A(_01864_),
    .B(_01865_),
    .Y(_01867_));
 sky130_fd_sc_hd__and2b_1 _17708_ (.A_N(_01866_),
    .B(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__xnor2_1 _17709_ (.A(_10517_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__and3_1 _17710_ (.A(_01770_),
    .B(_01751_),
    .C(_01869_),
    .X(_01870_));
 sky130_fd_sc_hd__a21oi_1 _17711_ (.A1(_01770_),
    .A2(_01751_),
    .B1(_01869_),
    .Y(_01871_));
 sky130_fd_sc_hd__or2_1 _17712_ (.A(_01870_),
    .B(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__or2_1 _17713_ (.A(_01753_),
    .B(_01754_),
    .X(_01873_));
 sky130_fd_sc_hd__a21boi_2 _17714_ (.A1(_01755_),
    .A2(_01757_),
    .B1_N(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__a21oi_1 _17715_ (.A1(_01872_),
    .A2(_01874_),
    .B1(_09937_),
    .Y(_01875_));
 sky130_fd_sc_hd__o21ai_4 _17716_ (.A1(_01872_),
    .A2(_01874_),
    .B1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__o311a_1 _17717_ (.A1(_09954_),
    .A2(_01768_),
    .A3(_01769_),
    .B1(_09978_),
    .C1(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__a21oi_1 _17718_ (.A1(_06146_),
    .A2(_09920_),
    .B1(_01877_),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_1 _17719_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01878_));
 sky130_fd_sc_hd__and2_1 _17720_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .X(_01879_));
 sky130_fd_sc_hd__o21ba_1 _17721_ (.A1(_01765_),
    .A2(_01767_),
    .B1_N(_01766_),
    .X(_01880_));
 sky130_fd_sc_hd__o21ai_1 _17722_ (.A1(_01878_),
    .A2(_01879_),
    .B1(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__o31a_1 _17723_ (.A1(_01878_),
    .A2(_01879_),
    .A3(_01880_),
    .B1(_06095_),
    .X(_01882_));
 sky130_fd_sc_hd__or2b_1 _17724_ (.A(_01809_),
    .B_N(_01776_),
    .X(_01883_));
 sky130_fd_sc_hd__o22a_1 _17725_ (.A1(_01783_),
    .A2(_01785_),
    .B1(_01786_),
    .B2(_01787_),
    .X(_01884_));
 sky130_fd_sc_hd__a21oi_2 _17726_ (.A1(_01807_),
    .A2(_01883_),
    .B1(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__and3_1 _17727_ (.A(_01807_),
    .B(_01883_),
    .C(_01884_),
    .X(_01886_));
 sky130_fd_sc_hd__nor2_1 _17728_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__a21o_1 _17729_ (.A1(_01788_),
    .A2(_01805_),
    .B1(_01803_),
    .X(_01888_));
 sky130_fd_sc_hd__or2b_1 _17730_ (.A(_01834_),
    .B_N(_01812_),
    .X(_01889_));
 sky130_fd_sc_hd__o22a_1 _17731_ (.A1(_10075_),
    .A2(_09378_),
    .B1(_09503_),
    .B2(_10208_),
    .X(_01890_));
 sky130_fd_sc_hd__or4_1 _17732_ (.A(_10075_),
    .B(_10208_),
    .C(_09378_),
    .D(_09503_),
    .X(_01891_));
 sky130_fd_sc_hd__or2b_1 _17733_ (.A(_01890_),
    .B_N(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__or2_1 _17734_ (.A(_09793_),
    .B(_09768_),
    .X(_01893_));
 sky130_fd_sc_hd__xnor2_1 _17735_ (.A(_01892_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(_01779_),
    .B(_01780_),
    .Y(_01895_));
 sky130_fd_sc_hd__o31a_1 _17737_ (.A1(_09526_),
    .A2(_09768_),
    .A3(_01781_),
    .B1(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__xnor2_1 _17738_ (.A(_01894_),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_1 _17739_ (.A(_09526_),
    .B(_10030_),
    .Y(_01898_));
 sky130_fd_sc_hd__xor2_1 _17740_ (.A(_01897_),
    .B(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__a21bo_1 _17741_ (.A1(_01793_),
    .A2(_01795_),
    .B1_N(_01792_),
    .X(_01900_));
 sky130_fd_sc_hd__nand2_2 _17742_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08554_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _17743_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08391_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _17744_ (.A(_08360_),
    .B(_09225_),
    .Y(_01903_));
 sky130_fd_sc_hd__a31o_1 _17745_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_08554_),
    .A3(_08391_),
    .B1(_01903_),
    .X(_01904_));
 sky130_fd_sc_hd__o21ai_1 _17746_ (.A1(_01791_),
    .A2(_01902_),
    .B1(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__or3_1 _17747_ (.A(_10205_),
    .B(_01901_),
    .C(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__o21ai_1 _17748_ (.A1(_10205_),
    .A2(_01901_),
    .B1(_01905_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _17749_ (.A(_01906_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__a21oi_1 _17750_ (.A1(_01817_),
    .A2(_01820_),
    .B1(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__and3_1 _17751_ (.A(_01817_),
    .B(_01820_),
    .C(_01908_),
    .X(_01910_));
 sky130_fd_sc_hd__nor2_1 _17752_ (.A(_01909_),
    .B(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__xnor2_1 _17753_ (.A(_01900_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__a21oi_1 _17754_ (.A1(_01789_),
    .A2(_01799_),
    .B1(_01797_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _17755_ (.A(_01912_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__and2_1 _17756_ (.A(_01912_),
    .B(_01913_),
    .X(_01915_));
 sky130_fd_sc_hd__nor2_1 _17757_ (.A(_01914_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_1 _17758_ (.A(_01899_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__a21o_1 _17759_ (.A1(_01832_),
    .A2(_01889_),
    .B1(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__nand3_1 _17760_ (.A(_01832_),
    .B(_01889_),
    .C(_01917_),
    .Y(_01919_));
 sky130_fd_sc_hd__nand2_1 _17761_ (.A(_01918_),
    .B(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__xnor2_1 _17762_ (.A(_01888_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__a21o_1 _17763_ (.A1(_01822_),
    .A2(_01830_),
    .B1(_01828_),
    .X(_01922_));
 sky130_fd_sc_hd__nand2_1 _17764_ (.A(_01838_),
    .B(_01844_),
    .Y(_01923_));
 sky130_fd_sc_hd__or2b_1 _17765_ (.A(_01845_),
    .B_N(_01837_),
    .X(_01924_));
 sky130_fd_sc_hd__or4_1 _17766_ (.A(_01700_),
    .B(_01698_),
    .C(_01816_),
    .D(_09446_),
    .X(_01925_));
 sky130_fd_sc_hd__a2bb2o_1 _17767_ (.A1_N(_01700_),
    .A2_N(_09446_),
    .B1(_09077_),
    .B2(_08556_),
    .X(_01926_));
 sky130_fd_sc_hd__nand2_1 _17768_ (.A(_01925_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__or3_1 _17769_ (.A(_01815_),
    .B(_10445_),
    .C(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__o21ai_1 _17770_ (.A1(_01815_),
    .A2(_10445_),
    .B1(_01927_),
    .Y(_01929_));
 sky130_fd_sc_hd__and2_1 _17771_ (.A(_01928_),
    .B(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__nor2_1 _17772_ (.A(_09671_),
    .B(_10104_),
    .Y(_01931_));
 sky130_fd_sc_hd__o22a_1 _17773_ (.A1(_09671_),
    .A2(_09706_),
    .B1(_10104_),
    .B2(_08856_),
    .X(_01932_));
 sky130_fd_sc_hd__a21o_1 _17774_ (.A1(_01823_),
    .A2(_01931_),
    .B1(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__nor2_1 _17775_ (.A(_01710_),
    .B(_09697_),
    .Y(_01934_));
 sky130_fd_sc_hd__xor2_1 _17776_ (.A(_01933_),
    .B(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__nand2_1 _17777_ (.A(_01707_),
    .B(_01823_),
    .Y(_01936_));
 sky130_fd_sc_hd__o31a_1 _17778_ (.A1(_01710_),
    .A2(_09696_),
    .A3(_01824_),
    .B1(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__nor2_1 _17779_ (.A(_01935_),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__and2_1 _17780_ (.A(_01935_),
    .B(_01937_),
    .X(_01939_));
 sky130_fd_sc_hd__nor2_1 _17781_ (.A(_01938_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__xnor2_1 _17782_ (.A(_01930_),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__a21o_1 _17783_ (.A1(_01923_),
    .A2(_01924_),
    .B1(_01941_),
    .X(_01942_));
 sky130_fd_sc_hd__nand3_1 _17784_ (.A(_01923_),
    .B(_01924_),
    .C(_01941_),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_1 _17785_ (.A(_01942_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__xnor2_1 _17786_ (.A(_01922_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__a2bb2o_1 _17787_ (.A1_N(_10461_),
    .A2_N(_01840_),
    .B1(_01843_),
    .B2(_01841_),
    .X(_01946_));
 sky130_fd_sc_hd__a21oi_1 _17788_ (.A1(_08868_),
    .A2(_08858_),
    .B1(_10473_),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _17789_ (.A(_01840_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_1 _17790_ (.A(_10228_),
    .B(_10461_),
    .Y(_01949_));
 sky130_fd_sc_hd__xnor2_1 _17791_ (.A(_01948_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__xor2_1 _17792_ (.A(_01838_),
    .B(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__nand2_1 _17793_ (.A(_01946_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__or2_1 _17794_ (.A(_01946_),
    .B(_01951_),
    .X(_01953_));
 sky130_fd_sc_hd__and2_1 _17795_ (.A(_01952_),
    .B(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__xnor2_1 _17796_ (.A(_01850_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__a21boi_1 _17797_ (.A1(_01846_),
    .A2(_01850_),
    .B1_N(_01847_),
    .Y(_01956_));
 sky130_fd_sc_hd__nor2_1 _17798_ (.A(_01955_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__and2_1 _17799_ (.A(_01955_),
    .B(_01956_),
    .X(_01958_));
 sky130_fd_sc_hd__nor2_1 _17800_ (.A(_01957_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__xnor2_1 _17801_ (.A(_01945_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__a21oi_1 _17802_ (.A1(_01835_),
    .A2(_01855_),
    .B1(_01853_),
    .Y(_01961_));
 sky130_fd_sc_hd__xor2_1 _17803_ (.A(_01960_),
    .B(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__xnor2_1 _17804_ (.A(_01921_),
    .B(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__nor2_1 _17805_ (.A(_01856_),
    .B(_01858_),
    .Y(_01964_));
 sky130_fd_sc_hd__a21oi_1 _17806_ (.A1(_01810_),
    .A2(_01859_),
    .B1(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__xor2_1 _17807_ (.A(_01963_),
    .B(_01965_),
    .X(_01966_));
 sky130_fd_sc_hd__xnor2_1 _17808_ (.A(_01887_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _17809_ (.A(_01860_),
    .B(_01862_),
    .Y(_01968_));
 sky130_fd_sc_hd__a21oi_1 _17810_ (.A1(_01775_),
    .A2(_01863_),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__or2_1 _17811_ (.A(_01967_),
    .B(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_1 _17812_ (.A(_01967_),
    .B(_01969_),
    .Y(_01971_));
 sky130_fd_sc_hd__and2_1 _17813_ (.A(_01970_),
    .B(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__nand2_1 _17814_ (.A(_01773_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__or2_1 _17815_ (.A(_01773_),
    .B(_01972_),
    .X(_01974_));
 sky130_fd_sc_hd__nand2_1 _17816_ (.A(_01973_),
    .B(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__a21oi_1 _17817_ (.A1(_10517_),
    .A2(_01867_),
    .B1(_01866_),
    .Y(_01976_));
 sky130_fd_sc_hd__or2_2 _17818_ (.A(_01975_),
    .B(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__nand2_1 _17819_ (.A(_01975_),
    .B(_01976_),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _17820_ (.A(_01977_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__or3b_1 _17821_ (.A(_01870_),
    .B(_01871_),
    .C_N(_01755_),
    .X(_01980_));
 sky130_fd_sc_hd__or2b_1 _17822_ (.A(_01980_),
    .B_N(_01756_),
    .X(_01981_));
 sky130_fd_sc_hd__o41a_1 _17823_ (.A1(_10387_),
    .A2(_10388_),
    .A3(_10505_),
    .A4(_01980_),
    .B1(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__o21ba_1 _17824_ (.A1(_01873_),
    .A2(_01870_),
    .B1_N(_01871_),
    .X(_01983_));
 sky130_fd_sc_hd__and3_1 _17825_ (.A(_01979_),
    .B(_01982_),
    .C(_01983_),
    .X(_01984_));
 sky130_fd_sc_hd__a21o_2 _17826_ (.A1(_01982_),
    .A2(_01983_),
    .B1(_01979_),
    .X(_01985_));
 sky130_fd_sc_hd__or3b_1 _17827_ (.A(_06094_),
    .B(_01984_),
    .C_N(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__a21bo_1 _17828_ (.A1(_01881_),
    .A2(_01882_),
    .B1_N(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _17829_ (.A0(\rbzero.wall_tracer.trackDistX[6] ),
    .A1(_01987_),
    .S(_09978_),
    .X(_01988_));
 sky130_fd_sc_hd__clkbuf_1 _17830_ (.A(_01988_),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _17831_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_1 _17832_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_01990_));
 sky130_fd_sc_hd__or2b_1 _17833_ (.A(_01989_),
    .B_N(_01990_),
    .X(_01991_));
 sky130_fd_sc_hd__o21ba_1 _17834_ (.A1(_01878_),
    .A2(_01880_),
    .B1_N(_01879_),
    .X(_01992_));
 sky130_fd_sc_hd__xnor2_1 _17835_ (.A(_01991_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__or2b_1 _17836_ (.A(_01920_),
    .B_N(_01888_),
    .X(_01994_));
 sky130_fd_sc_hd__o22a_1 _17837_ (.A1(_01894_),
    .A2(_01896_),
    .B1(_01897_),
    .B2(_01898_),
    .X(_01995_));
 sky130_fd_sc_hd__a21oi_2 _17838_ (.A1(_01918_),
    .A2(_01994_),
    .B1(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__and3_1 _17839_ (.A(_01918_),
    .B(_01994_),
    .C(_01995_),
    .X(_01997_));
 sky130_fd_sc_hd__nor2_1 _17840_ (.A(_01996_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__a21o_1 _17841_ (.A1(_01899_),
    .A2(_01916_),
    .B1(_01914_),
    .X(_01999_));
 sky130_fd_sc_hd__or2b_1 _17842_ (.A(_01944_),
    .B_N(_01922_),
    .X(_02000_));
 sky130_fd_sc_hd__and3_1 _17843_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08543_),
    .C(_08323_),
    .X(_02001_));
 sky130_fd_sc_hd__nand2_1 _17844_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08554_),
    .Y(_02002_));
 sky130_fd_sc_hd__nor2_1 _17845_ (.A(_10205_),
    .B(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _17846_ (.A(_02001_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__or2_1 _17847_ (.A(_02001_),
    .B(_02003_),
    .X(_02005_));
 sky130_fd_sc_hd__nand2_1 _17848_ (.A(_02004_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(_10208_),
    .B(_09768_),
    .Y(_02007_));
 sky130_fd_sc_hd__xor2_1 _17850_ (.A(_02006_),
    .B(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__o31a_1 _17851_ (.A1(_09793_),
    .A2(_09768_),
    .A3(_01890_),
    .B1(_01891_),
    .X(_02009_));
 sky130_fd_sc_hd__xor2_1 _17852_ (.A(_02008_),
    .B(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__and2_1 _17853_ (.A(_09793_),
    .B(_10030_),
    .X(_02011_));
 sky130_fd_sc_hd__xor2_1 _17854_ (.A(_02010_),
    .B(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__o21ai_1 _17855_ (.A1(_01791_),
    .A2(_01902_),
    .B1(_01906_),
    .Y(_02013_));
 sky130_fd_sc_hd__or3_1 _17856_ (.A(_01815_),
    .B(_01676_),
    .C(_01902_),
    .X(_02014_));
 sky130_fd_sc_hd__o21ai_1 _17857_ (.A1(_01815_),
    .A2(_01676_),
    .B1(_01902_),
    .Y(_02015_));
 sky130_fd_sc_hd__and2_1 _17858_ (.A(_02014_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__nor2_1 _17859_ (.A(_08360_),
    .B(_09511_),
    .Y(_02017_));
 sky130_fd_sc_hd__xnor2_1 _17860_ (.A(_02016_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__a21oi_1 _17861_ (.A1(_01925_),
    .A2(_01928_),
    .B1(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__and3_1 _17862_ (.A(_01925_),
    .B(_01928_),
    .C(_02018_),
    .X(_02020_));
 sky130_fd_sc_hd__nor2_1 _17863_ (.A(_02019_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__xnor2_1 _17864_ (.A(_02013_),
    .B(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__a21oi_1 _17865_ (.A1(_01900_),
    .A2(_01911_),
    .B1(_01909_),
    .Y(_02023_));
 sky130_fd_sc_hd__nor2_1 _17866_ (.A(_02022_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__and2_1 _17867_ (.A(_02022_),
    .B(_02023_),
    .X(_02025_));
 sky130_fd_sc_hd__nor2_1 _17868_ (.A(_02024_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__xnor2_1 _17869_ (.A(_02012_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__a21o_1 _17870_ (.A1(_01942_),
    .A2(_02000_),
    .B1(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__nand3_1 _17871_ (.A(_01942_),
    .B(_02000_),
    .C(_02027_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand2_1 _17872_ (.A(_02028_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__xnor2_1 _17873_ (.A(_01999_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__or2_1 _17874_ (.A(_10228_),
    .B(_01948_),
    .X(_02032_));
 sky130_fd_sc_hd__or2_1 _17875_ (.A(_10461_),
    .B(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__nor2_1 _17876_ (.A(_10228_),
    .B(_10473_),
    .Y(_02034_));
 sky130_fd_sc_hd__mux2_1 _17877_ (.A0(_10228_),
    .A1(_02034_),
    .S(_01948_),
    .X(_02035_));
 sky130_fd_sc_hd__xnor2_2 _17878_ (.A(_01838_),
    .B(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__a21o_1 _17879_ (.A1(_01840_),
    .A2(_02033_),
    .B1(_02036_),
    .X(_02037_));
 sky130_fd_sc_hd__nand3_1 _17880_ (.A(_01840_),
    .B(_02033_),
    .C(_02036_),
    .Y(_02038_));
 sky130_fd_sc_hd__and2_1 _17881_ (.A(_02037_),
    .B(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__xnor2_1 _17882_ (.A(_01850_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__a21boi_1 _17883_ (.A1(_01850_),
    .A2(_01954_),
    .B1_N(_01847_),
    .Y(_02041_));
 sky130_fd_sc_hd__nor2_1 _17884_ (.A(_02040_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__and2_1 _17885_ (.A(_02040_),
    .B(_02041_),
    .X(_02043_));
 sky130_fd_sc_hd__nor2_1 _17886_ (.A(_02042_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__a21o_1 _17887_ (.A1(_01930_),
    .A2(_01940_),
    .B1(_01938_),
    .X(_02045_));
 sky130_fd_sc_hd__nand2_1 _17888_ (.A(_01838_),
    .B(_01950_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_1 _17889_ (.A(_01700_),
    .B(_09565_),
    .Y(_02047_));
 sky130_fd_sc_hd__nor2_1 _17890_ (.A(_01698_),
    .B(_09446_),
    .Y(_02048_));
 sky130_fd_sc_hd__xnor2_1 _17891_ (.A(_02047_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__or3_1 _17892_ (.A(_01816_),
    .B(_10445_),
    .C(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__o21ai_1 _17893_ (.A1(_01816_),
    .A2(_10445_),
    .B1(_02049_),
    .Y(_02051_));
 sky130_fd_sc_hd__and2_1 _17894_ (.A(_02050_),
    .B(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__nor2_1 _17895_ (.A(_08856_),
    .B(_10461_),
    .Y(_02053_));
 sky130_fd_sc_hd__xnor2_1 _17896_ (.A(_01931_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _17897_ (.A(_01710_),
    .B(_09706_),
    .Y(_02055_));
 sky130_fd_sc_hd__xor2_1 _17898_ (.A(_02054_),
    .B(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _17899_ (.A(_01823_),
    .B(_01931_),
    .Y(_02057_));
 sky130_fd_sc_hd__o31a_1 _17900_ (.A1(_01710_),
    .A2(_09697_),
    .A3(_01933_),
    .B1(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__xor2_1 _17901_ (.A(_02056_),
    .B(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__xnor2_1 _17902_ (.A(_02052_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__a21o_1 _17903_ (.A1(_02046_),
    .A2(_01952_),
    .B1(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__nand3_1 _17904_ (.A(_02046_),
    .B(_01952_),
    .C(_02060_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _17905_ (.A(_02061_),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__xnor2_1 _17906_ (.A(_02045_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__xnor2_1 _17907_ (.A(_02044_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__a21oi_1 _17908_ (.A1(_01945_),
    .A2(_01959_),
    .B1(_01957_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _17909_ (.A(_02065_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__and2_1 _17910_ (.A(_02065_),
    .B(_02066_),
    .X(_02068_));
 sky130_fd_sc_hd__nor2_1 _17911_ (.A(_02067_),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__xnor2_1 _17912_ (.A(_02031_),
    .B(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_1 _17913_ (.A(_01960_),
    .B(_01961_),
    .Y(_02071_));
 sky130_fd_sc_hd__a21oi_1 _17914_ (.A1(_01921_),
    .A2(_01962_),
    .B1(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__xor2_1 _17915_ (.A(_02070_),
    .B(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__xnor2_1 _17916_ (.A(_01998_),
    .B(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__nor2_1 _17917_ (.A(_01963_),
    .B(_01965_),
    .Y(_02075_));
 sky130_fd_sc_hd__a21oi_1 _17918_ (.A1(_01887_),
    .A2(_01966_),
    .B1(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__nor2_1 _17919_ (.A(_02074_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__and2_1 _17920_ (.A(_02074_),
    .B(_02076_),
    .X(_02078_));
 sky130_fd_sc_hd__nor2_1 _17921_ (.A(_02077_),
    .B(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _17922_ (.A(_01885_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__a21o_2 _17923_ (.A1(_01970_),
    .A2(_01973_),
    .B1(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__and3_2 _17924_ (.A(_01970_),
    .B(_01973_),
    .C(_02080_),
    .X(_02082_));
 sky130_fd_sc_hd__inv_2 _17925_ (.A(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _17926_ (.A(_02081_),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__a21oi_1 _17927_ (.A1(_01977_),
    .A2(_01985_),
    .B1(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__a31o_1 _17928_ (.A1(_01977_),
    .A2(_01985_),
    .A3(_02084_),
    .B1(_06094_),
    .X(_02086_));
 sky130_fd_sc_hd__or2_1 _17929_ (.A(_02085_),
    .B(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__o211a_1 _17930_ (.A1(_09954_),
    .A2(_01993_),
    .B1(_02087_),
    .C1(_09945_),
    .X(_02088_));
 sky130_fd_sc_hd__a21oi_1 _17931_ (.A1(_06143_),
    .A2(_09919_),
    .B1(_02088_),
    .Y(_00546_));
 sky130_fd_sc_hd__or2b_1 _17932_ (.A(_02030_),
    .B_N(_01999_),
    .X(_02089_));
 sky130_fd_sc_hd__o2bb2a_1 _17933_ (.A1_N(_02010_),
    .A2_N(_02011_),
    .B1(_02008_),
    .B2(_02009_),
    .X(_02090_));
 sky130_fd_sc_hd__a21oi_2 _17934_ (.A1(_02028_),
    .A2(_02089_),
    .B1(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__and3_1 _17935_ (.A(_02028_),
    .B(_02089_),
    .C(_02090_),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_1 _17936_ (.A(_02091_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__a21bo_1 _17937_ (.A1(_01850_),
    .A2(_02039_),
    .B1_N(_01847_),
    .X(_02094_));
 sky130_fd_sc_hd__nand2_1 _17938_ (.A(_01840_),
    .B(_02032_),
    .Y(_02095_));
 sky130_fd_sc_hd__xnor2_2 _17939_ (.A(_02036_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__xor2_1 _17940_ (.A(_01850_),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__and2_1 _17941_ (.A(_02094_),
    .B(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__nor2_1 _17942_ (.A(_02094_),
    .B(_02097_),
    .Y(_02099_));
 sky130_fd_sc_hd__nor2_1 _17943_ (.A(_02098_),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_1 _17944_ (.A(_02056_),
    .B(_02058_),
    .Y(_02101_));
 sky130_fd_sc_hd__a21o_1 _17945_ (.A1(_02052_),
    .A2(_02059_),
    .B1(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__nand2_1 _17946_ (.A(_01838_),
    .B(_02035_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_1 _17947_ (.A(_02103_),
    .B(_02037_),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _17948_ (.A(_01698_),
    .B(_09703_),
    .Y(_02105_));
 sky130_fd_sc_hd__o22a_1 _17949_ (.A1(_01698_),
    .A2(_09565_),
    .B1(_09703_),
    .B2(_01700_),
    .X(_02106_));
 sky130_fd_sc_hd__a21o_1 _17950_ (.A1(_02047_),
    .A2(_02105_),
    .B1(_02106_),
    .X(_02107_));
 sky130_fd_sc_hd__or3_1 _17951_ (.A(_10445_),
    .B(_09446_),
    .C(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__o21ai_1 _17952_ (.A1(_10445_),
    .A2(_09446_),
    .B1(_02107_),
    .Y(_02109_));
 sky130_fd_sc_hd__and2_1 _17953_ (.A(_02108_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__nand2_1 _17954_ (.A(_10115_),
    .B(_10116_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor3_1 _17955_ (.A(_08856_),
    .B(_09671_),
    .C(_10473_),
    .Y(_02112_));
 sky130_fd_sc_hd__o22a_1 _17956_ (.A1(_08856_),
    .A2(_10473_),
    .B1(_10461_),
    .B2(_09671_),
    .X(_02113_));
 sky130_fd_sc_hd__a21oi_1 _17957_ (.A1(_02111_),
    .A2(_02112_),
    .B1(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _17958_ (.A(_01710_),
    .B(_10104_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _17959_ (.A(_02114_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__or2_1 _17960_ (.A(_02114_),
    .B(_02115_),
    .X(_02117_));
 sky130_fd_sc_hd__nand2_1 _17961_ (.A(_02116_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__nand2_1 _17962_ (.A(_01931_),
    .B(_02053_),
    .Y(_02119_));
 sky130_fd_sc_hd__o31a_1 _17963_ (.A1(_01710_),
    .A2(_09706_),
    .A3(_02054_),
    .B1(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__nor2_1 _17964_ (.A(_02118_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__and2_1 _17965_ (.A(_02118_),
    .B(_02120_),
    .X(_02122_));
 sky130_fd_sc_hd__nor2_1 _17966_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__xor2_1 _17967_ (.A(_02110_),
    .B(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__xnor2_1 _17968_ (.A(_02104_),
    .B(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__xnor2_1 _17969_ (.A(_02102_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__xnor2_1 _17970_ (.A(_02100_),
    .B(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__a21oi_1 _17971_ (.A1(_02044_),
    .A2(_02064_),
    .B1(_02042_),
    .Y(_02128_));
 sky130_fd_sc_hd__xor2_1 _17972_ (.A(_02127_),
    .B(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__a21o_1 _17973_ (.A1(_02012_),
    .A2(_02026_),
    .B1(_02024_),
    .X(_02130_));
 sky130_fd_sc_hd__or2b_1 _17974_ (.A(_02063_),
    .B_N(_02045_),
    .X(_02131_));
 sky130_fd_sc_hd__or2_2 _17975_ (.A(_08360_),
    .B(_09378_),
    .X(_02132_));
 sky130_fd_sc_hd__or2b_1 _17976_ (.A(_09503_),
    .B_N(_08303_),
    .X(_02133_));
 sky130_fd_sc_hd__xnor2_2 _17977_ (.A(_02132_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__nor2_1 _17978_ (.A(_10075_),
    .B(_09637_),
    .Y(_02135_));
 sky130_fd_sc_hd__xor2_2 _17979_ (.A(_02134_),
    .B(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__o31a_1 _17980_ (.A1(_10208_),
    .A2(_09768_),
    .A3(_02006_),
    .B1(_02004_),
    .X(_02137_));
 sky130_fd_sc_hd__xor2_2 _17981_ (.A(_02136_),
    .B(_02137_),
    .X(_02138_));
 sky130_fd_sc_hd__and2_1 _17982_ (.A(_10208_),
    .B(_10030_),
    .X(_02139_));
 sky130_fd_sc_hd__xor2_2 _17983_ (.A(_02138_),
    .B(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__a21bo_1 _17984_ (.A1(_02016_),
    .A2(_02017_),
    .B1_N(_02014_),
    .X(_02141_));
 sky130_fd_sc_hd__nand2_1 _17985_ (.A(_02047_),
    .B(_02048_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _17986_ (.A(_01815_),
    .B(_01790_),
    .Y(_02143_));
 sky130_fd_sc_hd__nor2_1 _17987_ (.A(_01816_),
    .B(_01676_),
    .Y(_02144_));
 sky130_fd_sc_hd__xnor2_1 _17988_ (.A(_02143_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__or3_1 _17989_ (.A(_08395_),
    .B(_01901_),
    .C(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__o21ai_1 _17990_ (.A1(_08395_),
    .A2(_01901_),
    .B1(_02145_),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_1 _17991_ (.A(_02146_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__a21o_1 _17992_ (.A1(_02142_),
    .A2(_02050_),
    .B1(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__nand3_1 _17993_ (.A(_02142_),
    .B(_02050_),
    .C(_02148_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_1 _17994_ (.A(_02149_),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__xor2_1 _17995_ (.A(_02141_),
    .B(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__a21oi_1 _17996_ (.A1(_02013_),
    .A2(_02021_),
    .B1(_02019_),
    .Y(_02153_));
 sky130_fd_sc_hd__nor2_1 _17997_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__and2_1 _17998_ (.A(_02152_),
    .B(_02153_),
    .X(_02155_));
 sky130_fd_sc_hd__nor2_1 _17999_ (.A(_02154_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__xnor2_1 _18000_ (.A(_02140_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__a21oi_1 _18001_ (.A1(_02061_),
    .A2(_02131_),
    .B1(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__and3_1 _18002_ (.A(_02061_),
    .B(_02131_),
    .C(_02157_),
    .X(_02159_));
 sky130_fd_sc_hd__or2_1 _18003_ (.A(_02158_),
    .B(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_02130_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__nand2_1 _18005_ (.A(_02129_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__or2_1 _18006_ (.A(_02129_),
    .B(_02161_),
    .X(_02163_));
 sky130_fd_sc_hd__nand2_1 _18007_ (.A(_02162_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_1 _18008_ (.A1(_02031_),
    .A2(_02069_),
    .B1(_02067_),
    .Y(_02165_));
 sky130_fd_sc_hd__xor2_1 _18009_ (.A(_02164_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__nand2_1 _18010_ (.A(_02093_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__or2_1 _18011_ (.A(_02093_),
    .B(_02166_),
    .X(_02168_));
 sky130_fd_sc_hd__nand2_1 _18012_ (.A(_02167_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__nor2_1 _18013_ (.A(_02070_),
    .B(_02072_),
    .Y(_02170_));
 sky130_fd_sc_hd__a21oi_2 _18014_ (.A1(_01998_),
    .A2(_02073_),
    .B1(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__xor2_1 _18015_ (.A(_02169_),
    .B(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__xnor2_1 _18016_ (.A(_01996_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__a21oi_2 _18017_ (.A1(_01885_),
    .A2(_02079_),
    .B1(_02077_),
    .Y(_02174_));
 sky130_fd_sc_hd__or2_1 _18018_ (.A(_02173_),
    .B(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__nand2_1 _18019_ (.A(_02173_),
    .B(_02174_),
    .Y(_02176_));
 sky130_fd_sc_hd__and2_1 _18020_ (.A(_02175_),
    .B(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__inv_2 _18021_ (.A(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__a311o_1 _18022_ (.A1(_01977_),
    .A2(_01985_),
    .A3(_02081_),
    .B1(_02082_),
    .C1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__a31o_1 _18023_ (.A1(_01977_),
    .A2(_01985_),
    .A3(_02081_),
    .B1(_02082_),
    .X(_02180_));
 sky130_fd_sc_hd__a21oi_1 _18024_ (.A1(_02178_),
    .A2(_02180_),
    .B1(_09938_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _18025_ (.A(_02179_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_1 _18026_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .X(_02183_));
 sky130_fd_sc_hd__nand2_1 _18027_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _18028_ (.A(_02183_),
    .B(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__o21a_1 _18029_ (.A1(_01989_),
    .A2(_01992_),
    .B1(_01990_),
    .X(_02186_));
 sky130_fd_sc_hd__or2_1 _18030_ (.A(_02185_),
    .B(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__a21oi_1 _18031_ (.A1(_02185_),
    .A2(_02186_),
    .B1(_10509_),
    .Y(_02188_));
 sky130_fd_sc_hd__a21oi_1 _18032_ (.A1(_02187_),
    .A2(_02188_),
    .B1(_09919_),
    .Y(_02189_));
 sky130_fd_sc_hd__o2bb2a_1 _18033_ (.A1_N(_02182_),
    .A2_N(_02189_),
    .B1(\rbzero.wall_tracer.trackDistX[8] ),
    .B2(_09946_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _18034_ (.A(_02169_),
    .B(_02171_),
    .X(_02190_));
 sky130_fd_sc_hd__nand2_1 _18035_ (.A(_01996_),
    .B(_02172_),
    .Y(_02191_));
 sky130_fd_sc_hd__a21o_1 _18036_ (.A1(_02100_),
    .A2(_02126_),
    .B1(_02098_),
    .X(_02192_));
 sky130_fd_sc_hd__a21o_1 _18037_ (.A1(_02110_),
    .A2(_02123_),
    .B1(_02121_),
    .X(_02193_));
 sky130_fd_sc_hd__or2b_1 _18038_ (.A(_02036_),
    .B_N(_02095_),
    .X(_02194_));
 sky130_fd_sc_hd__nand2_1 _18039_ (.A(_02103_),
    .B(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _18040_ (.A(_08292_),
    .B(_09572_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _18041_ (.A(_01700_),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__xnor2_1 _18042_ (.A(_02105_),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _18043_ (.A(_10445_),
    .B(_09565_),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _18044_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__nand2_1 _18045_ (.A(_02111_),
    .B(_02112_),
    .Y(_02201_));
 sky130_fd_sc_hd__a21oi_1 _18046_ (.A1(_08856_),
    .A2(_09671_),
    .B1(_10473_),
    .Y(_02202_));
 sky130_fd_sc_hd__or2b_1 _18047_ (.A(_02112_),
    .B_N(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__or2_1 _18048_ (.A(_01710_),
    .B(_10461_),
    .X(_02204_));
 sky130_fd_sc_hd__xnor2_1 _18049_ (.A(_02203_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__a21oi_1 _18050_ (.A1(_02201_),
    .A2(_02116_),
    .B1(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__and3_1 _18051_ (.A(_02201_),
    .B(_02116_),
    .C(_02205_),
    .X(_02207_));
 sky130_fd_sc_hd__nor2_1 _18052_ (.A(_02206_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__xor2_1 _18053_ (.A(_02200_),
    .B(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__and2_1 _18054_ (.A(_02195_),
    .B(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__nor2_1 _18055_ (.A(_02195_),
    .B(_02209_),
    .Y(_02211_));
 sky130_fd_sc_hd__nor2_1 _18056_ (.A(_02210_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__xnor2_1 _18057_ (.A(_02193_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__mux2_1 _18058_ (.A0(_01848_),
    .A1(_01847_),
    .S(_02096_),
    .X(_02214_));
 sky130_fd_sc_hd__xnor2_1 _18059_ (.A(_02213_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__xnor2_1 _18060_ (.A(_02192_),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__a21o_1 _18061_ (.A1(_02140_),
    .A2(_02156_),
    .B1(_02154_),
    .X(_02217_));
 sky130_fd_sc_hd__or2b_1 _18062_ (.A(_02125_),
    .B_N(_02102_),
    .X(_02218_));
 sky130_fd_sc_hd__a21bo_1 _18063_ (.A1(_02104_),
    .A2(_02124_),
    .B1_N(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__a22o_1 _18064_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_08389_),
    .B1(_08391_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_02220_));
 sky130_fd_sc_hd__nand2_1 _18065_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08391_),
    .Y(_02221_));
 sky130_fd_sc_hd__or2_1 _18066_ (.A(_02132_),
    .B(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__nand2_1 _18067_ (.A(_02220_),
    .B(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__or2b_1 _18068_ (.A(_09768_),
    .B_N(_08303_),
    .X(_02224_));
 sky130_fd_sc_hd__xnor2_2 _18069_ (.A(_02223_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__or2_1 _18070_ (.A(_02132_),
    .B(_02133_),
    .X(_02226_));
 sky130_fd_sc_hd__o31a_1 _18071_ (.A1(_10075_),
    .A2(_09768_),
    .A3(_02134_),
    .B1(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__xor2_2 _18072_ (.A(_02225_),
    .B(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__and2_1 _18073_ (.A(_10075_),
    .B(_10030_),
    .X(_02229_));
 sky130_fd_sc_hd__xor2_2 _18074_ (.A(_02228_),
    .B(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__or2b_1 _18075_ (.A(_02151_),
    .B_N(_02141_),
    .X(_02231_));
 sky130_fd_sc_hd__a21bo_1 _18076_ (.A1(_02143_),
    .A2(_02144_),
    .B1_N(_02146_),
    .X(_02232_));
 sky130_fd_sc_hd__a21bo_1 _18077_ (.A1(_02047_),
    .A2(_02105_),
    .B1_N(_02108_),
    .X(_02233_));
 sky130_fd_sc_hd__or4_1 _18078_ (.A(_01816_),
    .B(_01676_),
    .C(_09446_),
    .D(_01790_),
    .X(_02234_));
 sky130_fd_sc_hd__o22ai_1 _18079_ (.A1(_01676_),
    .A2(_09446_),
    .B1(_01790_),
    .B2(_01816_),
    .Y(_02235_));
 sky130_fd_sc_hd__nand2_1 _18080_ (.A(_02234_),
    .B(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__nor2_1 _18081_ (.A(_01815_),
    .B(_01901_),
    .Y(_02237_));
 sky130_fd_sc_hd__xnor2_1 _18082_ (.A(_02236_),
    .B(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__and2_1 _18083_ (.A(_02233_),
    .B(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__or2_1 _18084_ (.A(_02233_),
    .B(_02238_),
    .X(_02240_));
 sky130_fd_sc_hd__and2b_1 _18085_ (.A_N(_02239_),
    .B(_02240_),
    .X(_02241_));
 sky130_fd_sc_hd__xnor2_1 _18086_ (.A(_02232_),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__a21oi_1 _18087_ (.A1(_02149_),
    .A2(_02231_),
    .B1(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__and3_1 _18088_ (.A(_02149_),
    .B(_02231_),
    .C(_02242_),
    .X(_02244_));
 sky130_fd_sc_hd__nor2_1 _18089_ (.A(_02243_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__xor2_1 _18090_ (.A(_02230_),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__xor2_1 _18091_ (.A(_02219_),
    .B(_02246_),
    .X(_02247_));
 sky130_fd_sc_hd__and2_1 _18092_ (.A(_02217_),
    .B(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__nor2_1 _18093_ (.A(_02217_),
    .B(_02247_),
    .Y(_02249_));
 sky130_fd_sc_hd__nor2_1 _18094_ (.A(_02248_),
    .B(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__xor2_1 _18095_ (.A(_02216_),
    .B(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__o21a_1 _18096_ (.A1(_02127_),
    .A2(_02128_),
    .B1(_02162_),
    .X(_02252_));
 sky130_fd_sc_hd__xnor2_1 _18097_ (.A(_02251_),
    .B(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__and2b_1 _18098_ (.A_N(_02160_),
    .B(_02130_),
    .X(_02254_));
 sky130_fd_sc_hd__o2bb2a_1 _18099_ (.A1_N(_02138_),
    .A2_N(_02139_),
    .B1(_02136_),
    .B2(_02137_),
    .X(_02255_));
 sky130_fd_sc_hd__o21ba_1 _18100_ (.A1(_02158_),
    .A2(_02254_),
    .B1_N(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__or3b_1 _18101_ (.A(_02158_),
    .B(_02254_),
    .C_N(_02255_),
    .X(_02257_));
 sky130_fd_sc_hd__and2b_1 _18102_ (.A_N(_02256_),
    .B(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__xor2_1 _18103_ (.A(_02253_),
    .B(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__o21a_1 _18104_ (.A1(_02164_),
    .A2(_02165_),
    .B1(_02167_),
    .X(_02260_));
 sky130_fd_sc_hd__xor2_1 _18105_ (.A(_02259_),
    .B(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__xnor2_1 _18106_ (.A(_02091_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__a21o_1 _18107_ (.A1(_02190_),
    .A2(_02191_),
    .B1(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__inv_2 _18108_ (.A(_02263_),
    .Y(_02264_));
 sky130_fd_sc_hd__and3_1 _18109_ (.A(_02190_),
    .B(_02191_),
    .C(_02262_),
    .X(_02265_));
 sky130_fd_sc_hd__nor2_1 _18110_ (.A(_02264_),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__inv_2 _18111_ (.A(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21oi_1 _18112_ (.A1(_02175_),
    .A2(_02179_),
    .B1(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__a31o_1 _18113_ (.A1(_02175_),
    .A2(_02179_),
    .A3(_02267_),
    .B1(_09937_),
    .X(_02269_));
 sky130_fd_sc_hd__or2_1 _18114_ (.A(_02268_),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__and2_1 _18115_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_02271_));
 sky130_fd_sc_hd__or2_1 _18116_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_02272_));
 sky130_fd_sc_hd__or2b_1 _18117_ (.A(_02271_),
    .B_N(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__nand2_1 _18118_ (.A(_02184_),
    .B(_02186_),
    .Y(_02274_));
 sky130_fd_sc_hd__and2_1 _18119_ (.A(_02183_),
    .B(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__xnor2_1 _18120_ (.A(_02273_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__a21oi_1 _18121_ (.A1(_09938_),
    .A2(_02276_),
    .B1(_09919_),
    .Y(_02277_));
 sky130_fd_sc_hd__o2bb2a_1 _18122_ (.A1_N(_02270_),
    .A2_N(_02277_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_09946_),
    .X(_00548_));
 sky130_fd_sc_hd__a21o_1 _18123_ (.A1(_02175_),
    .A2(_02263_),
    .B1(_02265_),
    .X(_02278_));
 sky130_fd_sc_hd__nor2_1 _18124_ (.A(_02259_),
    .B(_02260_),
    .Y(_02279_));
 sky130_fd_sc_hd__a21oi_1 _18125_ (.A1(_02091_),
    .A2(_02261_),
    .B1(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__o2bb2a_1 _18126_ (.A1_N(_02228_),
    .A2_N(_02229_),
    .B1(_02225_),
    .B2(_02227_),
    .X(_02281_));
 sky130_fd_sc_hd__xnor2_1 _18127_ (.A(_02280_),
    .B(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__or2b_1 _18128_ (.A(_02253_),
    .B_N(_02258_),
    .X(_02283_));
 sky130_fd_sc_hd__o21a_1 _18129_ (.A1(_02251_),
    .A2(_02252_),
    .B1(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__nor2_1 _18130_ (.A(_01710_),
    .B(_10473_),
    .Y(_02285_));
 sky130_fd_sc_hd__a21oi_1 _18131_ (.A1(_02200_),
    .A2(_02208_),
    .B1(_02206_),
    .Y(_02286_));
 sky130_fd_sc_hd__o22a_1 _18132_ (.A1(_01698_),
    .A2(_02196_),
    .B1(_10115_),
    .B2(_01700_),
    .X(_02287_));
 sky130_fd_sc_hd__or4_1 _18133_ (.A(_01700_),
    .B(_01698_),
    .C(_02196_),
    .D(_10115_),
    .X(_02288_));
 sky130_fd_sc_hd__and2b_1 _18134_ (.A_N(_02287_),
    .B(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__nor2_1 _18135_ (.A(_10445_),
    .B(_09703_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _18136_ (.A(_02105_),
    .B(_02197_),
    .Y(_02291_));
 sky130_fd_sc_hd__o31a_1 _18137_ (.A1(_10445_),
    .A2(_09565_),
    .A3(_02198_),
    .B1(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__o31a_1 _18138_ (.A1(_01815_),
    .A2(_01901_),
    .A3(_02236_),
    .B1(_02234_),
    .X(_02293_));
 sky130_fd_sc_hd__nor2_1 _18139_ (.A(_01816_),
    .B(_01901_),
    .Y(_02294_));
 sky130_fd_sc_hd__xor2_1 _18140_ (.A(_02293_),
    .B(_02294_),
    .X(_02295_));
 sky130_fd_sc_hd__nor2_1 _18141_ (.A(_01815_),
    .B(_02002_),
    .Y(_02296_));
 sky130_fd_sc_hd__xnor2_1 _18142_ (.A(_02221_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__or2_1 _18143_ (.A(_02223_),
    .B(_02224_),
    .X(_02298_));
 sky130_fd_sc_hd__o211a_1 _18144_ (.A1(_08360_),
    .A2(_09768_),
    .B1(_02222_),
    .C1(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__a211oi_1 _18145_ (.A1(_02222_),
    .A2(_02298_),
    .B1(_08360_),
    .C1(_09768_),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _18146_ (.A(_02299_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__xnor2_1 _18147_ (.A(_02297_),
    .B(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hd__xnor2_1 _18148_ (.A(_02295_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__xnor2_1 _18149_ (.A(_02292_),
    .B(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__xnor2_1 _18150_ (.A(_02290_),
    .B(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__xnor2_1 _18151_ (.A(_02289_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__xnor2_1 _18152_ (.A(_02286_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__xnor2_1 _18153_ (.A(_02285_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__a21o_1 _18154_ (.A1(_02230_),
    .A2(_02245_),
    .B1(_02243_),
    .X(_02309_));
 sky130_fd_sc_hd__or2_1 _18155_ (.A(_09446_),
    .B(_01790_),
    .X(_02310_));
 sky130_fd_sc_hd__a21oi_1 _18156_ (.A1(_02232_),
    .A2(_02241_),
    .B1(_02239_),
    .Y(_02311_));
 sky130_fd_sc_hd__xnor2_1 _18157_ (.A(_02310_),
    .B(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _18158_ (.A(_08303_),
    .B(_09755_),
    .Y(_02313_));
 sky130_fd_sc_hd__xnor2_1 _18159_ (.A(_02312_),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__xnor2_1 _18160_ (.A(_02309_),
    .B(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _18161_ (.A(_01676_),
    .B(_09565_),
    .Y(_02316_));
 sky130_fd_sc_hd__xnor2_1 _18162_ (.A(_02195_),
    .B(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__xnor2_1 _18163_ (.A(_02315_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__xnor2_1 _18164_ (.A(_02308_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__or2_1 _18165_ (.A(_01848_),
    .B(_02096_),
    .X(_02320_));
 sky130_fd_sc_hd__a32o_1 _18166_ (.A1(_10238_),
    .A2(_01730_),
    .A3(_02096_),
    .B1(_02320_),
    .B2(_02213_),
    .X(_02321_));
 sky130_fd_sc_hd__a21oi_1 _18167_ (.A1(_02193_),
    .A2(_02212_),
    .B1(_02210_),
    .Y(_02322_));
 sky130_fd_sc_hd__xnor2_1 _18168_ (.A(_02321_),
    .B(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__xnor2_1 _18169_ (.A(_02319_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__a21o_1 _18170_ (.A1(_02202_),
    .A2(_02204_),
    .B1(_02112_),
    .X(_02325_));
 sky130_fd_sc_hd__a21oi_1 _18171_ (.A1(_02219_),
    .A2(_02246_),
    .B1(_02248_),
    .Y(_02326_));
 sky130_fd_sc_hd__xnor2_1 _18172_ (.A(_02325_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__xnor2_1 _18173_ (.A(_02324_),
    .B(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__and2b_1 _18174_ (.A_N(_02216_),
    .B(_02250_),
    .X(_02329_));
 sky130_fd_sc_hd__a21o_1 _18175_ (.A1(_02192_),
    .A2(_02215_),
    .B1(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__xor2_1 _18176_ (.A(_02256_),
    .B(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__xnor2_1 _18177_ (.A(_02328_),
    .B(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__xnor2_1 _18178_ (.A(_02284_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__xnor2_1 _18179_ (.A(_02282_),
    .B(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__o211a_1 _18180_ (.A1(_02179_),
    .A2(_02267_),
    .B1(_02278_),
    .C1(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__a311o_1 _18181_ (.A1(_02175_),
    .A2(_02179_),
    .A3(_02263_),
    .B1(_02265_),
    .C1(_02334_),
    .X(_02336_));
 sky130_fd_sc_hd__or3b_1 _18182_ (.A(_09938_),
    .B(_02335_),
    .C_N(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__a21oi_1 _18183_ (.A1(_02272_),
    .A2(_02275_),
    .B1(_02271_),
    .Y(_02338_));
 sky130_fd_sc_hd__xor2_1 _18184_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .X(_02339_));
 sky130_fd_sc_hd__xnor2_1 _18185_ (.A(_02338_),
    .B(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__a21oi_1 _18186_ (.A1(_09938_),
    .A2(_02340_),
    .B1(_09919_),
    .Y(_02341_));
 sky130_fd_sc_hd__o2bb2a_1 _18187_ (.A1_N(_02337_),
    .A2_N(_02341_),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_09946_),
    .X(_00549_));
 sky130_fd_sc_hd__and2_1 _18188_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_02342_));
 sky130_fd_sc_hd__nor2_1 _18189_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_02343_));
 sky130_fd_sc_hd__o21a_1 _18190_ (.A1(_06094_),
    .A2(_09069_),
    .B1(_06284_),
    .X(_02344_));
 sky130_fd_sc_hd__buf_4 _18191_ (.A(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__buf_4 _18192_ (.A(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__o31a_1 _18193_ (.A1(_10509_),
    .A2(_02342_),
    .A3(_02343_),
    .B1(_02346_),
    .X(_02347_));
 sky130_fd_sc_hd__clkbuf_4 _18194_ (.A(_02345_),
    .X(_02348_));
 sky130_fd_sc_hd__o2bb2a_1 _18195_ (.A1_N(_02347_),
    .A2_N(_09940_),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .B2(_02348_),
    .X(_00550_));
 sky130_fd_sc_hd__or2_1 _18196_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_02349_));
 sky130_fd_sc_hd__nand2_1 _18197_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_02350_));
 sky130_fd_sc_hd__and4_1 _18198_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .C(_02349_),
    .D(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__a22oi_1 _18199_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(\rbzero.wall_tracer.stepDistY[-11] ),
    .B1(_02349_),
    .B2(_02350_),
    .Y(_02352_));
 sky130_fd_sc_hd__o31a_1 _18200_ (.A1(_10509_),
    .A2(_02351_),
    .A3(_02352_),
    .B1(_02346_),
    .X(_02353_));
 sky130_fd_sc_hd__o2bb2a_1 _18201_ (.A1_N(_02353_),
    .A2_N(_09948_),
    .B1(\rbzero.wall_tracer.trackDistY[-10] ),
    .B2(_02348_),
    .X(_00551_));
 sky130_fd_sc_hd__a21oi_1 _18202_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(\rbzero.wall_tracer.stepDistY[-10] ),
    .B1(_02351_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _18203_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_02355_));
 sky130_fd_sc_hd__and2_1 _18204_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_02356_));
 sky130_fd_sc_hd__nor3_1 _18205_ (.A(_02354_),
    .B(_02355_),
    .C(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__o21a_1 _18206_ (.A1(_02355_),
    .A2(_02356_),
    .B1(_02354_),
    .X(_02358_));
 sky130_fd_sc_hd__o31a_1 _18207_ (.A1(_10509_),
    .A2(_02357_),
    .A3(_02358_),
    .B1(_02346_),
    .X(_02359_));
 sky130_fd_sc_hd__o2bb2a_1 _18208_ (.A1_N(_02359_),
    .A2_N(_09960_),
    .B1(\rbzero.wall_tracer.trackDistY[-9] ),
    .B2(_02348_),
    .X(_00552_));
 sky130_fd_sc_hd__or2_1 _18209_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_02360_));
 sky130_fd_sc_hd__nand2_1 _18210_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .Y(_02361_));
 sky130_fd_sc_hd__o21bai_1 _18211_ (.A1(_02354_),
    .A2(_02355_),
    .B1_N(_02356_),
    .Y(_02362_));
 sky130_fd_sc_hd__and3_1 _18212_ (.A(_02360_),
    .B(_02361_),
    .C(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__a21oi_1 _18213_ (.A1(_02360_),
    .A2(_02361_),
    .B1(_02362_),
    .Y(_02364_));
 sky130_fd_sc_hd__o31a_1 _18214_ (.A1(_10509_),
    .A2(_02363_),
    .A3(_02364_),
    .B1(_02346_),
    .X(_02365_));
 sky130_fd_sc_hd__o2bb2a_1 _18215_ (.A1_N(_02365_),
    .A2_N(_09967_),
    .B1(\rbzero.wall_tracer.trackDistY[-8] ),
    .B2(_02348_),
    .X(_00553_));
 sky130_fd_sc_hd__nor2_1 _18216_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _18217_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02367_));
 sky130_fd_sc_hd__or2b_1 _18218_ (.A(_02366_),
    .B_N(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__a21boi_1 _18219_ (.A1(_02360_),
    .A2(_02362_),
    .B1_N(_02361_),
    .Y(_02369_));
 sky130_fd_sc_hd__nor2_1 _18220_ (.A(_02368_),
    .B(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__a21o_1 _18221_ (.A1(_02368_),
    .A2(_02369_),
    .B1(_09974_),
    .X(_02371_));
 sky130_fd_sc_hd__o21ai_1 _18222_ (.A1(_02370_),
    .A2(_02371_),
    .B1(_09976_),
    .Y(_02372_));
 sky130_fd_sc_hd__mux2_1 _18223_ (.A0(\rbzero.wall_tracer.trackDistY[-7] ),
    .A1(_02372_),
    .S(_02345_),
    .X(_02373_));
 sky130_fd_sc_hd__clkbuf_1 _18224_ (.A(_02373_),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _18225_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_02374_));
 sky130_fd_sc_hd__nand2_1 _18226_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .Y(_02375_));
 sky130_fd_sc_hd__o21ai_1 _18227_ (.A1(_02366_),
    .A2(_02369_),
    .B1(_02367_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21oi_1 _18228_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__a31o_1 _18229_ (.A1(_02374_),
    .A2(_02375_),
    .A3(_02376_),
    .B1(_06287_),
    .X(_02378_));
 sky130_fd_sc_hd__clkbuf_4 _18230_ (.A(_02344_),
    .X(_02379_));
 sky130_fd_sc_hd__o21a_1 _18231_ (.A1(_02377_),
    .A2(_02378_),
    .B1(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__o2bb2a_1 _18232_ (.A1_N(_02380_),
    .A2_N(_09985_),
    .B1(\rbzero.wall_tracer.trackDistY[-6] ),
    .B2(_02348_),
    .X(_00555_));
 sky130_fd_sc_hd__nor2_1 _18233_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02381_));
 sky130_fd_sc_hd__nand2_1 _18234_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02382_));
 sky130_fd_sc_hd__or2b_1 _18235_ (.A(_02381_),
    .B_N(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__a21boi_1 _18236_ (.A1(_02374_),
    .A2(_02376_),
    .B1_N(_02375_),
    .Y(_02384_));
 sky130_fd_sc_hd__nor2_1 _18237_ (.A(_02383_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__a21o_1 _18238_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_09974_),
    .X(_02386_));
 sky130_fd_sc_hd__o21ai_1 _18239_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_09993_),
    .Y(_02387_));
 sky130_fd_sc_hd__mux2_1 _18240_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(_02387_),
    .S(_02345_),
    .X(_02388_));
 sky130_fd_sc_hd__clkbuf_1 _18241_ (.A(_02388_),
    .X(_00556_));
 sky130_fd_sc_hd__or2_1 _18242_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(_02389_));
 sky130_fd_sc_hd__nand2_1 _18243_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02390_));
 sky130_fd_sc_hd__o21ai_1 _18244_ (.A1(_02381_),
    .A2(_02384_),
    .B1(_02382_),
    .Y(_02391_));
 sky130_fd_sc_hd__and3_1 _18245_ (.A(_02389_),
    .B(_02390_),
    .C(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__a21oi_1 _18246_ (.A1(_02389_),
    .A2(_02390_),
    .B1(_02391_),
    .Y(_02393_));
 sky130_fd_sc_hd__o31a_1 _18247_ (.A1(_10509_),
    .A2(_02392_),
    .A3(_02393_),
    .B1(_02346_),
    .X(_02394_));
 sky130_fd_sc_hd__o2bb2a_1 _18248_ (.A1_N(_02394_),
    .A2_N(_10001_),
    .B1(\rbzero.wall_tracer.trackDistY[-4] ),
    .B2(_02348_),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _18249_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02395_));
 sky130_fd_sc_hd__nand2_1 _18250_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02396_));
 sky130_fd_sc_hd__or2b_1 _18251_ (.A(_02395_),
    .B_N(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__a21boi_1 _18252_ (.A1(_02389_),
    .A2(_02391_),
    .B1_N(_02390_),
    .Y(_02398_));
 sky130_fd_sc_hd__xnor2_1 _18253_ (.A(_02397_),
    .B(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__o21a_1 _18254_ (.A1(_06288_),
    .A2(_02399_),
    .B1(_02379_),
    .X(_02400_));
 sky130_fd_sc_hd__o2bb2a_1 _18255_ (.A1_N(_02400_),
    .A2_N(_10010_),
    .B1(\rbzero.wall_tracer.trackDistY[-3] ),
    .B2(_02348_),
    .X(_00558_));
 sky130_fd_sc_hd__or2_1 _18256_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_02401_));
 sky130_fd_sc_hd__nand2_1 _18257_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02402_));
 sky130_fd_sc_hd__o21ai_1 _18258_ (.A1(_02395_),
    .A2(_02398_),
    .B1(_02396_),
    .Y(_02403_));
 sky130_fd_sc_hd__and3_1 _18259_ (.A(_02401_),
    .B(_02402_),
    .C(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__a21oi_1 _18260_ (.A1(_02401_),
    .A2(_02402_),
    .B1(_02403_),
    .Y(_02405_));
 sky130_fd_sc_hd__o31a_1 _18261_ (.A1(_10509_),
    .A2(_02404_),
    .A3(_02405_),
    .B1(_02346_),
    .X(_02406_));
 sky130_fd_sc_hd__o2bb2a_1 _18262_ (.A1_N(_02406_),
    .A2_N(_10018_),
    .B1(\rbzero.wall_tracer.trackDistY[-2] ),
    .B2(_02348_),
    .X(_00559_));
 sky130_fd_sc_hd__nor2_1 _18263_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_02407_));
 sky130_fd_sc_hd__and2_1 _18264_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .X(_02408_));
 sky130_fd_sc_hd__or2_1 _18265_ (.A(_02407_),
    .B(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__a21boi_1 _18266_ (.A1(_02401_),
    .A2(_02403_),
    .B1_N(_02402_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor2_1 _18267_ (.A(_02409_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__a21o_1 _18268_ (.A1(_02409_),
    .A2(_02410_),
    .B1(_09974_),
    .X(_02412_));
 sky130_fd_sc_hd__o21ai_1 _18269_ (.A1(_02411_),
    .A2(_02412_),
    .B1(_10026_),
    .Y(_02413_));
 sky130_fd_sc_hd__mux2_1 _18270_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(_02413_),
    .S(_02345_),
    .X(_02414_));
 sky130_fd_sc_hd__clkbuf_1 _18271_ (.A(_02414_),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _18272_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .X(_02415_));
 sky130_fd_sc_hd__nand2_1 _18273_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_02416_));
 sky130_fd_sc_hd__a211oi_1 _18274_ (.A1(_02415_),
    .A2(_02416_),
    .B1(_02408_),
    .C1(_02411_),
    .Y(_02417_));
 sky130_fd_sc_hd__o211a_1 _18275_ (.A1(_02408_),
    .A2(_02411_),
    .B1(_02415_),
    .C1(_02416_),
    .X(_02418_));
 sky130_fd_sc_hd__o31a_1 _18276_ (.A1(_10509_),
    .A2(_02417_),
    .A3(_02418_),
    .B1(_02346_),
    .X(_02419_));
 sky130_fd_sc_hd__o2bb2a_1 _18277_ (.A1_N(_02419_),
    .A2_N(_10153_),
    .B1(\rbzero.wall_tracer.trackDistY[0] ),
    .B2(_02348_),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_1 _18278_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_02420_));
 sky130_fd_sc_hd__or2_1 _18279_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_02421_));
 sky130_fd_sc_hd__a21o_1 _18280_ (.A1(\rbzero.wall_tracer.trackDistY[0] ),
    .A2(\rbzero.wall_tracer.stepDistY[0] ),
    .B1(_02418_),
    .X(_02422_));
 sky130_fd_sc_hd__and3_1 _18281_ (.A(_02420_),
    .B(_02421_),
    .C(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__a21o_1 _18282_ (.A1(_02420_),
    .A2(_02421_),
    .B1(_02422_),
    .X(_02424_));
 sky130_fd_sc_hd__or3b_1 _18283_ (.A(_09974_),
    .B(_02423_),
    .C_N(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__nand2_1 _18284_ (.A(_10269_),
    .B(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__mux2_1 _18285_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(_02426_),
    .S(_02345_),
    .X(_02427_));
 sky130_fd_sc_hd__clkbuf_1 _18286_ (.A(_02427_),
    .X(_00562_));
 sky130_fd_sc_hd__inv_2 _18287_ (.A(_02420_),
    .Y(_02428_));
 sky130_fd_sc_hd__nand2_1 _18288_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_02429_));
 sky130_fd_sc_hd__or2_1 _18289_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_02430_));
 sky130_fd_sc_hd__o211ai_2 _18290_ (.A1(_02428_),
    .A2(_02423_),
    .B1(_02429_),
    .C1(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__a211o_1 _18291_ (.A1(_02429_),
    .A2(_02430_),
    .B1(_02428_),
    .C1(_02423_),
    .X(_02432_));
 sky130_fd_sc_hd__nand2_1 _18292_ (.A(_02431_),
    .B(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__o21a_1 _18293_ (.A1(_06288_),
    .A2(_02433_),
    .B1(_02379_),
    .X(_02434_));
 sky130_fd_sc_hd__o2bb2a_1 _18294_ (.A1_N(_02434_),
    .A2_N(_10391_),
    .B1(\rbzero.wall_tracer.trackDistY[2] ),
    .B2(_02348_),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _18295_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_02435_));
 sky130_fd_sc_hd__nor2_1 _18296_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_02436_));
 sky130_fd_sc_hd__o211a_1 _18297_ (.A1(_02435_),
    .A2(_02436_),
    .B1(_02429_),
    .C1(_02431_),
    .X(_02437_));
 sky130_fd_sc_hd__a211oi_2 _18298_ (.A1(_02429_),
    .A2(_02431_),
    .B1(_02435_),
    .C1(_02436_),
    .Y(_02438_));
 sky130_fd_sc_hd__o31a_1 _18299_ (.A1(_09954_),
    .A2(_02437_),
    .A3(_02438_),
    .B1(_02346_),
    .X(_02439_));
 sky130_fd_sc_hd__o2bb2a_1 _18300_ (.A1_N(_02439_),
    .A2_N(_10508_),
    .B1(\rbzero.wall_tracer.trackDistY[3] ),
    .B2(_02379_),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _18301_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .Y(_02440_));
 sky130_fd_sc_hd__or2_1 _18302_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_02441_));
 sky130_fd_sc_hd__o211a_1 _18303_ (.A1(_02435_),
    .A2(_02438_),
    .B1(_02440_),
    .C1(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__a211oi_1 _18304_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02435_),
    .C1(_02438_),
    .Y(_02443_));
 sky130_fd_sc_hd__o31a_1 _18305_ (.A1(_09954_),
    .A2(_02442_),
    .A3(_02443_),
    .B1(_02345_),
    .X(_02444_));
 sky130_fd_sc_hd__o2bb2a_1 _18306_ (.A1_N(_02444_),
    .A2_N(_01759_),
    .B1(\rbzero.wall_tracer.trackDistY[4] ),
    .B2(_02379_),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _18307_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_02445_));
 sky130_fd_sc_hd__and2_1 _18308_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_02446_));
 sky130_fd_sc_hd__a21oi_1 _18309_ (.A1(\rbzero.wall_tracer.trackDistY[4] ),
    .A2(\rbzero.wall_tracer.stepDistY[4] ),
    .B1(_02442_),
    .Y(_02447_));
 sky130_fd_sc_hd__o21a_1 _18310_ (.A1(_02445_),
    .A2(_02446_),
    .B1(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__nor3_1 _18311_ (.A(_02445_),
    .B(_02446_),
    .C(_02447_),
    .Y(_02449_));
 sky130_fd_sc_hd__o31a_1 _18312_ (.A1(_09954_),
    .A2(_02448_),
    .A3(_02449_),
    .B1(_02345_),
    .X(_02450_));
 sky130_fd_sc_hd__o2bb2a_1 _18313_ (.A1_N(_02450_),
    .A2_N(_01876_),
    .B1(\rbzero.wall_tracer.trackDistY[5] ),
    .B2(_02379_),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_1 _18314_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02451_));
 sky130_fd_sc_hd__and2_1 _18315_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .X(_02452_));
 sky130_fd_sc_hd__o21ba_1 _18316_ (.A1(_02445_),
    .A2(_02447_),
    .B1_N(_02446_),
    .X(_02453_));
 sky130_fd_sc_hd__o21ai_1 _18317_ (.A1(_02451_),
    .A2(_02452_),
    .B1(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__o31a_1 _18318_ (.A1(_02451_),
    .A2(_02452_),
    .A3(_02453_),
    .B1(_06095_),
    .X(_02455_));
 sky130_fd_sc_hd__a21bo_1 _18319_ (.A1(_02454_),
    .A2(_02455_),
    .B1_N(_01986_),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _18320_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(_02456_),
    .S(_02345_),
    .X(_02457_));
 sky130_fd_sc_hd__clkbuf_1 _18321_ (.A(_02457_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _18322_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02458_));
 sky130_fd_sc_hd__nand2_1 _18323_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02459_));
 sky130_fd_sc_hd__or2b_1 _18324_ (.A(_02458_),
    .B_N(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__o21ba_1 _18325_ (.A1(_02451_),
    .A2(_02453_),
    .B1_N(_02452_),
    .X(_02461_));
 sky130_fd_sc_hd__nor2_1 _18326_ (.A(_02460_),
    .B(_02461_),
    .Y(_02462_));
 sky130_fd_sc_hd__a21o_1 _18327_ (.A1(_02460_),
    .A2(_02461_),
    .B1(_09974_),
    .X(_02463_));
 sky130_fd_sc_hd__o21ai_1 _18328_ (.A1(_02462_),
    .A2(_02463_),
    .B1(_02087_),
    .Y(_02464_));
 sky130_fd_sc_hd__mux2_1 _18329_ (.A0(\rbzero.wall_tracer.trackDistY[7] ),
    .A1(_02464_),
    .S(_02345_),
    .X(_02465_));
 sky130_fd_sc_hd__clkbuf_1 _18330_ (.A(_02465_),
    .X(_00568_));
 sky130_fd_sc_hd__or2_1 _18331_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .X(_02466_));
 sky130_fd_sc_hd__nand2_1 _18332_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_02467_));
 sky130_fd_sc_hd__nand2_1 _18333_ (.A(_02466_),
    .B(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__o21a_1 _18334_ (.A1(_02458_),
    .A2(_02461_),
    .B1(_02459_),
    .X(_02469_));
 sky130_fd_sc_hd__nor2_1 _18335_ (.A(_02468_),
    .B(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__a21o_1 _18336_ (.A1(_02468_),
    .A2(_02469_),
    .B1(_09915_),
    .X(_02471_));
 sky130_fd_sc_hd__o21a_1 _18337_ (.A1(_02470_),
    .A2(_02471_),
    .B1(_02379_),
    .X(_02472_));
 sky130_fd_sc_hd__o2bb2a_1 _18338_ (.A1_N(_02472_),
    .A2_N(_02182_),
    .B1(\rbzero.wall_tracer.trackDistY[8] ),
    .B2(_02379_),
    .X(_00569_));
 sky130_fd_sc_hd__and2_1 _18339_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_02473_));
 sky130_fd_sc_hd__nor2_1 _18340_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_02474_));
 sky130_fd_sc_hd__nor2_1 _18341_ (.A(_02473_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__nand2_1 _18342_ (.A(_02467_),
    .B(_02469_),
    .Y(_02476_));
 sky130_fd_sc_hd__and2_1 _18343_ (.A(_02466_),
    .B(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__xnor2_1 _18344_ (.A(_02475_),
    .B(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__o21a_1 _18345_ (.A1(_06288_),
    .A2(_02478_),
    .B1(_02346_),
    .X(_02479_));
 sky130_fd_sc_hd__o2bb2a_1 _18346_ (.A1_N(_02479_),
    .A2_N(_02270_),
    .B1(\rbzero.wall_tracer.trackDistY[9] ),
    .B2(_02379_),
    .X(_00570_));
 sky130_fd_sc_hd__a31o_1 _18347_ (.A1(_02466_),
    .A2(_02475_),
    .A3(_02476_),
    .B1(_02473_),
    .X(_02480_));
 sky130_fd_sc_hd__xor2_1 _18348_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .X(_02481_));
 sky130_fd_sc_hd__xnor2_1 _18349_ (.A(_02480_),
    .B(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__o21a_1 _18350_ (.A1(_06288_),
    .A2(_02482_),
    .B1(_02346_),
    .X(_02483_));
 sky130_fd_sc_hd__o2bb2a_1 _18351_ (.A1_N(_02483_),
    .A2_N(_02337_),
    .B1(\rbzero.wall_tracer.trackDistY[10] ),
    .B2(_02379_),
    .X(_00571_));
 sky130_fd_sc_hd__buf_4 _18352_ (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_4 _18353_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02485_));
 sky130_fd_sc_hd__inv_2 _18354_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .Y(_02486_));
 sky130_fd_sc_hd__clkbuf_4 _18355_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_02487_));
 sky130_fd_sc_hd__clkbuf_4 _18356_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .X(_02488_));
 sky130_fd_sc_hd__and3b_1 _18357_ (.A_N(_02487_),
    .B(_02488_),
    .C(\rbzero.spi_registers.spi_done ),
    .X(_02489_));
 sky130_fd_sc_hd__and4_1 _18358_ (.A(_02485_),
    .B(_02486_),
    .C(_04108_),
    .D(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_4 _18359_ (.A(_02490_),
    .X(_02491_));
 sky130_fd_sc_hd__buf_4 _18360_ (.A(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _18361_ (.A0(\rbzero.spi_registers.new_texadd3[0] ),
    .A1(_02484_),
    .S(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _18362_ (.A(_02493_),
    .X(_00572_));
 sky130_fd_sc_hd__clkbuf_4 _18363_ (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _18364_ (.A0(\rbzero.spi_registers.new_texadd3[1] ),
    .A1(_02494_),
    .S(_02492_),
    .X(_02495_));
 sky130_fd_sc_hd__clkbuf_1 _18365_ (.A(_02495_),
    .X(_00573_));
 sky130_fd_sc_hd__clkbuf_4 _18366_ (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _18367_ (.A0(\rbzero.spi_registers.new_texadd3[2] ),
    .A1(_02496_),
    .S(_02492_),
    .X(_02497_));
 sky130_fd_sc_hd__clkbuf_1 _18368_ (.A(_02497_),
    .X(_00574_));
 sky130_fd_sc_hd__buf_4 _18369_ (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _18370_ (.A0(\rbzero.spi_registers.new_texadd3[3] ),
    .A1(_02498_),
    .S(_02492_),
    .X(_02499_));
 sky130_fd_sc_hd__clkbuf_1 _18371_ (.A(_02499_),
    .X(_00575_));
 sky130_fd_sc_hd__buf_4 _18372_ (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _18373_ (.A0(\rbzero.spi_registers.new_texadd3[4] ),
    .A1(_02500_),
    .S(_02492_),
    .X(_02501_));
 sky130_fd_sc_hd__clkbuf_1 _18374_ (.A(_02501_),
    .X(_00576_));
 sky130_fd_sc_hd__clkbuf_4 _18375_ (.A(\rbzero.spi_registers.spi_buffer[5] ),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _18376_ (.A0(\rbzero.spi_registers.new_texadd3[5] ),
    .A1(_02502_),
    .S(_02492_),
    .X(_02503_));
 sky130_fd_sc_hd__clkbuf_1 _18377_ (.A(_02503_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _18378_ (.A0(\rbzero.spi_registers.new_texadd3[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02492_),
    .X(_02504_));
 sky130_fd_sc_hd__clkbuf_1 _18379_ (.A(_02504_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _18380_ (.A0(\rbzero.spi_registers.new_texadd3[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02492_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _18381_ (.A(_02505_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _18382_ (.A0(\rbzero.spi_registers.new_texadd3[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02492_),
    .X(_02506_));
 sky130_fd_sc_hd__clkbuf_1 _18383_ (.A(_02506_),
    .X(_00580_));
 sky130_fd_sc_hd__buf_4 _18384_ (.A(_02491_),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _18385_ (.A0(\rbzero.spi_registers.new_texadd3[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__clkbuf_1 _18386_ (.A(_02508_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _18387_ (.A0(\rbzero.spi_registers.new_texadd3[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02507_),
    .X(_02509_));
 sky130_fd_sc_hd__clkbuf_1 _18388_ (.A(_02509_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _18389_ (.A0(\rbzero.spi_registers.new_texadd3[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_02507_),
    .X(_02510_));
 sky130_fd_sc_hd__clkbuf_1 _18390_ (.A(_02510_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _18391_ (.A0(\rbzero.spi_registers.new_texadd3[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_02507_),
    .X(_02511_));
 sky130_fd_sc_hd__clkbuf_1 _18392_ (.A(_02511_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _18393_ (.A0(\rbzero.spi_registers.new_texadd3[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_02507_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _18394_ (.A(_02512_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _18395_ (.A0(\rbzero.spi_registers.new_texadd3[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_02507_),
    .X(_02513_));
 sky130_fd_sc_hd__clkbuf_1 _18396_ (.A(_02513_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _18397_ (.A0(\rbzero.spi_registers.new_texadd3[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_02507_),
    .X(_02514_));
 sky130_fd_sc_hd__clkbuf_1 _18398_ (.A(_02514_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _18399_ (.A0(\rbzero.spi_registers.new_texadd3[16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_02507_),
    .X(_02515_));
 sky130_fd_sc_hd__clkbuf_1 _18400_ (.A(_02515_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _18401_ (.A0(\rbzero.spi_registers.new_texadd3[17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_02507_),
    .X(_02516_));
 sky130_fd_sc_hd__clkbuf_1 _18402_ (.A(_02516_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _18403_ (.A0(\rbzero.spi_registers.new_texadd3[18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_02507_),
    .X(_02517_));
 sky130_fd_sc_hd__clkbuf_1 _18404_ (.A(_02517_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _18405_ (.A0(\rbzero.spi_registers.new_texadd3[19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_02491_),
    .X(_02518_));
 sky130_fd_sc_hd__clkbuf_1 _18406_ (.A(_02518_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _18407_ (.A0(\rbzero.spi_registers.new_texadd3[20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_02491_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_1 _18408_ (.A(_02519_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _18409_ (.A0(\rbzero.spi_registers.new_texadd3[21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_02491_),
    .X(_02520_));
 sky130_fd_sc_hd__clkbuf_1 _18410_ (.A(_02520_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _18411_ (.A0(\rbzero.spi_registers.new_texadd3[22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_02491_),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _18412_ (.A(_02521_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _18413_ (.A0(\rbzero.spi_registers.new_texadd3[23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_02491_),
    .X(_02522_));
 sky130_fd_sc_hd__clkbuf_1 _18414_ (.A(_02522_),
    .X(_00595_));
 sky130_fd_sc_hd__nor2_1 _18415_ (.A(_05249_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _18416_ (.A(_05249_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02524_));
 sky130_fd_sc_hd__and2b_1 _18417_ (.A_N(_02523_),
    .B(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__clkbuf_4 _18418_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_02526_));
 sky130_fd_sc_hd__nor2_1 _18419_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2_1 _18420_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .Y(_02528_));
 sky130_fd_sc_hd__nand2_1 _18421_ (.A(_05246_),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_02529_));
 sky130_fd_sc_hd__or2_1 _18422_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_02530_));
 sky130_fd_sc_hd__nand2_1 _18423_ (.A(_02529_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__o21a_1 _18424_ (.A1(_02528_),
    .A2(_02531_),
    .B1(_02529_),
    .X(_02532_));
 sky130_fd_sc_hd__nand2_1 _18425_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02533_));
 sky130_fd_sc_hd__o21ai_1 _18426_ (.A1(_02527_),
    .A2(_02532_),
    .B1(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__a21o_1 _18427_ (.A1(_02526_),
    .A2(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B1(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__o21ai_1 _18428_ (.A1(_02526_),
    .A2(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B1(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__xnor2_1 _18429_ (.A(_02525_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__buf_2 _18430_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_02538_));
 sky130_fd_sc_hd__clkbuf_4 _18431_ (.A(_08261_),
    .X(_02539_));
 sky130_fd_sc_hd__a22o_1 _18432_ (.A1(_02538_),
    .A2(_02539_),
    .B1(_09886_),
    .B2(\rbzero.wall_tracer.rayAddendX[-5] ),
    .X(_02540_));
 sky130_fd_sc_hd__a21o_1 _18433_ (.A1(_09885_),
    .A2(_02537_),
    .B1(_02540_),
    .X(_00596_));
 sky130_fd_sc_hd__xnor2_1 _18434_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .Y(_02541_));
 sky130_fd_sc_hd__o21ai_1 _18435_ (.A1(_02523_),
    .A2(_02536_),
    .B1(_02524_),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_1 _18436_ (.A(_02541_),
    .B(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__clkbuf_4 _18437_ (.A(_08261_),
    .X(_02544_));
 sky130_fd_sc_hd__a211o_1 _18438_ (.A1(_02541_),
    .A2(_02542_),
    .B1(_02543_),
    .C1(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__nand2_1 _18439_ (.A(_05246_),
    .B(_02538_),
    .Y(_02546_));
 sky130_fd_sc_hd__or2_1 _18440_ (.A(_05246_),
    .B(_02538_),
    .X(_02547_));
 sky130_fd_sc_hd__a31o_1 _18441_ (.A1(_02544_),
    .A2(_02546_),
    .A3(_02547_),
    .B1(_09884_),
    .X(_02548_));
 sky130_fd_sc_hd__a22o_1 _18442_ (.A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_09894_),
    .B1(_02545_),
    .B2(_02548_),
    .X(_00597_));
 sky130_fd_sc_hd__or2_1 _18443_ (.A(_04566_),
    .B(_09878_),
    .X(_02549_));
 sky130_fd_sc_hd__buf_4 _18444_ (.A(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__buf_4 _18445_ (.A(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__nor2_1 _18446_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02552_));
 sky130_fd_sc_hd__and2_1 _18447_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .X(_02553_));
 sky130_fd_sc_hd__a21o_1 _18448_ (.A1(\rbzero.debug_overlay.vplaneX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B1(_02542_),
    .X(_02554_));
 sky130_fd_sc_hd__o21ai_1 _18449_ (.A1(\rbzero.debug_overlay.vplaneX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B1(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__o21ai_1 _18450_ (.A1(_02552_),
    .A2(_02553_),
    .B1(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__o311a_1 _18451_ (.A1(_02552_),
    .A2(_02553_),
    .A3(_02555_),
    .B1(_02556_),
    .C1(_04576_),
    .X(_02557_));
 sky130_fd_sc_hd__or3_1 _18452_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_05246_),
    .C(_02538_),
    .X(_02558_));
 sky130_fd_sc_hd__o21ai_1 _18453_ (.A1(_05246_),
    .A2(_02538_),
    .B1(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_02559_));
 sky130_fd_sc_hd__a31o_1 _18454_ (.A1(_02539_),
    .A2(_02558_),
    .A3(_02559_),
    .B1(_09881_),
    .X(_02560_));
 sky130_fd_sc_hd__o22a_1 _18455_ (.A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A2(_02551_),
    .B1(_02557_),
    .B2(_02560_),
    .X(_00598_));
 sky130_fd_sc_hd__nor2_1 _18456_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_02561_));
 sky130_fd_sc_hd__and2_1 _18457_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02562_));
 sky130_fd_sc_hd__nand2_1 _18458_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02563_));
 sky130_fd_sc_hd__o21ai_1 _18459_ (.A1(_02552_),
    .A2(_02555_),
    .B1(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__or3_1 _18460_ (.A(_02561_),
    .B(_02562_),
    .C(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__o21ai_1 _18461_ (.A1(_02561_),
    .A2(_02562_),
    .B1(_02564_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21oi_1 _18462_ (.A1(_02565_),
    .A2(_02566_),
    .B1(_08262_),
    .Y(_02567_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(_02526_),
    .B(_02558_),
    .Y(_02568_));
 sky130_fd_sc_hd__or2_1 _18464_ (.A(_02526_),
    .B(_02558_),
    .X(_02569_));
 sky130_fd_sc_hd__a31o_1 _18465_ (.A1(_02539_),
    .A2(_02568_),
    .A3(_02569_),
    .B1(_09881_),
    .X(_02570_));
 sky130_fd_sc_hd__o22a_1 _18466_ (.A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A2(_02551_),
    .B1(_02567_),
    .B2(_02570_),
    .X(_00599_));
 sky130_fd_sc_hd__buf_6 _18467_ (.A(_09884_),
    .X(_02571_));
 sky130_fd_sc_hd__or2_1 _18468_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02572_));
 sky130_fd_sc_hd__nand2_1 _18469_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_02573_));
 sky130_fd_sc_hd__nor2_1 _18470_ (.A(_02562_),
    .B(_02564_),
    .Y(_02574_));
 sky130_fd_sc_hd__nor2_1 _18471_ (.A(_02561_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__nand3_1 _18472_ (.A(_02572_),
    .B(_02573_),
    .C(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__a21o_1 _18473_ (.A1(_02572_),
    .A2(_02573_),
    .B1(_02575_),
    .X(_02577_));
 sky130_fd_sc_hd__inv_2 _18474_ (.A(_02538_),
    .Y(_02578_));
 sky130_fd_sc_hd__o31a_1 _18475_ (.A1(_02526_),
    .A2(\rbzero.debug_overlay.vplaneX[-7] ),
    .A3(_05246_),
    .B1(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__xor2_1 _18476_ (.A(_05249_),
    .B(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__a22o_1 _18477_ (.A1(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A2(_09880_),
    .B1(_02580_),
    .B2(_02539_),
    .X(_02581_));
 sky130_fd_sc_hd__a31o_1 _18478_ (.A1(_02571_),
    .A2(_02576_),
    .A3(_02577_),
    .B1(_02581_),
    .X(_00600_));
 sky130_fd_sc_hd__a21bo_1 _18479_ (.A1(_02572_),
    .A2(_02575_),
    .B1_N(_02573_),
    .X(_02582_));
 sky130_fd_sc_hd__buf_2 _18480_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_02583_));
 sky130_fd_sc_hd__nor2_1 _18481_ (.A(_02583_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_02584_));
 sky130_fd_sc_hd__and2_1 _18482_ (.A(_02583_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_02585_));
 sky130_fd_sc_hd__or2_1 _18483_ (.A(_02584_),
    .B(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__xnor2_1 _18484_ (.A(_02582_),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__or2_1 _18485_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(_05246_),
    .X(_02588_));
 sky130_fd_sc_hd__nand2_1 _18486_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(_05246_),
    .Y(_02589_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_02588_),
    .B(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__nor2_1 _18488_ (.A(_05249_),
    .B(_02569_),
    .Y(_02591_));
 sky130_fd_sc_hd__a21oi_1 _18489_ (.A1(_05249_),
    .A2(_02538_),
    .B1(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__xnor2_1 _18490_ (.A(_02590_),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__mux2_1 _18491_ (.A0(_02587_),
    .A1(_02593_),
    .S(_04566_),
    .X(_02594_));
 sky130_fd_sc_hd__mux2_1 _18492_ (.A0(\rbzero.wall_tracer.rayAddendX[0] ),
    .A1(_02594_),
    .S(_02550_),
    .X(_02595_));
 sky130_fd_sc_hd__clkbuf_1 _18493_ (.A(_02595_),
    .X(_00601_));
 sky130_fd_sc_hd__nand2_1 _18494_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_02596_));
 sky130_fd_sc_hd__or2_1 _18495_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02597_));
 sky130_fd_sc_hd__o21a_1 _18496_ (.A1(_02583_),
    .A2(\rbzero.wall_tracer.rayAddendX[0] ),
    .B1(_02582_),
    .X(_02598_));
 sky130_fd_sc_hd__a211o_1 _18497_ (.A1(_02596_),
    .A2(_02597_),
    .B1(_02598_),
    .C1(_02585_),
    .X(_02599_));
 sky130_fd_sc_hd__o211ai_2 _18498_ (.A1(_02585_),
    .A2(_02598_),
    .B1(_02597_),
    .C1(_02596_),
    .Y(_02600_));
 sky130_fd_sc_hd__a21oi_1 _18499_ (.A1(_05249_),
    .A2(_02538_),
    .B1(_02590_),
    .Y(_02601_));
 sky130_fd_sc_hd__nor2_1 _18500_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_02602_));
 sky130_fd_sc_hd__and2_1 _18501_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_02603_));
 sky130_fd_sc_hd__nor2_1 _18502_ (.A(_02602_),
    .B(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__xnor2_1 _18503_ (.A(_02588_),
    .B(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__o21a_1 _18504_ (.A1(_02591_),
    .A2(_02601_),
    .B1(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__inv_2 _18505_ (.A(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__or3_1 _18506_ (.A(_02591_),
    .B(_02605_),
    .C(_02601_),
    .X(_02608_));
 sky130_fd_sc_hd__a32o_1 _18507_ (.A1(_02544_),
    .A2(_02607_),
    .A3(_02608_),
    .B1(_09886_),
    .B2(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02609_));
 sky130_fd_sc_hd__a31o_1 _18508_ (.A1(_02571_),
    .A2(_02599_),
    .A3(_02600_),
    .B1(_02609_),
    .X(_00602_));
 sky130_fd_sc_hd__buf_2 _18509_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_02610_));
 sky130_fd_sc_hd__buf_2 _18510_ (.A(_02610_),
    .X(_02611_));
 sky130_fd_sc_hd__clkbuf_4 _18511_ (.A(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__xnor2_1 _18512_ (.A(_02612_),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_02613_));
 sky130_fd_sc_hd__a21oi_1 _18513_ (.A1(_02596_),
    .A2(_02600_),
    .B1(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__a311oi_1 _18514_ (.A1(_02596_),
    .A2(_02600_),
    .A3(_02613_),
    .B1(_02614_),
    .C1(_08262_),
    .Y(_02615_));
 sky130_fd_sc_hd__xor2_1 _18515_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(_02526_),
    .X(_02616_));
 sky130_fd_sc_hd__o31ai_1 _18516_ (.A1(_02588_),
    .A2(_02602_),
    .A3(_02603_),
    .B1(_02607_),
    .Y(_02617_));
 sky130_fd_sc_hd__xnor2_1 _18517_ (.A(_02616_),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__xnor2_1 _18518_ (.A(_02602_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__a21o_1 _18519_ (.A1(_08262_),
    .A2(_02619_),
    .B1(_09886_),
    .X(_02620_));
 sky130_fd_sc_hd__o22a_1 _18520_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(_02551_),
    .B1(_02615_),
    .B2(_02620_),
    .X(_00603_));
 sky130_fd_sc_hd__nand2_1 _18521_ (.A(_02616_),
    .B(_02617_),
    .Y(_02621_));
 sky130_fd_sc_hd__or2_1 _18522_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05249_),
    .X(_02622_));
 sky130_fd_sc_hd__nand2_1 _18523_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05249_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_1 _18524_ (.A(_02622_),
    .B(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__or3_1 _18525_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(_02526_),
    .C(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__o21ai_1 _18526_ (.A1(\rbzero.debug_overlay.vplaneX[-2] ),
    .A2(_02526_),
    .B1(_02624_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand2_1 _18527_ (.A(_02625_),
    .B(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__o21ai_1 _18528_ (.A1(_02606_),
    .A2(_02616_),
    .B1(_02602_),
    .Y(_02628_));
 sky130_fd_sc_hd__a31o_1 _18529_ (.A1(_02621_),
    .A2(_02627_),
    .A3(_02628_),
    .B1(_04568_),
    .X(_02629_));
 sky130_fd_sc_hd__a21o_1 _18530_ (.A1(_02621_),
    .A2(_02628_),
    .B1(_02627_),
    .X(_02630_));
 sky130_fd_sc_hd__and2b_1 _18531_ (.A_N(_02629_),
    .B(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__and4_1 _18532_ (.A(_04186_),
    .B(_04770_),
    .C(_05200_),
    .D(_09865_),
    .X(_02632_));
 sky130_fd_sc_hd__and4_2 _18533_ (.A(_04571_),
    .B(_04568_),
    .C(_05173_),
    .D(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__o21ai_1 _18534_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[1] ),
    .B1(_02610_),
    .Y(_02634_));
 sky130_fd_sc_hd__o21bai_1 _18535_ (.A1(_02610_),
    .A2(\rbzero.wall_tracer.rayAddendX[2] ),
    .B1_N(_02600_),
    .Y(_02635_));
 sky130_fd_sc_hd__and2_1 _18536_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02636_));
 sky130_fd_sc_hd__nor2_1 _18537_ (.A(_02610_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02637_));
 sky130_fd_sc_hd__a211o_1 _18538_ (.A1(_02634_),
    .A2(_02635_),
    .B1(_02636_),
    .C1(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__o211ai_1 _18539_ (.A1(_02636_),
    .A2(_02637_),
    .B1(_02634_),
    .C1(_02635_),
    .Y(_02639_));
 sky130_fd_sc_hd__a32o_1 _18540_ (.A1(_02633_),
    .A2(_02638_),
    .A3(_02639_),
    .B1(_09880_),
    .B2(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02640_));
 sky130_fd_sc_hd__or2_1 _18541_ (.A(_02631_),
    .B(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__clkbuf_1 _18542_ (.A(_02641_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _18543_ (.A(_02612_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02642_));
 sky130_fd_sc_hd__xor2_1 _18544_ (.A(_02610_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_02643_));
 sky130_fd_sc_hd__a21oi_1 _18545_ (.A1(_02642_),
    .A2(_02638_),
    .B1(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__a31o_1 _18546_ (.A1(_02642_),
    .A2(_02638_),
    .A3(_02643_),
    .B1(_04566_),
    .X(_02645_));
 sky130_fd_sc_hd__or2_1 _18547_ (.A(_02583_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_02646_));
 sky130_fd_sc_hd__nand2_1 _18548_ (.A(_02583_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .Y(_02647_));
 sky130_fd_sc_hd__nand2_1 _18549_ (.A(_02646_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__a21o_1 _18550_ (.A1(_02625_),
    .A2(_02630_),
    .B1(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__nand3_1 _18551_ (.A(_02625_),
    .B(_02630_),
    .C(_02648_),
    .Y(_02650_));
 sky130_fd_sc_hd__and2_1 _18552_ (.A(_02649_),
    .B(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__xnor2_1 _18553_ (.A(_02622_),
    .B(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hd__o22a_1 _18554_ (.A1(_02644_),
    .A2(_02645_),
    .B1(_02652_),
    .B2(_04568_),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _18555_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02653_),
    .S(_02550_),
    .X(_02654_));
 sky130_fd_sc_hd__clkbuf_1 _18556_ (.A(_02654_),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _18557_ (.A(_02610_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02655_));
 sky130_fd_sc_hd__or2_1 _18558_ (.A(_02610_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_02656_));
 sky130_fd_sc_hd__and2_1 _18559_ (.A(_02655_),
    .B(_02656_),
    .X(_02657_));
 sky130_fd_sc_hd__and2b_1 _18560_ (.A_N(_02638_),
    .B(_02643_),
    .X(_02658_));
 sky130_fd_sc_hd__o21ai_1 _18561_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02611_),
    .Y(_02659_));
 sky130_fd_sc_hd__inv_2 _18562_ (.A(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__or3_1 _18563_ (.A(_02657_),
    .B(_02658_),
    .C(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__o21ai_1 _18564_ (.A1(_02658_),
    .A2(_02660_),
    .B1(_02657_),
    .Y(_02662_));
 sky130_fd_sc_hd__nor2_1 _18565_ (.A(_02610_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .Y(_02663_));
 sky130_fd_sc_hd__and2_1 _18566_ (.A(_02610_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_02664_));
 sky130_fd_sc_hd__o21a_1 _18567_ (.A1(_02663_),
    .A2(_02664_),
    .B1(_02646_),
    .X(_02665_));
 sky130_fd_sc_hd__nor3_1 _18568_ (.A(_02646_),
    .B(_02663_),
    .C(_02664_),
    .Y(_02666_));
 sky130_fd_sc_hd__nor2_1 _18569_ (.A(_02665_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__a22o_1 _18570_ (.A1(_02630_),
    .A2(_02648_),
    .B1(_02649_),
    .B2(_02622_),
    .X(_02668_));
 sky130_fd_sc_hd__xnor2_1 _18571_ (.A(_02667_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a22o_1 _18572_ (.A1(\rbzero.wall_tracer.rayAddendX[5] ),
    .A2(_09880_),
    .B1(_02669_),
    .B2(_02539_),
    .X(_02670_));
 sky130_fd_sc_hd__a31o_1 _18573_ (.A1(_09888_),
    .A2(_02661_),
    .A3(_02662_),
    .B1(_02670_),
    .X(_00606_));
 sky130_fd_sc_hd__xnor2_1 _18574_ (.A(_02610_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_02671_));
 sky130_fd_sc_hd__nand3_1 _18575_ (.A(_02655_),
    .B(_02662_),
    .C(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__a21o_1 _18576_ (.A1(_02655_),
    .A2(_02662_),
    .B1(_02671_),
    .X(_02673_));
 sky130_fd_sc_hd__or2_1 _18577_ (.A(_02611_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_02674_));
 sky130_fd_sc_hd__nand2_1 _18578_ (.A(_02611_),
    .B(\rbzero.debug_overlay.vplaneX[-2] ),
    .Y(_02675_));
 sky130_fd_sc_hd__a21o_1 _18579_ (.A1(_02674_),
    .A2(_02675_),
    .B1(_02663_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_1 _18580_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(_02663_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_1 _18581_ (.A(_02676_),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__o21bai_1 _18582_ (.A1(_02665_),
    .A2(_02668_),
    .B1_N(_02666_),
    .Y(_02679_));
 sky130_fd_sc_hd__xnor2_1 _18583_ (.A(_02678_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__a22o_1 _18584_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(_09880_),
    .B1(_02680_),
    .B2(_02539_),
    .X(_02681_));
 sky130_fd_sc_hd__a31o_1 _18585_ (.A1(_09888_),
    .A2(_02672_),
    .A3(_02673_),
    .B1(_02681_),
    .X(_00607_));
 sky130_fd_sc_hd__nand2_1 _18586_ (.A(_02611_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_02682_));
 sky130_fd_sc_hd__or2_1 _18587_ (.A(_02611_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02683_));
 sky130_fd_sc_hd__inv_2 _18588_ (.A(_02671_),
    .Y(_02684_));
 sky130_fd_sc_hd__o21a_1 _18589_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .B1(_02611_),
    .X(_02685_));
 sky130_fd_sc_hd__a311o_1 _18590_ (.A1(_02657_),
    .A2(_02658_),
    .A3(_02684_),
    .B1(_02685_),
    .C1(_02660_),
    .X(_02686_));
 sky130_fd_sc_hd__a21o_1 _18591_ (.A1(_02682_),
    .A2(_02683_),
    .B1(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__nand3_1 _18592_ (.A(_02682_),
    .B(_02683_),
    .C(_02686_),
    .Y(_02688_));
 sky130_fd_sc_hd__inv_2 _18593_ (.A(_02677_),
    .Y(_02689_));
 sky130_fd_sc_hd__and3_1 _18594_ (.A(_02676_),
    .B(_02677_),
    .C(_02679_),
    .X(_02690_));
 sky130_fd_sc_hd__nor2_1 _18595_ (.A(_02611_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .Y(_02691_));
 sky130_fd_sc_hd__and2_1 _18596_ (.A(_02611_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_02692_));
 sky130_fd_sc_hd__o21ai_1 _18597_ (.A1(_02691_),
    .A2(_02692_),
    .B1(_02674_),
    .Y(_02693_));
 sky130_fd_sc_hd__or3_1 _18598_ (.A(_02674_),
    .B(_02691_),
    .C(_02692_),
    .X(_02694_));
 sky130_fd_sc_hd__o211ai_2 _18599_ (.A1(_02689_),
    .A2(_02690_),
    .B1(_02693_),
    .C1(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__a211o_1 _18600_ (.A1(_02693_),
    .A2(_02694_),
    .B1(_02689_),
    .C1(_02690_),
    .X(_02696_));
 sky130_fd_sc_hd__a32o_1 _18601_ (.A1(_02544_),
    .A2(_02695_),
    .A3(_02696_),
    .B1(_09886_),
    .B2(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02697_));
 sky130_fd_sc_hd__a31o_1 _18602_ (.A1(_09888_),
    .A2(_02687_),
    .A3(_02688_),
    .B1(_02697_),
    .X(_00608_));
 sky130_fd_sc_hd__nand2_1 _18603_ (.A(_02612_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_02698_));
 sky130_fd_sc_hd__or2_1 _18604_ (.A(_02611_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_02699_));
 sky130_fd_sc_hd__nand2_1 _18605_ (.A(_02698_),
    .B(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hd__a21oi_1 _18606_ (.A1(_02682_),
    .A2(_02688_),
    .B1(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__a31o_1 _18607_ (.A1(_02682_),
    .A2(_02688_),
    .A3(_02700_),
    .B1(_08261_),
    .X(_02702_));
 sky130_fd_sc_hd__nor2_1 _18608_ (.A(_02701_),
    .B(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__inv_2 _18609_ (.A(_02583_),
    .Y(_02704_));
 sky130_fd_sc_hd__a21oi_1 _18610_ (.A1(_02583_),
    .A2(\rbzero.debug_overlay.vplaneX[-1] ),
    .B1(_02612_),
    .Y(_02705_));
 sky130_fd_sc_hd__a21oi_1 _18611_ (.A1(_02612_),
    .A2(_02583_),
    .B1(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__a21oi_1 _18612_ (.A1(_02704_),
    .A2(_02691_),
    .B1(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__a21o_1 _18613_ (.A1(_02694_),
    .A2(_02695_),
    .B1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__nand3_1 _18614_ (.A(_02694_),
    .B(_02695_),
    .C(_02707_),
    .Y(_02709_));
 sky130_fd_sc_hd__a31o_1 _18615_ (.A1(_02539_),
    .A2(_02708_),
    .A3(_02709_),
    .B1(_09881_),
    .X(_02710_));
 sky130_fd_sc_hd__o22a_1 _18616_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(_02551_),
    .B1(_02703_),
    .B2(_02710_),
    .X(_00609_));
 sky130_fd_sc_hd__or2_1 _18617_ (.A(_02612_),
    .B(_02583_),
    .X(_02711_));
 sky130_fd_sc_hd__mux2_1 _18618_ (.A0(_02711_),
    .A1(_02705_),
    .S(_02708_),
    .X(_02712_));
 sky130_fd_sc_hd__or2_1 _18619_ (.A(_02612_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_02713_));
 sky130_fd_sc_hd__nand2_1 _18620_ (.A(_02612_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_02714_));
 sky130_fd_sc_hd__nand2_1 _18621_ (.A(_02713_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__o211a_1 _18622_ (.A1(_02688_),
    .A2(_02700_),
    .B1(_02698_),
    .C1(_02682_),
    .X(_02716_));
 sky130_fd_sc_hd__xnor2_1 _18623_ (.A(_02715_),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__o2bb2a_1 _18624_ (.A1_N(_02633_),
    .A2_N(_02717_),
    .B1(\rbzero.wall_tracer.rayAddendX[9] ),
    .B2(_02550_),
    .X(_02718_));
 sky130_fd_sc_hd__o21a_1 _18625_ (.A1(_04576_),
    .A2(_02712_),
    .B1(_02718_),
    .X(_00610_));
 sky130_fd_sc_hd__or2_1 _18626_ (.A(_02715_),
    .B(_02716_),
    .X(_02719_));
 sky130_fd_sc_hd__xnor2_1 _18627_ (.A(_02612_),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_02720_));
 sky130_fd_sc_hd__a21oi_1 _18628_ (.A1(_02714_),
    .A2(_02719_),
    .B1(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__a311oi_1 _18629_ (.A1(_02714_),
    .A2(_02719_),
    .A3(_02720_),
    .B1(_02721_),
    .C1(_08262_),
    .Y(_02722_));
 sky130_fd_sc_hd__inv_2 _18630_ (.A(_02612_),
    .Y(_02723_));
 sky130_fd_sc_hd__or2_1 _18631_ (.A(_02583_),
    .B(_02708_),
    .X(_02724_));
 sky130_fd_sc_hd__a31o_1 _18632_ (.A1(_02723_),
    .A2(_08261_),
    .A3(_02724_),
    .B1(_09881_),
    .X(_02725_));
 sky130_fd_sc_hd__o22a_1 _18633_ (.A1(\rbzero.wall_tracer.rayAddendX[10] ),
    .A2(_02551_),
    .B1(_02722_),
    .B2(_02725_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _18634_ (.A0(\rbzero.debug_overlay.playerY[0] ),
    .A1(_06187_),
    .S(_06095_),
    .X(_02726_));
 sky130_fd_sc_hd__mux2_1 _18635_ (.A0(_02726_),
    .A1(_06229_),
    .S(_06286_),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_1 _18636_ (.A(_02727_),
    .X(_00612_));
 sky130_fd_sc_hd__or2_1 _18637_ (.A(_06229_),
    .B(_06378_),
    .X(_02728_));
 sky130_fd_sc_hd__inv_2 _18638_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .Y(_02729_));
 sky130_fd_sc_hd__nor2_1 _18639_ (.A(_02729_),
    .B(_09937_),
    .Y(_02730_));
 sky130_fd_sc_hd__a31o_1 _18640_ (.A1(_09937_),
    .A2(_06379_),
    .A3(_02728_),
    .B1(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__mux2_1 _18641_ (.A0(_02731_),
    .A1(\rbzero.map_rom.c6 ),
    .S(_06286_),
    .X(_02732_));
 sky130_fd_sc_hd__clkbuf_1 _18642_ (.A(_02732_),
    .X(_00613_));
 sky130_fd_sc_hd__or2_1 _18643_ (.A(_06380_),
    .B(_06381_),
    .X(_02733_));
 sky130_fd_sc_hd__and3_1 _18644_ (.A(_09938_),
    .B(_06382_),
    .C(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__a21o_1 _18645_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_06288_),
    .B1(_06286_),
    .X(_02735_));
 sky130_fd_sc_hd__o2bb2a_1 _18646_ (.A1_N(_06193_),
    .A2_N(_06286_),
    .B1(_02734_),
    .B2(_02735_),
    .X(_00614_));
 sky130_fd_sc_hd__nand2_1 _18647_ (.A(_06376_),
    .B(_06384_),
    .Y(_02736_));
 sky130_fd_sc_hd__xnor2_1 _18648_ (.A(_06383_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__mux2_1 _18649_ (.A0(\rbzero.debug_overlay.playerY[3] ),
    .A1(_02737_),
    .S(_06095_),
    .X(_02738_));
 sky130_fd_sc_hd__mux2_1 _18650_ (.A0(_02738_),
    .A1(\rbzero.map_rom.a6 ),
    .S(_06285_),
    .X(_02739_));
 sky130_fd_sc_hd__clkbuf_1 _18651_ (.A(_02739_),
    .X(_00615_));
 sky130_fd_sc_hd__a21oi_1 _18652_ (.A1(_06376_),
    .A2(_06385_),
    .B1(_06375_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand2_1 _18653_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .B(_06287_),
    .Y(_02741_));
 sky130_fd_sc_hd__o31ai_1 _18654_ (.A1(_09915_),
    .A2(_06386_),
    .A3(_02740_),
    .B1(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__mux2_1 _18655_ (.A0(_02742_),
    .A1(\rbzero.map_rom.i_row[4] ),
    .S(_06285_),
    .X(_02743_));
 sky130_fd_sc_hd__clkbuf_1 _18656_ (.A(_02743_),
    .X(_00616_));
 sky130_fd_sc_hd__a21oi_1 _18657_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(_06372_),
    .B1(_06386_),
    .Y(_02744_));
 sky130_fd_sc_hd__xnor2_1 _18658_ (.A(_06374_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__mux2_1 _18659_ (.A0(\rbzero.debug_overlay.playerY[5] ),
    .A1(_02745_),
    .S(_06095_),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _18660_ (.A0(_02746_),
    .A1(\rbzero.wall_tracer.mapY[5] ),
    .S(_06285_),
    .X(_02747_));
 sky130_fd_sc_hd__clkbuf_1 _18661_ (.A(_02747_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _18662_ (.A0(\rbzero.debug_overlay.playerX[0] ),
    .A1(_06204_),
    .S(_06095_),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _18663_ (.A0(_02748_),
    .A1(_06220_),
    .S(_09919_),
    .X(_02749_));
 sky130_fd_sc_hd__clkbuf_1 _18664_ (.A(_02749_),
    .X(_00618_));
 sky130_fd_sc_hd__nor2_1 _18665_ (.A(_06220_),
    .B(_09904_),
    .Y(_02750_));
 sky130_fd_sc_hd__or2_1 _18666_ (.A(_09905_),
    .B(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__nor2_1 _18667_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_09937_),
    .Y(_02752_));
 sky130_fd_sc_hd__a211o_1 _18668_ (.A1(_09938_),
    .A2(_02751_),
    .B1(_02752_),
    .C1(_09919_),
    .X(_02753_));
 sky130_fd_sc_hd__o21ai_1 _18669_ (.A1(_06183_),
    .A2(_09946_),
    .B1(_02753_),
    .Y(_00619_));
 sky130_fd_sc_hd__or3_1 _18670_ (.A(_09902_),
    .B(_09905_),
    .C(_09906_),
    .X(_02754_));
 sky130_fd_sc_hd__nor2_1 _18671_ (.A(_04804_),
    .B(_09937_),
    .Y(_02755_));
 sky130_fd_sc_hd__a31o_1 _18672_ (.A1(_09937_),
    .A2(_09907_),
    .A3(_02754_),
    .B1(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__mux2_1 _18673_ (.A0(_02756_),
    .A1(_06184_),
    .S(_09916_),
    .X(_02757_));
 sky130_fd_sc_hd__clkbuf_1 _18674_ (.A(_02757_),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _18675_ (.A(_09901_),
    .B(_09909_),
    .Y(_02758_));
 sky130_fd_sc_hd__xnor2_1 _18676_ (.A(_09908_),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__mux2_1 _18677_ (.A0(\rbzero.debug_overlay.playerX[3] ),
    .A1(_02759_),
    .S(_06095_),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _18678_ (.A0(_06223_),
    .A1(_02760_),
    .S(_09978_),
    .X(_02761_));
 sky130_fd_sc_hd__clkbuf_1 _18679_ (.A(_02761_),
    .X(_00621_));
 sky130_fd_sc_hd__a21oi_1 _18680_ (.A1(_09901_),
    .A2(_09910_),
    .B1(_09900_),
    .Y(_02762_));
 sky130_fd_sc_hd__nand2_1 _18681_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_06287_),
    .Y(_02763_));
 sky130_fd_sc_hd__o31ai_1 _18682_ (.A1(_09915_),
    .A2(_09911_),
    .A3(_02762_),
    .B1(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__mux2_1 _18683_ (.A0(\rbzero.map_rom.i_col[4] ),
    .A1(_02764_),
    .S(_09978_),
    .X(_02765_));
 sky130_fd_sc_hd__clkbuf_1 _18684_ (.A(_02765_),
    .X(_00622_));
 sky130_fd_sc_hd__a21oi_1 _18685_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(_09266_),
    .B1(_09911_),
    .Y(_02766_));
 sky130_fd_sc_hd__xnor2_1 _18686_ (.A(_09899_),
    .B(_02766_),
    .Y(_02767_));
 sky130_fd_sc_hd__mux2_1 _18687_ (.A0(\rbzero.debug_overlay.playerX[5] ),
    .A1(_02767_),
    .S(_06095_),
    .X(_02768_));
 sky130_fd_sc_hd__mux2_1 _18688_ (.A0(\rbzero.wall_tracer.mapX[5] ),
    .A1(_02768_),
    .S(_09944_),
    .X(_02769_));
 sky130_fd_sc_hd__clkbuf_1 _18689_ (.A(_02769_),
    .X(_00623_));
 sky130_fd_sc_hd__inv_2 _18690_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .Y(_02770_));
 sky130_fd_sc_hd__nor2b_2 _18691_ (.A(\rbzero.spi_registers.sclk_buffer[2] ),
    .B_N(\rbzero.spi_registers.sclk_buffer[1] ),
    .Y(_02771_));
 sky130_fd_sc_hd__inv_2 _18692_ (.A(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__nor2b_2 _18693_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B_N(\rbzero.spi_registers.spi_cmd[2] ),
    .Y(_02773_));
 sky130_fd_sc_hd__or2_1 _18694_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02774_));
 sky130_fd_sc_hd__a21oi_2 _18695_ (.A1(_02487_),
    .A2(_02774_),
    .B1(_02488_),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2_2 _18696_ (.A(_02485_),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .Y(_02776_));
 sky130_fd_sc_hd__and3b_1 _18697_ (.A_N(\rbzero.spi_registers.spi_cmd[2] ),
    .B(\rbzero.spi_registers.spi_cmd[3] ),
    .C(_02776_),
    .X(_02777_));
 sky130_fd_sc_hd__a311oi_4 _18698_ (.A1(_02485_),
    .A2(\rbzero.spi_registers.spi_cmd[0] ),
    .A3(_02773_),
    .B1(_02775_),
    .C1(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand3_2 _18699_ (.A(_02485_),
    .B(_02486_),
    .C(_02773_),
    .Y(_02779_));
 sky130_fd_sc_hd__nand2_1 _18700_ (.A(_02779_),
    .B(_02778_),
    .Y(_02780_));
 sky130_fd_sc_hd__o211a_1 _18701_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(\rbzero.spi_registers.spi_counter[1] ),
    .B1(_02775_),
    .C1(_02776_),
    .X(_02781_));
 sky130_fd_sc_hd__or3_1 _18702_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .C(_02488_),
    .X(_02782_));
 sky130_fd_sc_hd__o21ai_1 _18703_ (.A1(_02487_),
    .A2(_02488_),
    .B1(\rbzero.spi_registers.spi_counter[2] ),
    .Y(_02783_));
 sky130_fd_sc_hd__a32o_1 _18704_ (.A1(\rbzero.spi_registers.spi_counter[1] ),
    .A2(_02782_),
    .A3(_02783_),
    .B1(_02775_),
    .B2(_02776_),
    .X(_02784_));
 sky130_fd_sc_hd__and2b_1 _18705_ (.A_N(_02781_),
    .B(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__and4bb_1 _18706_ (.A_N(\rbzero.spi_registers.spi_counter[1] ),
    .B_N(_02780_),
    .C(_02770_),
    .D(\rbzero.spi_registers.spi_counter[2] ),
    .X(_02786_));
 sky130_fd_sc_hd__a31oi_1 _18707_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02780_),
    .A3(_02785_),
    .B1(_02786_),
    .Y(_02787_));
 sky130_fd_sc_hd__or2_1 _18708_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(\rbzero.spi_registers.spi_counter[5] ),
    .X(_02788_));
 sky130_fd_sc_hd__a21oi_1 _18709_ (.A1(_02485_),
    .A2(_02773_),
    .B1(_02777_),
    .Y(_02789_));
 sky130_fd_sc_hd__o22a_1 _18710_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_02789_),
    .B1(_02778_),
    .B2(\rbzero.spi_registers.spi_counter[3] ),
    .X(_02790_));
 sky130_fd_sc_hd__a21bo_1 _18711_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_02789_),
    .B1_N(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__a2111o_1 _18712_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(_02778_),
    .B1(_02787_),
    .C1(_02788_),
    .D1(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__a21o_1 _18713_ (.A1(_02771_),
    .A2(_02792_),
    .B1(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02793_));
 sky130_fd_sc_hd__nor2_2 _18714_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_04187_),
    .Y(_02794_));
 sky130_fd_sc_hd__o211a_1 _18715_ (.A1(_02770_),
    .A2(_02772_),
    .B1(_02793_),
    .C1(_02794_),
    .X(_00624_));
 sky130_fd_sc_hd__o21ai_2 _18716_ (.A1(_02772_),
    .A2(_02792_),
    .B1(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__a21oi_1 _18717_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02771_),
    .B1(\rbzero.spi_registers.spi_counter[1] ),
    .Y(_02796_));
 sky130_fd_sc_hd__and3_1 _18718_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .C(_02771_),
    .X(_02797_));
 sky130_fd_sc_hd__nor3_1 _18719_ (.A(_02795_),
    .B(_02796_),
    .C(_02797_),
    .Y(_00625_));
 sky130_fd_sc_hd__xnor2_1 _18720_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__nor2_1 _18721_ (.A(_02795_),
    .B(_02798_),
    .Y(_00626_));
 sky130_fd_sc_hd__a21oi_1 _18722_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(_02797_),
    .B1(\rbzero.spi_registers.spi_counter[3] ),
    .Y(_02799_));
 sky130_fd_sc_hd__and3_1 _18723_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(\rbzero.spi_registers.spi_counter[2] ),
    .C(_02797_),
    .X(_02800_));
 sky130_fd_sc_hd__nor3_1 _18724_ (.A(_02795_),
    .B(_02799_),
    .C(_02800_),
    .Y(_00627_));
 sky130_fd_sc_hd__and2_1 _18725_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__or2_1 _18726_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02800_),
    .X(_02802_));
 sky130_fd_sc_hd__nor3b_1 _18727_ (.A(_02801_),
    .B(_02795_),
    .C_N(_02802_),
    .Y(_00628_));
 sky130_fd_sc_hd__and3_1 _18728_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(\rbzero.spi_registers.spi_counter[4] ),
    .C(_02800_),
    .X(_02803_));
 sky130_fd_sc_hd__o21ai_1 _18729_ (.A1(\rbzero.spi_registers.spi_counter[5] ),
    .A2(_02801_),
    .B1(_02794_),
    .Y(_02804_));
 sky130_fd_sc_hd__nor2_1 _18730_ (.A(_02803_),
    .B(_02804_),
    .Y(_00629_));
 sky130_fd_sc_hd__or2_1 _18731_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(_02803_),
    .X(_02805_));
 sky130_fd_sc_hd__nand2_1 _18732_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(_02803_),
    .Y(_02806_));
 sky130_fd_sc_hd__and3_1 _18733_ (.A(_02794_),
    .B(_02805_),
    .C(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__clkbuf_1 _18734_ (.A(_02807_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_4 _18735_ (.A(_08244_),
    .X(_02808_));
 sky130_fd_sc_hd__and2_1 _18736_ (.A(net56),
    .B(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _18737_ (.A(_02809_),
    .X(_00631_));
 sky130_fd_sc_hd__and2_1 _18738_ (.A(\rbzero.pov.sclk_buffer[0] ),
    .B(_02808_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_1 _18739_ (.A(_02810_),
    .X(_00632_));
 sky130_fd_sc_hd__and2_1 _18740_ (.A(\rbzero.pov.sclk_buffer[1] ),
    .B(_02808_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_1 _18741_ (.A(_02811_),
    .X(_00633_));
 sky130_fd_sc_hd__or4_2 _18742_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(\rbzero.spi_registers.spi_counter[3] ),
    .C(\rbzero.spi_registers.spi_counter[2] ),
    .D(_02788_),
    .X(_02812_));
 sky130_fd_sc_hd__and3_1 _18743_ (.A(_02794_),
    .B(_02771_),
    .C(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__buf_2 _18744_ (.A(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__buf_4 _18745_ (.A(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _18746_ (.A0(_02484_),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__clkbuf_1 _18747_ (.A(_02816_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _18748_ (.A0(_02494_),
    .A1(_02484_),
    .S(_02815_),
    .X(_02817_));
 sky130_fd_sc_hd__clkbuf_1 _18749_ (.A(_02817_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _18750_ (.A0(_02496_),
    .A1(_02494_),
    .S(_02815_),
    .X(_02818_));
 sky130_fd_sc_hd__clkbuf_1 _18751_ (.A(_02818_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _18752_ (.A0(_02498_),
    .A1(_02496_),
    .S(_02815_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _18753_ (.A(_02819_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _18754_ (.A0(_02500_),
    .A1(_02498_),
    .S(_02815_),
    .X(_02820_));
 sky130_fd_sc_hd__clkbuf_1 _18755_ (.A(_02820_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _18756_ (.A0(_02502_),
    .A1(_02500_),
    .S(_02815_),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_1 _18757_ (.A(_02821_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _18758_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(_02502_),
    .S(_02815_),
    .X(_02822_));
 sky130_fd_sc_hd__clkbuf_1 _18759_ (.A(_02822_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _18760_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02815_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_1 _18761_ (.A(_02823_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _18762_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02815_),
    .X(_02824_));
 sky130_fd_sc_hd__clkbuf_1 _18763_ (.A(_02824_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _18764_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02815_),
    .X(_02825_));
 sky130_fd_sc_hd__clkbuf_1 _18765_ (.A(_02825_),
    .X(_00643_));
 sky130_fd_sc_hd__buf_4 _18766_ (.A(_02814_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _18767_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__clkbuf_1 _18768_ (.A(_02827_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _18769_ (.A0(\rbzero.spi_registers.spi_buffer[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02826_),
    .X(_02828_));
 sky130_fd_sc_hd__clkbuf_1 _18770_ (.A(_02828_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _18771_ (.A0(\rbzero.spi_registers.spi_buffer[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_02826_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _18772_ (.A(_02829_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _18773_ (.A0(\rbzero.spi_registers.spi_buffer[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_02826_),
    .X(_02830_));
 sky130_fd_sc_hd__clkbuf_1 _18774_ (.A(_02830_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18775_ (.A0(\rbzero.spi_registers.spi_buffer[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_02826_),
    .X(_02831_));
 sky130_fd_sc_hd__clkbuf_1 _18776_ (.A(_02831_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _18777_ (.A0(\rbzero.spi_registers.spi_buffer[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_02826_),
    .X(_02832_));
 sky130_fd_sc_hd__clkbuf_1 _18778_ (.A(_02832_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18779_ (.A0(\rbzero.spi_registers.spi_buffer[16] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_02826_),
    .X(_02833_));
 sky130_fd_sc_hd__clkbuf_1 _18780_ (.A(_02833_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _18781_ (.A0(\rbzero.spi_registers.spi_buffer[17] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_02826_),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_1 _18782_ (.A(_02834_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _18783_ (.A0(\rbzero.spi_registers.spi_buffer[18] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_02826_),
    .X(_02835_));
 sky130_fd_sc_hd__clkbuf_1 _18784_ (.A(_02835_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _18785_ (.A0(\rbzero.spi_registers.spi_buffer[19] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_02826_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _18786_ (.A(_02836_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18787_ (.A0(\rbzero.spi_registers.spi_buffer[20] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_02814_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _18788_ (.A(_02837_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _18789_ (.A0(\rbzero.spi_registers.spi_buffer[21] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_02814_),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _18790_ (.A(_02838_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _18791_ (.A0(\rbzero.spi_registers.spi_buffer[22] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_02814_),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _18792_ (.A(_02839_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _18793_ (.A0(\rbzero.spi_registers.spi_buffer[23] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_02814_),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _18794_ (.A(_02840_),
    .X(_00657_));
 sky130_fd_sc_hd__nor4_4 _18795_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_04544_),
    .C(_02772_),
    .D(_02812_),
    .Y(_02841_));
 sky130_fd_sc_hd__mux2_1 _18796_ (.A0(\rbzero.spi_registers.spi_cmd[0] ),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _18797_ (.A(_02842_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _18798_ (.A0(_02485_),
    .A1(\rbzero.spi_registers.spi_cmd[0] ),
    .S(_02841_),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _18799_ (.A(_02843_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _18800_ (.A0(_02487_),
    .A1(_02485_),
    .S(_02841_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _18801_ (.A(_02844_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _18802_ (.A0(_02488_),
    .A1(_02487_),
    .S(_02841_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _18803_ (.A(_02845_),
    .X(_00661_));
 sky130_fd_sc_hd__and2_1 _18804_ (.A(net44),
    .B(_02808_),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _18805_ (.A(_02846_),
    .X(_00662_));
 sky130_fd_sc_hd__and2_1 _18806_ (.A(\rbzero.spi_registers.mosi_buffer[0] ),
    .B(_02808_),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _18807_ (.A(_02847_),
    .X(_00663_));
 sky130_fd_sc_hd__and2_1 _18808_ (.A(net43),
    .B(_02808_),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _18809_ (.A(_02848_),
    .X(_00664_));
 sky130_fd_sc_hd__and2_1 _18810_ (.A(\rbzero.spi_registers.ss_buffer[0] ),
    .B(_02808_),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _18811_ (.A(_02849_),
    .X(_00665_));
 sky130_fd_sc_hd__buf_4 _18812_ (.A(_08244_),
    .X(_02850_));
 sky130_fd_sc_hd__and2_1 _18813_ (.A(net46),
    .B(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _18814_ (.A(_02851_),
    .X(_00666_));
 sky130_fd_sc_hd__and2_1 _18815_ (.A(\rbzero.spi_registers.sclk_buffer[0] ),
    .B(_02850_),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _18816_ (.A(_02852_),
    .X(_00667_));
 sky130_fd_sc_hd__and2_1 _18817_ (.A(\rbzero.spi_registers.sclk_buffer[1] ),
    .B(_02850_),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _18818_ (.A(_02853_),
    .X(_00668_));
 sky130_fd_sc_hd__and3_1 _18819_ (.A(_05177_),
    .B(_04775_),
    .C(_04782_),
    .X(_02854_));
 sky130_fd_sc_hd__and2b_2 _18820_ (.A_N(_05746_),
    .B(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__and3_1 _18821_ (.A(\gpout0.vpos[2] ),
    .B(_05745_),
    .C(\gpout0.vpos[0] ),
    .X(_02856_));
 sky130_fd_sc_hd__and3_2 _18822_ (.A(_05739_),
    .B(_02632_),
    .C(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__and4_1 _18823_ (.A(_04817_),
    .B(_05742_),
    .C(_02855_),
    .D(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__buf_6 _18824_ (.A(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__buf_6 _18825_ (.A(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__buf_4 _18826_ (.A(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__nand2_4 _18827_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__and3_1 _18828_ (.A(_05739_),
    .B(_09866_),
    .C(_02856_),
    .X(_02863_));
 sky130_fd_sc_hd__and4_2 _18829_ (.A(_04817_),
    .B(_05742_),
    .C(_02855_),
    .D(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__and2_2 _18830_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__or2_1 _18831_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__buf_4 _18832_ (.A(_08244_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_4 _18833_ (.A(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__o211a_1 _18834_ (.A1(\rbzero.spi_registers.new_other[6] ),
    .A2(_02862_),
    .B1(_02866_),
    .C1(_02868_),
    .X(_00669_));
 sky130_fd_sc_hd__or2_1 _18835_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .B(_02865_),
    .X(_02869_));
 sky130_fd_sc_hd__o211a_1 _18836_ (.A1(net515),
    .A2(_02862_),
    .B1(_02869_),
    .C1(_02868_),
    .X(_00670_));
 sky130_fd_sc_hd__or2_1 _18837_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .B(_02865_),
    .X(_02870_));
 sky130_fd_sc_hd__o211a_1 _18838_ (.A1(net516),
    .A2(_02862_),
    .B1(_02870_),
    .C1(_02868_),
    .X(_00671_));
 sky130_fd_sc_hd__or2_1 _18839_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .B(_02865_),
    .X(_02871_));
 sky130_fd_sc_hd__o211a_1 _18840_ (.A1(\rbzero.spi_registers.new_other[9] ),
    .A2(_02862_),
    .B1(_02871_),
    .C1(_02868_),
    .X(_00672_));
 sky130_fd_sc_hd__or2_1 _18841_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_02865_),
    .X(_02872_));
 sky130_fd_sc_hd__o211a_1 _18842_ (.A1(net513),
    .A2(_02862_),
    .B1(_02872_),
    .C1(_02868_),
    .X(_00673_));
 sky130_fd_sc_hd__or2_1 _18843_ (.A(\rbzero.map_overlay.i_othery[0] ),
    .B(_02865_),
    .X(_02873_));
 sky130_fd_sc_hd__o211a_1 _18844_ (.A1(\rbzero.spi_registers.new_other[0] ),
    .A2(_02862_),
    .B1(_02873_),
    .C1(_02868_),
    .X(_00674_));
 sky130_fd_sc_hd__or2_1 _18845_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(_02865_),
    .X(_02874_));
 sky130_fd_sc_hd__o211a_1 _18846_ (.A1(net517),
    .A2(_02862_),
    .B1(_02874_),
    .C1(_02868_),
    .X(_00675_));
 sky130_fd_sc_hd__or2_1 _18847_ (.A(\rbzero.map_overlay.i_othery[2] ),
    .B(_02865_),
    .X(_02875_));
 sky130_fd_sc_hd__buf_6 _18848_ (.A(_08244_),
    .X(_02876_));
 sky130_fd_sc_hd__buf_2 _18849_ (.A(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__o211a_1 _18850_ (.A1(net519),
    .A2(_02862_),
    .B1(_02875_),
    .C1(_02877_),
    .X(_00676_));
 sky130_fd_sc_hd__or2_1 _18851_ (.A(\rbzero.map_overlay.i_othery[3] ),
    .B(_02865_),
    .X(_02878_));
 sky130_fd_sc_hd__o211a_1 _18852_ (.A1(\rbzero.spi_registers.new_other[3] ),
    .A2(_02862_),
    .B1(_02878_),
    .C1(_02877_),
    .X(_00677_));
 sky130_fd_sc_hd__or2_1 _18853_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .B(_02865_),
    .X(_02879_));
 sky130_fd_sc_hd__o211a_1 _18854_ (.A1(\rbzero.spi_registers.new_other[4] ),
    .A2(_02862_),
    .B1(_02879_),
    .C1(_02877_),
    .X(_00678_));
 sky130_fd_sc_hd__inv_2 _18855_ (.A(\rbzero.spi_registers.got_new_vinf ),
    .Y(_02880_));
 sky130_fd_sc_hd__nand4_4 _18856_ (.A(_04817_),
    .B(_05742_),
    .C(_02855_),
    .D(_02857_),
    .Y(_02881_));
 sky130_fd_sc_hd__a21o_1 _18857_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_02864_),
    .B1(\rbzero.row_render.vinf ),
    .X(_02882_));
 sky130_fd_sc_hd__buf_4 _18858_ (.A(_08245_),
    .X(_02883_));
 sky130_fd_sc_hd__o311a_1 _18859_ (.A1(net514),
    .A2(_02880_),
    .A3(_02881_),
    .B1(_02882_),
    .C1(_02883_),
    .X(_00679_));
 sky130_fd_sc_hd__nand2_2 _18860_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_02860_),
    .Y(_02884_));
 sky130_fd_sc_hd__clkbuf_4 _18861_ (.A(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__and2_1 _18862_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_02864_),
    .X(_02886_));
 sky130_fd_sc_hd__buf_2 _18863_ (.A(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__or2_1 _18864_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__o211a_1 _18865_ (.A1(\rbzero.spi_registers.new_mapd[10] ),
    .A2(_02885_),
    .B1(_02888_),
    .C1(_02877_),
    .X(_00680_));
 sky130_fd_sc_hd__or2_1 _18866_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .B(_02887_),
    .X(_02889_));
 sky130_fd_sc_hd__o211a_1 _18867_ (.A1(\rbzero.spi_registers.new_mapd[11] ),
    .A2(_02885_),
    .B1(_02889_),
    .C1(_02877_),
    .X(_00681_));
 sky130_fd_sc_hd__or2_1 _18868_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_02887_),
    .X(_02890_));
 sky130_fd_sc_hd__o211a_1 _18869_ (.A1(\rbzero.spi_registers.new_mapd[12] ),
    .A2(_02885_),
    .B1(_02890_),
    .C1(_02877_),
    .X(_00682_));
 sky130_fd_sc_hd__or2_1 _18870_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_02887_),
    .X(_02891_));
 sky130_fd_sc_hd__o211a_1 _18871_ (.A1(\rbzero.spi_registers.new_mapd[13] ),
    .A2(_02885_),
    .B1(_02891_),
    .C1(_02877_),
    .X(_00683_));
 sky130_fd_sc_hd__or2_1 _18872_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .B(_02887_),
    .X(_02892_));
 sky130_fd_sc_hd__o211a_1 _18873_ (.A1(\rbzero.spi_registers.new_mapd[14] ),
    .A2(_02885_),
    .B1(_02892_),
    .C1(_02877_),
    .X(_00684_));
 sky130_fd_sc_hd__or2_1 _18874_ (.A(\rbzero.map_overlay.i_mapdx[5] ),
    .B(_02887_),
    .X(_02893_));
 sky130_fd_sc_hd__o211a_1 _18875_ (.A1(\rbzero.spi_registers.new_mapd[15] ),
    .A2(_02885_),
    .B1(_02893_),
    .C1(_02877_),
    .X(_00685_));
 sky130_fd_sc_hd__or2_1 _18876_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(_02887_),
    .X(_02894_));
 sky130_fd_sc_hd__o211a_1 _18877_ (.A1(\rbzero.spi_registers.new_mapd[4] ),
    .A2(_02885_),
    .B1(_02894_),
    .C1(_02877_),
    .X(_00686_));
 sky130_fd_sc_hd__or2_1 _18878_ (.A(\rbzero.map_overlay.i_mapdy[1] ),
    .B(_02887_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_4 _18879_ (.A(_02876_),
    .X(_02896_));
 sky130_fd_sc_hd__o211a_1 _18880_ (.A1(\rbzero.spi_registers.new_mapd[5] ),
    .A2(_02885_),
    .B1(_02895_),
    .C1(_02896_),
    .X(_00687_));
 sky130_fd_sc_hd__or2_1 _18881_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(_02887_),
    .X(_02897_));
 sky130_fd_sc_hd__o211a_1 _18882_ (.A1(\rbzero.spi_registers.new_mapd[6] ),
    .A2(_02885_),
    .B1(_02897_),
    .C1(_02896_),
    .X(_00688_));
 sky130_fd_sc_hd__or2_1 _18883_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(_02887_),
    .X(_02898_));
 sky130_fd_sc_hd__o211a_1 _18884_ (.A1(\rbzero.spi_registers.new_mapd[7] ),
    .A2(_02885_),
    .B1(_02898_),
    .C1(_02896_),
    .X(_00689_));
 sky130_fd_sc_hd__or2_1 _18885_ (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .B(_02886_),
    .X(_02899_));
 sky130_fd_sc_hd__o211a_1 _18886_ (.A1(\rbzero.spi_registers.new_mapd[8] ),
    .A2(_02884_),
    .B1(_02899_),
    .C1(_02896_),
    .X(_00690_));
 sky130_fd_sc_hd__or2_1 _18887_ (.A(\rbzero.map_overlay.i_mapdy[5] ),
    .B(_02886_),
    .X(_02900_));
 sky130_fd_sc_hd__o211a_1 _18888_ (.A1(\rbzero.spi_registers.new_mapd[9] ),
    .A2(_02884_),
    .B1(_02900_),
    .C1(_02896_),
    .X(_00691_));
 sky130_fd_sc_hd__or2_1 _18889_ (.A(\rbzero.mapdxw[0] ),
    .B(_02886_),
    .X(_02901_));
 sky130_fd_sc_hd__o211a_1 _18890_ (.A1(\rbzero.spi_registers.new_mapd[2] ),
    .A2(_02884_),
    .B1(_02901_),
    .C1(_02896_),
    .X(_00692_));
 sky130_fd_sc_hd__or2_1 _18891_ (.A(\rbzero.mapdxw[1] ),
    .B(_02886_),
    .X(_02902_));
 sky130_fd_sc_hd__o211a_1 _18892_ (.A1(\rbzero.spi_registers.new_mapd[3] ),
    .A2(_02884_),
    .B1(_02902_),
    .C1(_02896_),
    .X(_00693_));
 sky130_fd_sc_hd__or2_1 _18893_ (.A(\rbzero.mapdyw[0] ),
    .B(_02886_),
    .X(_02903_));
 sky130_fd_sc_hd__o211a_1 _18894_ (.A1(\rbzero.spi_registers.new_mapd[0] ),
    .A2(_02884_),
    .B1(_02903_),
    .C1(_02896_),
    .X(_00694_));
 sky130_fd_sc_hd__or2_1 _18895_ (.A(\rbzero.mapdyw[1] ),
    .B(_02886_),
    .X(_02904_));
 sky130_fd_sc_hd__o211a_1 _18896_ (.A1(\rbzero.spi_registers.new_mapd[1] ),
    .A2(_02884_),
    .B1(_02904_),
    .C1(_02896_),
    .X(_00695_));
 sky130_fd_sc_hd__nand2_2 _18897_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02861_),
    .Y(_02905_));
 sky130_fd_sc_hd__and2_1 _18898_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_02859_),
    .X(_02906_));
 sky130_fd_sc_hd__or2_1 _18899_ (.A(\rbzero.floor_leak[0] ),
    .B(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__o211a_1 _18900_ (.A1(\rbzero.spi_registers.new_leak[0] ),
    .A2(_02905_),
    .B1(_02907_),
    .C1(_02896_),
    .X(_00696_));
 sky130_fd_sc_hd__or2_1 _18901_ (.A(\rbzero.floor_leak[1] ),
    .B(_02906_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_4 _18902_ (.A(_02876_),
    .X(_02909_));
 sky130_fd_sc_hd__o211a_1 _18903_ (.A1(\rbzero.spi_registers.new_leak[1] ),
    .A2(_02905_),
    .B1(_02908_),
    .C1(_02909_),
    .X(_00697_));
 sky130_fd_sc_hd__or2_1 _18904_ (.A(\rbzero.floor_leak[2] ),
    .B(_02906_),
    .X(_02910_));
 sky130_fd_sc_hd__o211a_1 _18905_ (.A1(\rbzero.spi_registers.new_leak[2] ),
    .A2(_02905_),
    .B1(_02910_),
    .C1(_02909_),
    .X(_00698_));
 sky130_fd_sc_hd__or2_1 _18906_ (.A(\rbzero.floor_leak[3] ),
    .B(_02906_),
    .X(_02911_));
 sky130_fd_sc_hd__o211a_1 _18907_ (.A1(\rbzero.spi_registers.new_leak[3] ),
    .A2(_02905_),
    .B1(_02911_),
    .C1(_02909_),
    .X(_00699_));
 sky130_fd_sc_hd__or2_1 _18908_ (.A(\rbzero.floor_leak[4] ),
    .B(_02906_),
    .X(_02912_));
 sky130_fd_sc_hd__o211a_1 _18909_ (.A1(\rbzero.spi_registers.new_leak[4] ),
    .A2(_02905_),
    .B1(_02912_),
    .C1(_02909_),
    .X(_00700_));
 sky130_fd_sc_hd__or2_1 _18910_ (.A(\rbzero.floor_leak[5] ),
    .B(_02906_),
    .X(_02913_));
 sky130_fd_sc_hd__o211a_1 _18911_ (.A1(\rbzero.spi_registers.new_leak[5] ),
    .A2(_02905_),
    .B1(_02913_),
    .C1(_02909_),
    .X(_00701_));
 sky130_fd_sc_hd__nand2_2 _18912_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_02861_),
    .Y(_02914_));
 sky130_fd_sc_hd__buf_6 _18913_ (.A(_04544_),
    .X(_02915_));
 sky130_fd_sc_hd__a31o_1 _18914_ (.A1(\rbzero.spi_registers.new_sky[0] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02861_),
    .B1(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__a21o_1 _18915_ (.A1(\rbzero.color_sky[0] ),
    .A2(_02914_),
    .B1(_02916_),
    .X(_00702_));
 sky130_fd_sc_hd__and2_1 _18916_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_02860_),
    .X(_02917_));
 sky130_fd_sc_hd__or2_1 _18917_ (.A(\rbzero.color_sky[1] ),
    .B(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__o211a_1 _18918_ (.A1(\rbzero.spi_registers.new_sky[1] ),
    .A2(_02914_),
    .B1(_02918_),
    .C1(_02909_),
    .X(_00703_));
 sky130_fd_sc_hd__a31o_1 _18919_ (.A1(\rbzero.spi_registers.new_sky[2] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02861_),
    .B1(_04545_),
    .X(_02919_));
 sky130_fd_sc_hd__a21o_1 _18920_ (.A1(\rbzero.color_sky[2] ),
    .A2(_02914_),
    .B1(_02919_),
    .X(_00704_));
 sky130_fd_sc_hd__or2_1 _18921_ (.A(\rbzero.color_sky[3] ),
    .B(_02917_),
    .X(_02920_));
 sky130_fd_sc_hd__o211a_1 _18922_ (.A1(\rbzero.spi_registers.new_sky[3] ),
    .A2(_02914_),
    .B1(_02920_),
    .C1(_02909_),
    .X(_00705_));
 sky130_fd_sc_hd__a31o_1 _18923_ (.A1(\rbzero.spi_registers.new_sky[4] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_02861_),
    .B1(_04545_),
    .X(_02921_));
 sky130_fd_sc_hd__a21o_1 _18924_ (.A1(\rbzero.color_sky[4] ),
    .A2(_02914_),
    .B1(_02921_),
    .X(_00706_));
 sky130_fd_sc_hd__or2_1 _18925_ (.A(\rbzero.color_sky[5] ),
    .B(_02917_),
    .X(_02922_));
 sky130_fd_sc_hd__o211a_1 _18926_ (.A1(\rbzero.spi_registers.new_sky[5] ),
    .A2(_02914_),
    .B1(_02922_),
    .C1(_02909_),
    .X(_00707_));
 sky130_fd_sc_hd__buf_4 _18927_ (.A(_02860_),
    .X(_02923_));
 sky130_fd_sc_hd__nand2_2 _18928_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__and2_1 _18929_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_02860_),
    .X(_02925_));
 sky130_fd_sc_hd__or2_1 _18930_ (.A(\rbzero.color_floor[0] ),
    .B(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__o211a_1 _18931_ (.A1(\rbzero.spi_registers.new_floor[0] ),
    .A2(_02924_),
    .B1(_02926_),
    .C1(_02909_),
    .X(_00708_));
 sky130_fd_sc_hd__a31o_1 _18932_ (.A1(\rbzero.spi_registers.new_floor[1] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02861_),
    .B1(_04545_),
    .X(_02927_));
 sky130_fd_sc_hd__a21o_1 _18933_ (.A1(\rbzero.color_floor[1] ),
    .A2(_02924_),
    .B1(_02927_),
    .X(_00709_));
 sky130_fd_sc_hd__or2_1 _18934_ (.A(\rbzero.color_floor[2] ),
    .B(_02925_),
    .X(_02928_));
 sky130_fd_sc_hd__o211a_1 _18935_ (.A1(\rbzero.spi_registers.new_floor[2] ),
    .A2(_02924_),
    .B1(_02928_),
    .C1(_02909_),
    .X(_00710_));
 sky130_fd_sc_hd__a31o_1 _18936_ (.A1(\rbzero.spi_registers.new_floor[3] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02861_),
    .B1(_04545_),
    .X(_02929_));
 sky130_fd_sc_hd__a21o_1 _18937_ (.A1(\rbzero.color_floor[3] ),
    .A2(_02924_),
    .B1(_02929_),
    .X(_00711_));
 sky130_fd_sc_hd__or2_1 _18938_ (.A(\rbzero.color_floor[4] ),
    .B(_02925_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_4 _18939_ (.A(_02876_),
    .X(_02931_));
 sky130_fd_sc_hd__o211a_1 _18940_ (.A1(\rbzero.spi_registers.new_floor[4] ),
    .A2(_02924_),
    .B1(_02930_),
    .C1(_02931_),
    .X(_00712_));
 sky130_fd_sc_hd__a31o_1 _18941_ (.A1(\rbzero.spi_registers.new_floor[5] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_02861_),
    .B1(_04545_),
    .X(_02932_));
 sky130_fd_sc_hd__a21o_1 _18942_ (.A1(\rbzero.color_floor[5] ),
    .A2(_02924_),
    .B1(_02932_),
    .X(_00713_));
 sky130_fd_sc_hd__nand2_2 _18943_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02861_),
    .Y(_02933_));
 sky130_fd_sc_hd__and2_1 _18944_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_02859_),
    .X(_02934_));
 sky130_fd_sc_hd__or2_1 _18945_ (.A(\rbzero.spi_registers.vshift[0] ),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__o211a_1 _18946_ (.A1(\rbzero.spi_registers.new_vshift[0] ),
    .A2(_02933_),
    .B1(_02935_),
    .C1(_02931_),
    .X(_00714_));
 sky130_fd_sc_hd__or2_1 _18947_ (.A(\rbzero.spi_registers.vshift[1] ),
    .B(_02934_),
    .X(_02936_));
 sky130_fd_sc_hd__o211a_1 _18948_ (.A1(\rbzero.spi_registers.new_vshift[1] ),
    .A2(_02933_),
    .B1(_02936_),
    .C1(_02931_),
    .X(_00715_));
 sky130_fd_sc_hd__or2_1 _18949_ (.A(\rbzero.spi_registers.vshift[2] ),
    .B(_02934_),
    .X(_02937_));
 sky130_fd_sc_hd__o211a_1 _18950_ (.A1(\rbzero.spi_registers.new_vshift[2] ),
    .A2(_02933_),
    .B1(_02937_),
    .C1(_02931_),
    .X(_00716_));
 sky130_fd_sc_hd__or2_1 _18951_ (.A(\rbzero.spi_registers.vshift[3] ),
    .B(_02934_),
    .X(_02938_));
 sky130_fd_sc_hd__o211a_1 _18952_ (.A1(\rbzero.spi_registers.new_vshift[3] ),
    .A2(_02933_),
    .B1(_02938_),
    .C1(_02931_),
    .X(_00717_));
 sky130_fd_sc_hd__or2_1 _18953_ (.A(\rbzero.spi_registers.vshift[4] ),
    .B(_02934_),
    .X(_02939_));
 sky130_fd_sc_hd__o211a_1 _18954_ (.A1(\rbzero.spi_registers.new_vshift[4] ),
    .A2(_02933_),
    .B1(_02939_),
    .C1(_02931_),
    .X(_00718_));
 sky130_fd_sc_hd__or2_1 _18955_ (.A(\rbzero.spi_registers.vshift[5] ),
    .B(_02934_),
    .X(_02940_));
 sky130_fd_sc_hd__o211a_1 _18956_ (.A1(\rbzero.spi_registers.new_vshift[5] ),
    .A2(_02933_),
    .B1(_02940_),
    .C1(_02931_),
    .X(_00719_));
 sky130_fd_sc_hd__nand2_2 _18957_ (.A(\rbzero.spi_registers.got_new_texadd0 ),
    .B(_02860_),
    .Y(_02941_));
 sky130_fd_sc_hd__clkbuf_4 _18958_ (.A(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__and2_1 _18959_ (.A(\rbzero.spi_registers.got_new_texadd0 ),
    .B(_02864_),
    .X(_02943_));
 sky130_fd_sc_hd__buf_2 _18960_ (.A(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__or2_1 _18961_ (.A(\rbzero.spi_registers.texadd0[0] ),
    .B(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__o211a_1 _18962_ (.A1(\rbzero.spi_registers.new_texadd0[0] ),
    .A2(_02942_),
    .B1(_02945_),
    .C1(_02931_),
    .X(_00720_));
 sky130_fd_sc_hd__or2_1 _18963_ (.A(\rbzero.spi_registers.texadd0[1] ),
    .B(_02944_),
    .X(_02946_));
 sky130_fd_sc_hd__o211a_1 _18964_ (.A1(\rbzero.spi_registers.new_texadd0[1] ),
    .A2(_02942_),
    .B1(_02946_),
    .C1(_02931_),
    .X(_00721_));
 sky130_fd_sc_hd__or2_1 _18965_ (.A(\rbzero.spi_registers.texadd0[2] ),
    .B(_02944_),
    .X(_02947_));
 sky130_fd_sc_hd__o211a_1 _18966_ (.A1(\rbzero.spi_registers.new_texadd0[2] ),
    .A2(_02942_),
    .B1(_02947_),
    .C1(_02931_),
    .X(_00722_));
 sky130_fd_sc_hd__or2_1 _18967_ (.A(\rbzero.spi_registers.texadd0[3] ),
    .B(_02944_),
    .X(_02948_));
 sky130_fd_sc_hd__clkbuf_4 _18968_ (.A(_02876_),
    .X(_02949_));
 sky130_fd_sc_hd__o211a_1 _18969_ (.A1(\rbzero.spi_registers.new_texadd0[3] ),
    .A2(_02942_),
    .B1(_02948_),
    .C1(_02949_),
    .X(_00723_));
 sky130_fd_sc_hd__or2_1 _18970_ (.A(\rbzero.spi_registers.texadd0[4] ),
    .B(_02944_),
    .X(_02950_));
 sky130_fd_sc_hd__o211a_1 _18971_ (.A1(\rbzero.spi_registers.new_texadd0[4] ),
    .A2(_02942_),
    .B1(_02950_),
    .C1(_02949_),
    .X(_00724_));
 sky130_fd_sc_hd__or2_1 _18972_ (.A(\rbzero.spi_registers.texadd0[5] ),
    .B(_02944_),
    .X(_02951_));
 sky130_fd_sc_hd__o211a_1 _18973_ (.A1(\rbzero.spi_registers.new_texadd0[5] ),
    .A2(_02942_),
    .B1(_02951_),
    .C1(_02949_),
    .X(_00725_));
 sky130_fd_sc_hd__or2_1 _18974_ (.A(\rbzero.spi_registers.texadd0[6] ),
    .B(_02944_),
    .X(_02952_));
 sky130_fd_sc_hd__o211a_1 _18975_ (.A1(\rbzero.spi_registers.new_texadd0[6] ),
    .A2(_02942_),
    .B1(_02952_),
    .C1(_02949_),
    .X(_00726_));
 sky130_fd_sc_hd__or2_1 _18976_ (.A(\rbzero.spi_registers.texadd0[7] ),
    .B(_02944_),
    .X(_02953_));
 sky130_fd_sc_hd__o211a_1 _18977_ (.A1(\rbzero.spi_registers.new_texadd0[7] ),
    .A2(_02942_),
    .B1(_02953_),
    .C1(_02949_),
    .X(_00727_));
 sky130_fd_sc_hd__or2_1 _18978_ (.A(\rbzero.spi_registers.texadd0[8] ),
    .B(_02944_),
    .X(_02954_));
 sky130_fd_sc_hd__o211a_1 _18979_ (.A1(\rbzero.spi_registers.new_texadd0[8] ),
    .A2(_02942_),
    .B1(_02954_),
    .C1(_02949_),
    .X(_00728_));
 sky130_fd_sc_hd__or2_1 _18980_ (.A(\rbzero.spi_registers.texadd0[9] ),
    .B(_02944_),
    .X(_02955_));
 sky130_fd_sc_hd__o211a_1 _18981_ (.A1(\rbzero.spi_registers.new_texadd0[9] ),
    .A2(_02942_),
    .B1(_02955_),
    .C1(_02949_),
    .X(_00729_));
 sky130_fd_sc_hd__clkbuf_4 _18982_ (.A(_02941_),
    .X(_02956_));
 sky130_fd_sc_hd__buf_2 _18983_ (.A(_02943_),
    .X(_02957_));
 sky130_fd_sc_hd__or2_1 _18984_ (.A(\rbzero.spi_registers.texadd0[10] ),
    .B(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__o211a_1 _18985_ (.A1(\rbzero.spi_registers.new_texadd0[10] ),
    .A2(_02956_),
    .B1(_02958_),
    .C1(_02949_),
    .X(_00730_));
 sky130_fd_sc_hd__or2_1 _18986_ (.A(\rbzero.spi_registers.texadd0[11] ),
    .B(_02957_),
    .X(_02959_));
 sky130_fd_sc_hd__o211a_1 _18987_ (.A1(\rbzero.spi_registers.new_texadd0[11] ),
    .A2(_02956_),
    .B1(_02959_),
    .C1(_02949_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_1 _18988_ (.A(\rbzero.spi_registers.texadd0[12] ),
    .B(_02957_),
    .X(_02960_));
 sky130_fd_sc_hd__o211a_1 _18989_ (.A1(\rbzero.spi_registers.new_texadd0[12] ),
    .A2(_02956_),
    .B1(_02960_),
    .C1(_02949_),
    .X(_00732_));
 sky130_fd_sc_hd__or2_1 _18990_ (.A(\rbzero.spi_registers.texadd0[13] ),
    .B(_02957_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_4 _18991_ (.A(_02876_),
    .X(_02962_));
 sky130_fd_sc_hd__o211a_1 _18992_ (.A1(\rbzero.spi_registers.new_texadd0[13] ),
    .A2(_02956_),
    .B1(_02961_),
    .C1(_02962_),
    .X(_00733_));
 sky130_fd_sc_hd__or2_1 _18993_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_02957_),
    .X(_02963_));
 sky130_fd_sc_hd__o211a_1 _18994_ (.A1(\rbzero.spi_registers.new_texadd0[14] ),
    .A2(_02956_),
    .B1(_02963_),
    .C1(_02962_),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _18995_ (.A(\rbzero.spi_registers.texadd0[15] ),
    .B(_02957_),
    .X(_02964_));
 sky130_fd_sc_hd__o211a_1 _18996_ (.A1(\rbzero.spi_registers.new_texadd0[15] ),
    .A2(_02956_),
    .B1(_02964_),
    .C1(_02962_),
    .X(_00735_));
 sky130_fd_sc_hd__or2_1 _18997_ (.A(\rbzero.spi_registers.texadd0[16] ),
    .B(_02957_),
    .X(_02965_));
 sky130_fd_sc_hd__o211a_1 _18998_ (.A1(\rbzero.spi_registers.new_texadd0[16] ),
    .A2(_02956_),
    .B1(_02965_),
    .C1(_02962_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _18999_ (.A(\rbzero.spi_registers.texadd0[17] ),
    .B(_02957_),
    .X(_02966_));
 sky130_fd_sc_hd__o211a_1 _19000_ (.A1(\rbzero.spi_registers.new_texadd0[17] ),
    .A2(_02956_),
    .B1(_02966_),
    .C1(_02962_),
    .X(_00737_));
 sky130_fd_sc_hd__or2_1 _19001_ (.A(\rbzero.spi_registers.texadd0[18] ),
    .B(_02957_),
    .X(_02967_));
 sky130_fd_sc_hd__o211a_1 _19002_ (.A1(\rbzero.spi_registers.new_texadd0[18] ),
    .A2(_02956_),
    .B1(_02967_),
    .C1(_02962_),
    .X(_00738_));
 sky130_fd_sc_hd__or2_1 _19003_ (.A(\rbzero.spi_registers.texadd0[19] ),
    .B(_02957_),
    .X(_02968_));
 sky130_fd_sc_hd__o211a_1 _19004_ (.A1(\rbzero.spi_registers.new_texadd0[19] ),
    .A2(_02956_),
    .B1(_02968_),
    .C1(_02962_),
    .X(_00739_));
 sky130_fd_sc_hd__or2_1 _19005_ (.A(\rbzero.spi_registers.texadd0[20] ),
    .B(_02943_),
    .X(_02969_));
 sky130_fd_sc_hd__o211a_1 _19006_ (.A1(\rbzero.spi_registers.new_texadd0[20] ),
    .A2(_02941_),
    .B1(_02969_),
    .C1(_02962_),
    .X(_00740_));
 sky130_fd_sc_hd__or2_1 _19007_ (.A(\rbzero.spi_registers.texadd0[21] ),
    .B(_02943_),
    .X(_02970_));
 sky130_fd_sc_hd__o211a_1 _19008_ (.A1(\rbzero.spi_registers.new_texadd0[21] ),
    .A2(_02941_),
    .B1(_02970_),
    .C1(_02962_),
    .X(_00741_));
 sky130_fd_sc_hd__or2_1 _19009_ (.A(\rbzero.spi_registers.texadd0[22] ),
    .B(_02943_),
    .X(_02971_));
 sky130_fd_sc_hd__o211a_1 _19010_ (.A1(\rbzero.spi_registers.new_texadd0[22] ),
    .A2(_02941_),
    .B1(_02971_),
    .C1(_02962_),
    .X(_00742_));
 sky130_fd_sc_hd__or2_1 _19011_ (.A(\rbzero.spi_registers.texadd0[23] ),
    .B(_02943_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_4 _19012_ (.A(_08244_),
    .X(_02973_));
 sky130_fd_sc_hd__clkbuf_4 _19013_ (.A(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__o211a_1 _19014_ (.A1(\rbzero.spi_registers.new_texadd0[23] ),
    .A2(_02941_),
    .B1(_02972_),
    .C1(_02974_),
    .X(_00743_));
 sky130_fd_sc_hd__nand2_2 _19015_ (.A(\rbzero.spi_registers.got_new_texadd1 ),
    .B(_02860_),
    .Y(_02975_));
 sky130_fd_sc_hd__clkbuf_4 _19016_ (.A(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__and2_2 _19017_ (.A(\rbzero.spi_registers.got_new_texadd1 ),
    .B(_02864_),
    .X(_02977_));
 sky130_fd_sc_hd__buf_2 _19018_ (.A(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__or2_1 _19019_ (.A(\rbzero.spi_registers.texadd1[0] ),
    .B(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__o211a_1 _19020_ (.A1(\rbzero.spi_registers.new_texadd1[0] ),
    .A2(_02976_),
    .B1(_02979_),
    .C1(_02974_),
    .X(_00744_));
 sky130_fd_sc_hd__or2_1 _19021_ (.A(\rbzero.spi_registers.texadd1[1] ),
    .B(_02978_),
    .X(_02980_));
 sky130_fd_sc_hd__o211a_1 _19022_ (.A1(\rbzero.spi_registers.new_texadd1[1] ),
    .A2(_02976_),
    .B1(_02980_),
    .C1(_02974_),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _19023_ (.A(\rbzero.spi_registers.texadd1[2] ),
    .B(_02978_),
    .X(_02981_));
 sky130_fd_sc_hd__o211a_1 _19024_ (.A1(\rbzero.spi_registers.new_texadd1[2] ),
    .A2(_02976_),
    .B1(_02981_),
    .C1(_02974_),
    .X(_00746_));
 sky130_fd_sc_hd__or2_1 _19025_ (.A(\rbzero.spi_registers.texadd1[3] ),
    .B(_02978_),
    .X(_02982_));
 sky130_fd_sc_hd__o211a_1 _19026_ (.A1(\rbzero.spi_registers.new_texadd1[3] ),
    .A2(_02976_),
    .B1(_02982_),
    .C1(_02974_),
    .X(_00747_));
 sky130_fd_sc_hd__or2_1 _19027_ (.A(\rbzero.spi_registers.texadd1[4] ),
    .B(_02978_),
    .X(_02983_));
 sky130_fd_sc_hd__o211a_1 _19028_ (.A1(\rbzero.spi_registers.new_texadd1[4] ),
    .A2(_02976_),
    .B1(_02983_),
    .C1(_02974_),
    .X(_00748_));
 sky130_fd_sc_hd__or2_1 _19029_ (.A(\rbzero.spi_registers.texadd1[5] ),
    .B(_02978_),
    .X(_02984_));
 sky130_fd_sc_hd__o211a_1 _19030_ (.A1(\rbzero.spi_registers.new_texadd1[5] ),
    .A2(_02976_),
    .B1(_02984_),
    .C1(_02974_),
    .X(_00749_));
 sky130_fd_sc_hd__or2_1 _19031_ (.A(\rbzero.spi_registers.texadd1[6] ),
    .B(_02978_),
    .X(_02985_));
 sky130_fd_sc_hd__o211a_1 _19032_ (.A1(\rbzero.spi_registers.new_texadd1[6] ),
    .A2(_02976_),
    .B1(_02985_),
    .C1(_02974_),
    .X(_00750_));
 sky130_fd_sc_hd__or2_1 _19033_ (.A(\rbzero.spi_registers.texadd1[7] ),
    .B(_02978_),
    .X(_02986_));
 sky130_fd_sc_hd__o211a_1 _19034_ (.A1(\rbzero.spi_registers.new_texadd1[7] ),
    .A2(_02976_),
    .B1(_02986_),
    .C1(_02974_),
    .X(_00751_));
 sky130_fd_sc_hd__or2_1 _19035_ (.A(\rbzero.spi_registers.texadd1[8] ),
    .B(_02978_),
    .X(_02987_));
 sky130_fd_sc_hd__o211a_1 _19036_ (.A1(\rbzero.spi_registers.new_texadd1[8] ),
    .A2(_02976_),
    .B1(_02987_),
    .C1(_02974_),
    .X(_00752_));
 sky130_fd_sc_hd__or2_1 _19037_ (.A(\rbzero.spi_registers.texadd1[9] ),
    .B(_02978_),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_4 _19038_ (.A(_02973_),
    .X(_02989_));
 sky130_fd_sc_hd__o211a_1 _19039_ (.A1(\rbzero.spi_registers.new_texadd1[9] ),
    .A2(_02976_),
    .B1(_02988_),
    .C1(_02989_),
    .X(_00753_));
 sky130_fd_sc_hd__clkbuf_4 _19040_ (.A(_02975_),
    .X(_02990_));
 sky130_fd_sc_hd__buf_2 _19041_ (.A(_02977_),
    .X(_02991_));
 sky130_fd_sc_hd__or2_1 _19042_ (.A(\rbzero.spi_registers.texadd1[10] ),
    .B(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__o211a_1 _19043_ (.A1(\rbzero.spi_registers.new_texadd1[10] ),
    .A2(_02990_),
    .B1(_02992_),
    .C1(_02989_),
    .X(_00754_));
 sky130_fd_sc_hd__or2_1 _19044_ (.A(\rbzero.spi_registers.texadd1[11] ),
    .B(_02991_),
    .X(_02993_));
 sky130_fd_sc_hd__o211a_1 _19045_ (.A1(\rbzero.spi_registers.new_texadd1[11] ),
    .A2(_02990_),
    .B1(_02993_),
    .C1(_02989_),
    .X(_00755_));
 sky130_fd_sc_hd__or2_1 _19046_ (.A(\rbzero.spi_registers.texadd1[12] ),
    .B(_02991_),
    .X(_02994_));
 sky130_fd_sc_hd__o211a_1 _19047_ (.A1(\rbzero.spi_registers.new_texadd1[12] ),
    .A2(_02990_),
    .B1(_02994_),
    .C1(_02989_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _19048_ (.A(\rbzero.spi_registers.texadd1[13] ),
    .B(_02991_),
    .X(_02995_));
 sky130_fd_sc_hd__o211a_1 _19049_ (.A1(\rbzero.spi_registers.new_texadd1[13] ),
    .A2(_02990_),
    .B1(_02995_),
    .C1(_02989_),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _19050_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .B(_02991_),
    .X(_02996_));
 sky130_fd_sc_hd__o211a_1 _19051_ (.A1(\rbzero.spi_registers.new_texadd1[14] ),
    .A2(_02990_),
    .B1(_02996_),
    .C1(_02989_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _19052_ (.A(\rbzero.spi_registers.texadd1[15] ),
    .B(_02991_),
    .X(_02997_));
 sky130_fd_sc_hd__o211a_1 _19053_ (.A1(\rbzero.spi_registers.new_texadd1[15] ),
    .A2(_02990_),
    .B1(_02997_),
    .C1(_02989_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _19054_ (.A(\rbzero.spi_registers.texadd1[16] ),
    .B(_02991_),
    .X(_02998_));
 sky130_fd_sc_hd__o211a_1 _19055_ (.A1(\rbzero.spi_registers.new_texadd1[16] ),
    .A2(_02990_),
    .B1(_02998_),
    .C1(_02989_),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _19056_ (.A(\rbzero.spi_registers.texadd1[17] ),
    .B(_02991_),
    .X(_02999_));
 sky130_fd_sc_hd__o211a_1 _19057_ (.A1(\rbzero.spi_registers.new_texadd1[17] ),
    .A2(_02990_),
    .B1(_02999_),
    .C1(_02989_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _19058_ (.A(\rbzero.spi_registers.texadd1[18] ),
    .B(_02991_),
    .X(_03000_));
 sky130_fd_sc_hd__o211a_1 _19059_ (.A1(\rbzero.spi_registers.new_texadd1[18] ),
    .A2(_02990_),
    .B1(_03000_),
    .C1(_02989_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _19060_ (.A(\rbzero.spi_registers.texadd1[19] ),
    .B(_02991_),
    .X(_03001_));
 sky130_fd_sc_hd__buf_4 _19061_ (.A(_02973_),
    .X(_03002_));
 sky130_fd_sc_hd__o211a_1 _19062_ (.A1(\rbzero.spi_registers.new_texadd1[19] ),
    .A2(_02990_),
    .B1(_03001_),
    .C1(_03002_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _19063_ (.A(\rbzero.spi_registers.texadd1[20] ),
    .B(_02977_),
    .X(_03003_));
 sky130_fd_sc_hd__o211a_1 _19064_ (.A1(\rbzero.spi_registers.new_texadd1[20] ),
    .A2(_02975_),
    .B1(_03003_),
    .C1(_03002_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _19065_ (.A(\rbzero.spi_registers.texadd1[21] ),
    .B(_02977_),
    .X(_03004_));
 sky130_fd_sc_hd__o211a_1 _19066_ (.A1(\rbzero.spi_registers.new_texadd1[21] ),
    .A2(_02975_),
    .B1(_03004_),
    .C1(_03002_),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _19067_ (.A(\rbzero.spi_registers.texadd1[22] ),
    .B(_02977_),
    .X(_03005_));
 sky130_fd_sc_hd__o211a_1 _19068_ (.A1(\rbzero.spi_registers.new_texadd1[22] ),
    .A2(_02975_),
    .B1(_03005_),
    .C1(_03002_),
    .X(_00766_));
 sky130_fd_sc_hd__or2_1 _19069_ (.A(\rbzero.spi_registers.texadd1[23] ),
    .B(_02977_),
    .X(_03006_));
 sky130_fd_sc_hd__o211a_1 _19070_ (.A1(\rbzero.spi_registers.new_texadd1[23] ),
    .A2(_02975_),
    .B1(_03006_),
    .C1(_03002_),
    .X(_00767_));
 sky130_fd_sc_hd__nand2_4 _19071_ (.A(\rbzero.spi_registers.got_new_texadd2 ),
    .B(_02860_),
    .Y(_03007_));
 sky130_fd_sc_hd__clkbuf_4 _19072_ (.A(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__and2_2 _19073_ (.A(\rbzero.spi_registers.got_new_texadd2 ),
    .B(_02864_),
    .X(_03009_));
 sky130_fd_sc_hd__buf_2 _19074_ (.A(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__or2_1 _19075_ (.A(\rbzero.spi_registers.texadd2[0] ),
    .B(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__o211a_1 _19076_ (.A1(\rbzero.spi_registers.new_texadd2[0] ),
    .A2(_03008_),
    .B1(_03011_),
    .C1(_03002_),
    .X(_00768_));
 sky130_fd_sc_hd__or2_1 _19077_ (.A(\rbzero.spi_registers.texadd2[1] ),
    .B(_03010_),
    .X(_03012_));
 sky130_fd_sc_hd__o211a_1 _19078_ (.A1(\rbzero.spi_registers.new_texadd2[1] ),
    .A2(_03008_),
    .B1(_03012_),
    .C1(_03002_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _19079_ (.A(\rbzero.spi_registers.texadd2[2] ),
    .B(_03010_),
    .X(_03013_));
 sky130_fd_sc_hd__o211a_1 _19080_ (.A1(\rbzero.spi_registers.new_texadd2[2] ),
    .A2(_03008_),
    .B1(_03013_),
    .C1(_03002_),
    .X(_00770_));
 sky130_fd_sc_hd__or2_1 _19081_ (.A(\rbzero.spi_registers.texadd2[3] ),
    .B(_03010_),
    .X(_03014_));
 sky130_fd_sc_hd__o211a_1 _19082_ (.A1(\rbzero.spi_registers.new_texadd2[3] ),
    .A2(_03008_),
    .B1(_03014_),
    .C1(_03002_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _19083_ (.A(\rbzero.spi_registers.texadd2[4] ),
    .B(_03010_),
    .X(_03015_));
 sky130_fd_sc_hd__o211a_1 _19084_ (.A1(\rbzero.spi_registers.new_texadd2[4] ),
    .A2(_03008_),
    .B1(_03015_),
    .C1(_03002_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _19085_ (.A(\rbzero.spi_registers.texadd2[5] ),
    .B(_03010_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_4 _19086_ (.A(_02973_),
    .X(_03017_));
 sky130_fd_sc_hd__o211a_1 _19087_ (.A1(\rbzero.spi_registers.new_texadd2[5] ),
    .A2(_03008_),
    .B1(_03016_),
    .C1(_03017_),
    .X(_00773_));
 sky130_fd_sc_hd__or2_1 _19088_ (.A(\rbzero.spi_registers.texadd2[6] ),
    .B(_03010_),
    .X(_03018_));
 sky130_fd_sc_hd__o211a_1 _19089_ (.A1(\rbzero.spi_registers.new_texadd2[6] ),
    .A2(_03008_),
    .B1(_03018_),
    .C1(_03017_),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _19090_ (.A(\rbzero.spi_registers.texadd2[7] ),
    .B(_03010_),
    .X(_03019_));
 sky130_fd_sc_hd__o211a_1 _19091_ (.A1(\rbzero.spi_registers.new_texadd2[7] ),
    .A2(_03008_),
    .B1(_03019_),
    .C1(_03017_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _19092_ (.A(\rbzero.spi_registers.texadd2[8] ),
    .B(_03010_),
    .X(_03020_));
 sky130_fd_sc_hd__o211a_1 _19093_ (.A1(\rbzero.spi_registers.new_texadd2[8] ),
    .A2(_03008_),
    .B1(_03020_),
    .C1(_03017_),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _19094_ (.A(\rbzero.spi_registers.texadd2[9] ),
    .B(_03010_),
    .X(_03021_));
 sky130_fd_sc_hd__o211a_1 _19095_ (.A1(\rbzero.spi_registers.new_texadd2[9] ),
    .A2(_03008_),
    .B1(_03021_),
    .C1(_03017_),
    .X(_00777_));
 sky130_fd_sc_hd__clkbuf_4 _19096_ (.A(_03007_),
    .X(_03022_));
 sky130_fd_sc_hd__buf_2 _19097_ (.A(_03009_),
    .X(_03023_));
 sky130_fd_sc_hd__or2_1 _19098_ (.A(\rbzero.spi_registers.texadd2[10] ),
    .B(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__o211a_1 _19099_ (.A1(\rbzero.spi_registers.new_texadd2[10] ),
    .A2(_03022_),
    .B1(_03024_),
    .C1(_03017_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _19100_ (.A(\rbzero.spi_registers.texadd2[11] ),
    .B(_03023_),
    .X(_03025_));
 sky130_fd_sc_hd__o211a_1 _19101_ (.A1(\rbzero.spi_registers.new_texadd2[11] ),
    .A2(_03022_),
    .B1(_03025_),
    .C1(_03017_),
    .X(_00779_));
 sky130_fd_sc_hd__or2_1 _19102_ (.A(\rbzero.spi_registers.texadd2[12] ),
    .B(_03023_),
    .X(_03026_));
 sky130_fd_sc_hd__o211a_1 _19103_ (.A1(\rbzero.spi_registers.new_texadd2[12] ),
    .A2(_03022_),
    .B1(_03026_),
    .C1(_03017_),
    .X(_00780_));
 sky130_fd_sc_hd__or2_1 _19104_ (.A(\rbzero.spi_registers.texadd2[13] ),
    .B(_03023_),
    .X(_03027_));
 sky130_fd_sc_hd__o211a_1 _19105_ (.A1(\rbzero.spi_registers.new_texadd2[13] ),
    .A2(_03022_),
    .B1(_03027_),
    .C1(_03017_),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _19106_ (.A(\rbzero.spi_registers.texadd2[14] ),
    .B(_03023_),
    .X(_03028_));
 sky130_fd_sc_hd__o211a_1 _19107_ (.A1(\rbzero.spi_registers.new_texadd2[14] ),
    .A2(_03022_),
    .B1(_03028_),
    .C1(_03017_),
    .X(_00782_));
 sky130_fd_sc_hd__or2_1 _19108_ (.A(\rbzero.spi_registers.texadd2[15] ),
    .B(_03023_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_4 _19109_ (.A(_02973_),
    .X(_03030_));
 sky130_fd_sc_hd__o211a_1 _19110_ (.A1(\rbzero.spi_registers.new_texadd2[15] ),
    .A2(_03022_),
    .B1(_03029_),
    .C1(_03030_),
    .X(_00783_));
 sky130_fd_sc_hd__or2_1 _19111_ (.A(\rbzero.spi_registers.texadd2[16] ),
    .B(_03023_),
    .X(_03031_));
 sky130_fd_sc_hd__o211a_1 _19112_ (.A1(\rbzero.spi_registers.new_texadd2[16] ),
    .A2(_03022_),
    .B1(_03031_),
    .C1(_03030_),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _19113_ (.A(\rbzero.spi_registers.texadd2[17] ),
    .B(_03023_),
    .X(_03032_));
 sky130_fd_sc_hd__o211a_1 _19114_ (.A1(\rbzero.spi_registers.new_texadd2[17] ),
    .A2(_03022_),
    .B1(_03032_),
    .C1(_03030_),
    .X(_00785_));
 sky130_fd_sc_hd__or2_1 _19115_ (.A(\rbzero.spi_registers.texadd2[18] ),
    .B(_03023_),
    .X(_03033_));
 sky130_fd_sc_hd__o211a_1 _19116_ (.A1(\rbzero.spi_registers.new_texadd2[18] ),
    .A2(_03022_),
    .B1(_03033_),
    .C1(_03030_),
    .X(_00786_));
 sky130_fd_sc_hd__or2_1 _19117_ (.A(\rbzero.spi_registers.texadd2[19] ),
    .B(_03023_),
    .X(_03034_));
 sky130_fd_sc_hd__o211a_1 _19118_ (.A1(\rbzero.spi_registers.new_texadd2[19] ),
    .A2(_03022_),
    .B1(_03034_),
    .C1(_03030_),
    .X(_00787_));
 sky130_fd_sc_hd__or2_1 _19119_ (.A(\rbzero.spi_registers.texadd2[20] ),
    .B(_03009_),
    .X(_03035_));
 sky130_fd_sc_hd__o211a_1 _19120_ (.A1(\rbzero.spi_registers.new_texadd2[20] ),
    .A2(_03007_),
    .B1(_03035_),
    .C1(_03030_),
    .X(_00788_));
 sky130_fd_sc_hd__or2_1 _19121_ (.A(\rbzero.spi_registers.texadd2[21] ),
    .B(_03009_),
    .X(_03036_));
 sky130_fd_sc_hd__o211a_1 _19122_ (.A1(\rbzero.spi_registers.new_texadd2[21] ),
    .A2(_03007_),
    .B1(_03036_),
    .C1(_03030_),
    .X(_00789_));
 sky130_fd_sc_hd__or2_1 _19123_ (.A(\rbzero.spi_registers.texadd2[22] ),
    .B(_03009_),
    .X(_03037_));
 sky130_fd_sc_hd__o211a_1 _19124_ (.A1(\rbzero.spi_registers.new_texadd2[22] ),
    .A2(_03007_),
    .B1(_03037_),
    .C1(_03030_),
    .X(_00790_));
 sky130_fd_sc_hd__or2_1 _19125_ (.A(\rbzero.spi_registers.texadd2[23] ),
    .B(_03009_),
    .X(_03038_));
 sky130_fd_sc_hd__o211a_1 _19126_ (.A1(\rbzero.spi_registers.new_texadd2[23] ),
    .A2(_03007_),
    .B1(_03038_),
    .C1(_03030_),
    .X(_00791_));
 sky130_fd_sc_hd__nand2_4 _19127_ (.A(\rbzero.spi_registers.got_new_texadd3 ),
    .B(_02860_),
    .Y(_03039_));
 sky130_fd_sc_hd__clkbuf_4 _19128_ (.A(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__and2_2 _19129_ (.A(\rbzero.spi_registers.got_new_texadd3 ),
    .B(_02864_),
    .X(_03041_));
 sky130_fd_sc_hd__buf_2 _19130_ (.A(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__or2_1 _19131_ (.A(\rbzero.spi_registers.texadd3[0] ),
    .B(_03042_),
    .X(_03043_));
 sky130_fd_sc_hd__o211a_1 _19132_ (.A1(\rbzero.spi_registers.new_texadd3[0] ),
    .A2(_03040_),
    .B1(_03043_),
    .C1(_03030_),
    .X(_00792_));
 sky130_fd_sc_hd__or2_1 _19133_ (.A(\rbzero.spi_registers.texadd3[1] ),
    .B(_03042_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_4 _19134_ (.A(_02973_),
    .X(_03045_));
 sky130_fd_sc_hd__o211a_1 _19135_ (.A1(\rbzero.spi_registers.new_texadd3[1] ),
    .A2(_03040_),
    .B1(_03044_),
    .C1(_03045_),
    .X(_00793_));
 sky130_fd_sc_hd__or2_1 _19136_ (.A(\rbzero.spi_registers.texadd3[2] ),
    .B(_03042_),
    .X(_03046_));
 sky130_fd_sc_hd__o211a_1 _19137_ (.A1(\rbzero.spi_registers.new_texadd3[2] ),
    .A2(_03040_),
    .B1(_03046_),
    .C1(_03045_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _19138_ (.A(\rbzero.spi_registers.texadd3[3] ),
    .B(_03042_),
    .X(_03047_));
 sky130_fd_sc_hd__o211a_1 _19139_ (.A1(\rbzero.spi_registers.new_texadd3[3] ),
    .A2(_03040_),
    .B1(_03047_),
    .C1(_03045_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _19140_ (.A(\rbzero.spi_registers.texadd3[4] ),
    .B(_03042_),
    .X(_03048_));
 sky130_fd_sc_hd__o211a_1 _19141_ (.A1(\rbzero.spi_registers.new_texadd3[4] ),
    .A2(_03040_),
    .B1(_03048_),
    .C1(_03045_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _19142_ (.A(\rbzero.spi_registers.texadd3[5] ),
    .B(_03042_),
    .X(_03049_));
 sky130_fd_sc_hd__o211a_1 _19143_ (.A1(\rbzero.spi_registers.new_texadd3[5] ),
    .A2(_03040_),
    .B1(_03049_),
    .C1(_03045_),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _19144_ (.A(\rbzero.spi_registers.texadd3[6] ),
    .B(_03042_),
    .X(_03050_));
 sky130_fd_sc_hd__o211a_1 _19145_ (.A1(\rbzero.spi_registers.new_texadd3[6] ),
    .A2(_03040_),
    .B1(_03050_),
    .C1(_03045_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _19146_ (.A(\rbzero.spi_registers.texadd3[7] ),
    .B(_03042_),
    .X(_03051_));
 sky130_fd_sc_hd__o211a_1 _19147_ (.A1(\rbzero.spi_registers.new_texadd3[7] ),
    .A2(_03040_),
    .B1(_03051_),
    .C1(_03045_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _19148_ (.A(\rbzero.spi_registers.texadd3[8] ),
    .B(_03042_),
    .X(_03052_));
 sky130_fd_sc_hd__o211a_1 _19149_ (.A1(\rbzero.spi_registers.new_texadd3[8] ),
    .A2(_03040_),
    .B1(_03052_),
    .C1(_03045_),
    .X(_00800_));
 sky130_fd_sc_hd__or2_1 _19150_ (.A(\rbzero.spi_registers.texadd3[9] ),
    .B(_03042_),
    .X(_03053_));
 sky130_fd_sc_hd__o211a_1 _19151_ (.A1(\rbzero.spi_registers.new_texadd3[9] ),
    .A2(_03040_),
    .B1(_03053_),
    .C1(_03045_),
    .X(_00801_));
 sky130_fd_sc_hd__clkbuf_4 _19152_ (.A(_03039_),
    .X(_03054_));
 sky130_fd_sc_hd__buf_2 _19153_ (.A(_03041_),
    .X(_03055_));
 sky130_fd_sc_hd__or2_1 _19154_ (.A(\rbzero.spi_registers.texadd3[10] ),
    .B(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__o211a_1 _19155_ (.A1(\rbzero.spi_registers.new_texadd3[10] ),
    .A2(_03054_),
    .B1(_03056_),
    .C1(_03045_),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _19156_ (.A(\rbzero.spi_registers.texadd3[11] ),
    .B(_03055_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_4 _19157_ (.A(_02973_),
    .X(_03058_));
 sky130_fd_sc_hd__o211a_1 _19158_ (.A1(\rbzero.spi_registers.new_texadd3[11] ),
    .A2(_03054_),
    .B1(_03057_),
    .C1(_03058_),
    .X(_00803_));
 sky130_fd_sc_hd__or2_1 _19159_ (.A(\rbzero.spi_registers.texadd3[12] ),
    .B(_03055_),
    .X(_03059_));
 sky130_fd_sc_hd__o211a_1 _19160_ (.A1(\rbzero.spi_registers.new_texadd3[12] ),
    .A2(_03054_),
    .B1(_03059_),
    .C1(_03058_),
    .X(_00804_));
 sky130_fd_sc_hd__or2_1 _19161_ (.A(\rbzero.spi_registers.texadd3[13] ),
    .B(_03055_),
    .X(_03060_));
 sky130_fd_sc_hd__o211a_1 _19162_ (.A1(\rbzero.spi_registers.new_texadd3[13] ),
    .A2(_03054_),
    .B1(_03060_),
    .C1(_03058_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _19163_ (.A(\rbzero.spi_registers.texadd3[14] ),
    .B(_03055_),
    .X(_03061_));
 sky130_fd_sc_hd__o211a_1 _19164_ (.A1(\rbzero.spi_registers.new_texadd3[14] ),
    .A2(_03054_),
    .B1(_03061_),
    .C1(_03058_),
    .X(_00806_));
 sky130_fd_sc_hd__or2_1 _19165_ (.A(\rbzero.spi_registers.texadd3[15] ),
    .B(_03055_),
    .X(_03062_));
 sky130_fd_sc_hd__o211a_1 _19166_ (.A1(\rbzero.spi_registers.new_texadd3[15] ),
    .A2(_03054_),
    .B1(_03062_),
    .C1(_03058_),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _19167_ (.A(\rbzero.spi_registers.texadd3[16] ),
    .B(_03055_),
    .X(_03063_));
 sky130_fd_sc_hd__o211a_1 _19168_ (.A1(\rbzero.spi_registers.new_texadd3[16] ),
    .A2(_03054_),
    .B1(_03063_),
    .C1(_03058_),
    .X(_00808_));
 sky130_fd_sc_hd__or2_1 _19169_ (.A(\rbzero.spi_registers.texadd3[17] ),
    .B(_03055_),
    .X(_03064_));
 sky130_fd_sc_hd__o211a_1 _19170_ (.A1(\rbzero.spi_registers.new_texadd3[17] ),
    .A2(_03054_),
    .B1(_03064_),
    .C1(_03058_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _19171_ (.A(\rbzero.spi_registers.texadd3[18] ),
    .B(_03055_),
    .X(_03065_));
 sky130_fd_sc_hd__o211a_1 _19172_ (.A1(\rbzero.spi_registers.new_texadd3[18] ),
    .A2(_03054_),
    .B1(_03065_),
    .C1(_03058_),
    .X(_00810_));
 sky130_fd_sc_hd__or2_1 _19173_ (.A(\rbzero.spi_registers.texadd3[19] ),
    .B(_03055_),
    .X(_03066_));
 sky130_fd_sc_hd__o211a_1 _19174_ (.A1(\rbzero.spi_registers.new_texadd3[19] ),
    .A2(_03054_),
    .B1(_03066_),
    .C1(_03058_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _19175_ (.A(\rbzero.spi_registers.texadd3[20] ),
    .B(_03041_),
    .X(_03067_));
 sky130_fd_sc_hd__o211a_1 _19176_ (.A1(\rbzero.spi_registers.new_texadd3[20] ),
    .A2(_03039_),
    .B1(_03067_),
    .C1(_03058_),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _19177_ (.A(\rbzero.spi_registers.texadd3[21] ),
    .B(_03041_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_4 _19178_ (.A(_02973_),
    .X(_03069_));
 sky130_fd_sc_hd__o211a_1 _19179_ (.A1(\rbzero.spi_registers.new_texadd3[21] ),
    .A2(_03039_),
    .B1(_03068_),
    .C1(_03069_),
    .X(_00813_));
 sky130_fd_sc_hd__or2_1 _19180_ (.A(\rbzero.spi_registers.texadd3[22] ),
    .B(_03041_),
    .X(_03070_));
 sky130_fd_sc_hd__o211a_1 _19181_ (.A1(\rbzero.spi_registers.new_texadd3[22] ),
    .A2(_03039_),
    .B1(_03070_),
    .C1(_03069_),
    .X(_00814_));
 sky130_fd_sc_hd__or2_1 _19182_ (.A(\rbzero.spi_registers.texadd3[23] ),
    .B(_03041_),
    .X(_03071_));
 sky130_fd_sc_hd__o211a_1 _19183_ (.A1(\rbzero.spi_registers.new_texadd3[23] ),
    .A2(_03039_),
    .B1(_03071_),
    .C1(_03069_),
    .X(_00815_));
 sky130_fd_sc_hd__clkinv_2 _19184_ (.A(_02792_),
    .Y(_03072_));
 sky130_fd_sc_hd__and4b_1 _19185_ (.A_N(\rbzero.spi_registers.spi_done ),
    .B(_02794_),
    .C(_02771_),
    .D(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _19186_ (.A(_03073_),
    .X(_00816_));
 sky130_fd_sc_hd__or3b_1 _19187_ (.A(_02487_),
    .B(_02488_),
    .C_N(\rbzero.spi_registers.spi_done ),
    .X(_03074_));
 sky130_fd_sc_hd__or3_1 _19188_ (.A(_04187_),
    .B(_02774_),
    .C(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_4 _19189_ (.A(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _19190_ (.A0(_02484_),
    .A1(\rbzero.spi_registers.new_sky[0] ),
    .S(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_1 _19191_ (.A(_03077_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _19192_ (.A0(_02494_),
    .A1(\rbzero.spi_registers.new_sky[1] ),
    .S(_03076_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _19193_ (.A(_03078_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _19194_ (.A0(_02496_),
    .A1(\rbzero.spi_registers.new_sky[2] ),
    .S(_03076_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _19195_ (.A(_03079_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _19196_ (.A0(_02498_),
    .A1(\rbzero.spi_registers.new_sky[3] ),
    .S(_03076_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _19197_ (.A(_03080_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _19198_ (.A0(_02500_),
    .A1(\rbzero.spi_registers.new_sky[4] ),
    .S(_03076_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _19199_ (.A(_03081_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _19200_ (.A0(_02502_),
    .A1(\rbzero.spi_registers.new_sky[5] ),
    .S(_03076_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _19201_ (.A(_03082_),
    .X(_00822_));
 sky130_fd_sc_hd__clkbuf_4 _19202_ (.A(_02881_),
    .X(_03083_));
 sky130_fd_sc_hd__inv_2 _19203_ (.A(_03076_),
    .Y(_03084_));
 sky130_fd_sc_hd__a31o_1 _19204_ (.A1(\rbzero.spi_registers.got_new_sky ),
    .A2(_02883_),
    .A3(_03083_),
    .B1(_03084_),
    .X(_00823_));
 sky130_fd_sc_hd__or4b_4 _19205_ (.A(_02485_),
    .B(_02486_),
    .C(_04187_),
    .D_N(\rbzero.spi_registers.spi_done ),
    .X(_03085_));
 sky130_fd_sc_hd__nor3_4 _19206_ (.A(_02487_),
    .B(_02488_),
    .C(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__mux2_1 _19207_ (.A0(\rbzero.spi_registers.new_floor[0] ),
    .A1(_02484_),
    .S(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _19208_ (.A(_03087_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _19209_ (.A0(\rbzero.spi_registers.new_floor[1] ),
    .A1(_02494_),
    .S(_03086_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_1 _19210_ (.A(_03088_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _19211_ (.A0(\rbzero.spi_registers.new_floor[2] ),
    .A1(_02496_),
    .S(_03086_),
    .X(_03089_));
 sky130_fd_sc_hd__clkbuf_1 _19212_ (.A(_03089_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _19213_ (.A0(\rbzero.spi_registers.new_floor[3] ),
    .A1(_02498_),
    .S(_03086_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _19214_ (.A(_03090_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _19215_ (.A0(\rbzero.spi_registers.new_floor[4] ),
    .A1(_02500_),
    .S(_03086_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _19216_ (.A(_03091_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _19217_ (.A0(\rbzero.spi_registers.new_floor[5] ),
    .A1(_02502_),
    .S(_03086_),
    .X(_03092_));
 sky130_fd_sc_hd__clkbuf_1 _19218_ (.A(_03092_),
    .X(_00829_));
 sky130_fd_sc_hd__a31o_1 _19219_ (.A1(\rbzero.spi_registers.got_new_floor ),
    .A2(_02883_),
    .A3(_03083_),
    .B1(_03086_),
    .X(_00830_));
 sky130_fd_sc_hd__or4b_2 _19220_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_04187_),
    .C(_03074_),
    .D_N(_02485_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_4 _19221_ (.A(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__mux2_1 _19222_ (.A0(_02484_),
    .A1(\rbzero.spi_registers.new_leak[0] ),
    .S(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_1 _19223_ (.A(_03095_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _19224_ (.A0(_02494_),
    .A1(\rbzero.spi_registers.new_leak[1] ),
    .S(_03094_),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _19225_ (.A(_03096_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _19226_ (.A0(_02496_),
    .A1(\rbzero.spi_registers.new_leak[2] ),
    .S(_03094_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _19227_ (.A(_03097_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _19228_ (.A0(_02498_),
    .A1(\rbzero.spi_registers.new_leak[3] ),
    .S(_03094_),
    .X(_03098_));
 sky130_fd_sc_hd__clkbuf_1 _19229_ (.A(_03098_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _19230_ (.A0(_02500_),
    .A1(\rbzero.spi_registers.new_leak[4] ),
    .S(_03094_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _19231_ (.A(_03099_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _19232_ (.A0(_02502_),
    .A1(\rbzero.spi_registers.new_leak[5] ),
    .S(_03094_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _19233_ (.A(_03100_),
    .X(_00836_));
 sky130_fd_sc_hd__inv_2 _19234_ (.A(_03094_),
    .Y(_03101_));
 sky130_fd_sc_hd__a31o_1 _19235_ (.A1(\rbzero.spi_registers.got_new_leak ),
    .A2(_02883_),
    .A3(_03083_),
    .B1(_03101_),
    .X(_00837_));
 sky130_fd_sc_hd__or3_1 _19236_ (.A(_04187_),
    .B(_02776_),
    .C(_03074_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_4 _19237_ (.A(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _19238_ (.A0(_02484_),
    .A1(\rbzero.spi_registers.new_other[0] ),
    .S(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _19239_ (.A(_03104_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _19240_ (.A0(_02494_),
    .A1(\rbzero.spi_registers.new_other[1] ),
    .S(_03103_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _19241_ (.A(_03105_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _19242_ (.A0(_02496_),
    .A1(\rbzero.spi_registers.new_other[2] ),
    .S(_03103_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _19243_ (.A(_03106_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _19244_ (.A0(_02498_),
    .A1(\rbzero.spi_registers.new_other[3] ),
    .S(_03103_),
    .X(_03107_));
 sky130_fd_sc_hd__clkbuf_1 _19245_ (.A(_03107_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _19246_ (.A0(_02500_),
    .A1(\rbzero.spi_registers.new_other[4] ),
    .S(_03103_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _19247_ (.A(_03108_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _19248_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(\rbzero.spi_registers.new_other[6] ),
    .S(_03103_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _19249_ (.A(_03109_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _19250_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.new_other[7] ),
    .S(_03103_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _19251_ (.A(_03110_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _19252_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.new_other[8] ),
    .S(_03103_),
    .X(_03111_));
 sky130_fd_sc_hd__clkbuf_1 _19253_ (.A(_03111_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _19254_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.new_other[9] ),
    .S(_03103_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _19255_ (.A(_03112_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _19256_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.new_other[10] ),
    .S(_03102_),
    .X(_03113_));
 sky130_fd_sc_hd__clkbuf_1 _19257_ (.A(_03113_),
    .X(_00847_));
 sky130_fd_sc_hd__inv_2 _19258_ (.A(_03103_),
    .Y(_03114_));
 sky130_fd_sc_hd__a31o_1 _19259_ (.A1(\rbzero.spi_registers.got_new_other ),
    .A2(_02883_),
    .A3(_03083_),
    .B1(_03114_),
    .X(_00848_));
 sky130_fd_sc_hd__nor2_1 _19260_ (.A(_02485_),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .Y(_03115_));
 sky130_fd_sc_hd__and4_1 _19261_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_08244_),
    .C(_02773_),
    .D(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_2 _19262_ (.A(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _19263_ (.A0(\rbzero.spi_registers.new_vshift[0] ),
    .A1(_02484_),
    .S(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _19264_ (.A(_03118_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _19265_ (.A0(\rbzero.spi_registers.new_vshift[1] ),
    .A1(_02494_),
    .S(_03117_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _19266_ (.A(_03119_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _19267_ (.A0(\rbzero.spi_registers.new_vshift[2] ),
    .A1(_02496_),
    .S(_03117_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _19268_ (.A(_03120_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _19269_ (.A0(\rbzero.spi_registers.new_vshift[3] ),
    .A1(_02498_),
    .S(_03117_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_1 _19270_ (.A(_03121_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _19271_ (.A0(\rbzero.spi_registers.new_vshift[4] ),
    .A1(_02500_),
    .S(_03117_),
    .X(_03122_));
 sky130_fd_sc_hd__clkbuf_1 _19272_ (.A(_03122_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _19273_ (.A0(\rbzero.spi_registers.new_vshift[5] ),
    .A1(_02502_),
    .S(_03117_),
    .X(_03123_));
 sky130_fd_sc_hd__clkbuf_1 _19274_ (.A(_03123_),
    .X(_00854_));
 sky130_fd_sc_hd__a31o_1 _19275_ (.A1(\rbzero.spi_registers.got_new_vshift ),
    .A2(_08246_),
    .A3(_03083_),
    .B1(_03117_),
    .X(_00855_));
 sky130_fd_sc_hd__nor3b_1 _19276_ (.A(_02488_),
    .B(_03085_),
    .C_N(_02487_),
    .Y(_03124_));
 sky130_fd_sc_hd__mux2_1 _19277_ (.A0(\rbzero.spi_registers.new_vinf ),
    .A1(_02484_),
    .S(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__clkbuf_1 _19278_ (.A(_03125_),
    .X(_00856_));
 sky130_fd_sc_hd__a31o_1 _19279_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_08246_),
    .A3(_03083_),
    .B1(_03124_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_2 _19280_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_04108_),
    .Y(_03126_));
 sky130_fd_sc_hd__nor2_4 _19281_ (.A(_02779_),
    .B(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__clkbuf_4 _19282_ (.A(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_1 _19283_ (.A0(\rbzero.spi_registers.new_mapd[0] ),
    .A1(_02484_),
    .S(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _19284_ (.A(_03129_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _19285_ (.A0(\rbzero.spi_registers.new_mapd[1] ),
    .A1(_02494_),
    .S(_03128_),
    .X(_03130_));
 sky130_fd_sc_hd__clkbuf_1 _19286_ (.A(_03130_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _19287_ (.A0(\rbzero.spi_registers.new_mapd[2] ),
    .A1(_02496_),
    .S(_03128_),
    .X(_03131_));
 sky130_fd_sc_hd__clkbuf_1 _19288_ (.A(_03131_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _19289_ (.A0(\rbzero.spi_registers.new_mapd[3] ),
    .A1(_02498_),
    .S(_03128_),
    .X(_03132_));
 sky130_fd_sc_hd__clkbuf_1 _19290_ (.A(_03132_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _19291_ (.A0(\rbzero.spi_registers.new_mapd[4] ),
    .A1(_02500_),
    .S(_03128_),
    .X(_03133_));
 sky130_fd_sc_hd__clkbuf_1 _19292_ (.A(_03133_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _19293_ (.A0(\rbzero.spi_registers.new_mapd[5] ),
    .A1(_02502_),
    .S(_03128_),
    .X(_03134_));
 sky130_fd_sc_hd__clkbuf_1 _19294_ (.A(_03134_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _19295_ (.A0(\rbzero.spi_registers.new_mapd[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03128_),
    .X(_03135_));
 sky130_fd_sc_hd__clkbuf_1 _19296_ (.A(_03135_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _19297_ (.A0(\rbzero.spi_registers.new_mapd[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03128_),
    .X(_03136_));
 sky130_fd_sc_hd__clkbuf_1 _19298_ (.A(_03136_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _19299_ (.A0(\rbzero.spi_registers.new_mapd[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03128_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_1 _19300_ (.A(_03137_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _19301_ (.A0(\rbzero.spi_registers.new_mapd[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03127_),
    .X(_03138_));
 sky130_fd_sc_hd__clkbuf_1 _19302_ (.A(_03138_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _19303_ (.A0(\rbzero.spi_registers.new_mapd[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03127_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_1 _19304_ (.A(_03139_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _19305_ (.A0(\rbzero.spi_registers.new_mapd[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03127_),
    .X(_03140_));
 sky130_fd_sc_hd__clkbuf_1 _19306_ (.A(_03140_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _19307_ (.A0(\rbzero.spi_registers.new_mapd[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03127_),
    .X(_03141_));
 sky130_fd_sc_hd__clkbuf_1 _19308_ (.A(_03141_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _19309_ (.A0(\rbzero.spi_registers.new_mapd[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03127_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_1 _19310_ (.A(_03142_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _19311_ (.A0(\rbzero.spi_registers.new_mapd[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03127_),
    .X(_03143_));
 sky130_fd_sc_hd__clkbuf_1 _19312_ (.A(_03143_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _19313_ (.A0(\rbzero.spi_registers.new_mapd[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03127_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_1 _19314_ (.A(_03144_),
    .X(_00873_));
 sky130_fd_sc_hd__a31o_1 _19315_ (.A1(\rbzero.spi_registers.got_new_mapd ),
    .A2(_08246_),
    .A3(_03083_),
    .B1(_03128_),
    .X(_00874_));
 sky130_fd_sc_hd__nor4b_4 _19316_ (.A(_02488_),
    .B(_02776_),
    .C(_03126_),
    .D_N(_02487_),
    .Y(_03145_));
 sky130_fd_sc_hd__buf_4 _19317_ (.A(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_1 _19318_ (.A0(\rbzero.spi_registers.new_texadd0[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_1 _19319_ (.A(_03147_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _19320_ (.A0(\rbzero.spi_registers.new_texadd0[1] ),
    .A1(_02494_),
    .S(_03146_),
    .X(_03148_));
 sky130_fd_sc_hd__clkbuf_1 _19321_ (.A(_03148_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _19322_ (.A0(\rbzero.spi_registers.new_texadd0[2] ),
    .A1(_02496_),
    .S(_03146_),
    .X(_03149_));
 sky130_fd_sc_hd__clkbuf_1 _19323_ (.A(_03149_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _19324_ (.A0(\rbzero.spi_registers.new_texadd0[3] ),
    .A1(_02498_),
    .S(_03146_),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_1 _19325_ (.A(_03150_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _19326_ (.A0(\rbzero.spi_registers.new_texadd0[4] ),
    .A1(_02500_),
    .S(_03146_),
    .X(_03151_));
 sky130_fd_sc_hd__clkbuf_1 _19327_ (.A(_03151_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _19328_ (.A0(\rbzero.spi_registers.new_texadd0[5] ),
    .A1(_02502_),
    .S(_03146_),
    .X(_03152_));
 sky130_fd_sc_hd__clkbuf_1 _19329_ (.A(_03152_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _19330_ (.A0(\rbzero.spi_registers.new_texadd0[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03146_),
    .X(_03153_));
 sky130_fd_sc_hd__clkbuf_1 _19331_ (.A(_03153_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _19332_ (.A0(\rbzero.spi_registers.new_texadd0[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03146_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_1 _19333_ (.A(_03154_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _19334_ (.A0(\rbzero.spi_registers.new_texadd0[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03146_),
    .X(_03155_));
 sky130_fd_sc_hd__clkbuf_1 _19335_ (.A(_03155_),
    .X(_00883_));
 sky130_fd_sc_hd__buf_4 _19336_ (.A(_03145_),
    .X(_03156_));
 sky130_fd_sc_hd__mux2_1 _19337_ (.A0(\rbzero.spi_registers.new_texadd0[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_1 _19338_ (.A(_03157_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _19339_ (.A0(\rbzero.spi_registers.new_texadd0[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03156_),
    .X(_03158_));
 sky130_fd_sc_hd__clkbuf_1 _19340_ (.A(_03158_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _19341_ (.A0(\rbzero.spi_registers.new_texadd0[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03156_),
    .X(_03159_));
 sky130_fd_sc_hd__clkbuf_1 _19342_ (.A(_03159_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _19343_ (.A0(\rbzero.spi_registers.new_texadd0[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03156_),
    .X(_03160_));
 sky130_fd_sc_hd__clkbuf_1 _19344_ (.A(_03160_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _19345_ (.A0(\rbzero.spi_registers.new_texadd0[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03156_),
    .X(_03161_));
 sky130_fd_sc_hd__clkbuf_1 _19346_ (.A(_03161_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _19347_ (.A0(\rbzero.spi_registers.new_texadd0[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03156_),
    .X(_03162_));
 sky130_fd_sc_hd__clkbuf_1 _19348_ (.A(_03162_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _19349_ (.A0(\rbzero.spi_registers.new_texadd0[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03156_),
    .X(_03163_));
 sky130_fd_sc_hd__clkbuf_1 _19350_ (.A(_03163_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _19351_ (.A0(\rbzero.spi_registers.new_texadd0[16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03156_),
    .X(_03164_));
 sky130_fd_sc_hd__clkbuf_1 _19352_ (.A(_03164_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _19353_ (.A0(\rbzero.spi_registers.new_texadd0[17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03156_),
    .X(_03165_));
 sky130_fd_sc_hd__clkbuf_1 _19354_ (.A(_03165_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _19355_ (.A0(\rbzero.spi_registers.new_texadd0[18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03156_),
    .X(_03166_));
 sky130_fd_sc_hd__clkbuf_1 _19356_ (.A(_03166_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _19357_ (.A0(\rbzero.spi_registers.new_texadd0[19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03145_),
    .X(_03167_));
 sky130_fd_sc_hd__clkbuf_1 _19358_ (.A(_03167_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _19359_ (.A0(\rbzero.spi_registers.new_texadd0[20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03145_),
    .X(_03168_));
 sky130_fd_sc_hd__clkbuf_1 _19360_ (.A(_03168_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _19361_ (.A0(\rbzero.spi_registers.new_texadd0[21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03145_),
    .X(_03169_));
 sky130_fd_sc_hd__clkbuf_1 _19362_ (.A(_03169_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _19363_ (.A0(\rbzero.spi_registers.new_texadd0[22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03145_),
    .X(_03170_));
 sky130_fd_sc_hd__clkbuf_1 _19364_ (.A(_03170_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _19365_ (.A0(\rbzero.spi_registers.new_texadd0[23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03145_),
    .X(_03171_));
 sky130_fd_sc_hd__clkbuf_1 _19366_ (.A(_03171_),
    .X(_00898_));
 sky130_fd_sc_hd__a31o_1 _19367_ (.A1(\rbzero.spi_registers.got_new_texadd0 ),
    .A2(_08246_),
    .A3(_03083_),
    .B1(_03146_),
    .X(_00899_));
 sky130_fd_sc_hd__and3_1 _19368_ (.A(_04108_),
    .B(_02489_),
    .C(_03115_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_4 _19369_ (.A(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__buf_4 _19370_ (.A(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _19371_ (.A0(\rbzero.spi_registers.new_texadd1[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_1 _19372_ (.A(_03175_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _19373_ (.A0(\rbzero.spi_registers.new_texadd1[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_03174_),
    .X(_03176_));
 sky130_fd_sc_hd__clkbuf_1 _19374_ (.A(_03176_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _19375_ (.A0(\rbzero.spi_registers.new_texadd1[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_03174_),
    .X(_03177_));
 sky130_fd_sc_hd__clkbuf_1 _19376_ (.A(_03177_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _19377_ (.A0(\rbzero.spi_registers.new_texadd1[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_03174_),
    .X(_03178_));
 sky130_fd_sc_hd__clkbuf_1 _19378_ (.A(_03178_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _19379_ (.A0(\rbzero.spi_registers.new_texadd1[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_03174_),
    .X(_03179_));
 sky130_fd_sc_hd__clkbuf_1 _19380_ (.A(_03179_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _19381_ (.A0(\rbzero.spi_registers.new_texadd1[5] ),
    .A1(_02502_),
    .S(_03174_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_1 _19382_ (.A(_03180_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _19383_ (.A0(\rbzero.spi_registers.new_texadd1[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03174_),
    .X(_03181_));
 sky130_fd_sc_hd__clkbuf_1 _19384_ (.A(_03181_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _19385_ (.A0(\rbzero.spi_registers.new_texadd1[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03174_),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_1 _19386_ (.A(_03182_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _19387_ (.A0(\rbzero.spi_registers.new_texadd1[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03174_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_1 _19388_ (.A(_03183_),
    .X(_00908_));
 sky130_fd_sc_hd__buf_4 _19389_ (.A(_03173_),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_1 _19390_ (.A0(\rbzero.spi_registers.new_texadd1[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_1 _19391_ (.A(_03185_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _19392_ (.A0(\rbzero.spi_registers.new_texadd1[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03184_),
    .X(_03186_));
 sky130_fd_sc_hd__clkbuf_1 _19393_ (.A(_03186_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _19394_ (.A0(\rbzero.spi_registers.new_texadd1[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03184_),
    .X(_03187_));
 sky130_fd_sc_hd__clkbuf_1 _19395_ (.A(_03187_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _19396_ (.A0(\rbzero.spi_registers.new_texadd1[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03184_),
    .X(_03188_));
 sky130_fd_sc_hd__clkbuf_1 _19397_ (.A(_03188_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _19398_ (.A0(\rbzero.spi_registers.new_texadd1[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03184_),
    .X(_03189_));
 sky130_fd_sc_hd__clkbuf_1 _19399_ (.A(_03189_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _19400_ (.A0(\rbzero.spi_registers.new_texadd1[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03184_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_1 _19401_ (.A(_03190_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _19402_ (.A0(\rbzero.spi_registers.new_texadd1[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03184_),
    .X(_03191_));
 sky130_fd_sc_hd__clkbuf_1 _19403_ (.A(_03191_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _19404_ (.A0(\rbzero.spi_registers.new_texadd1[16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03184_),
    .X(_03192_));
 sky130_fd_sc_hd__clkbuf_1 _19405_ (.A(_03192_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _19406_ (.A0(\rbzero.spi_registers.new_texadd1[17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03184_),
    .X(_03193_));
 sky130_fd_sc_hd__clkbuf_1 _19407_ (.A(_03193_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _19408_ (.A0(\rbzero.spi_registers.new_texadd1[18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03184_),
    .X(_03194_));
 sky130_fd_sc_hd__clkbuf_1 _19409_ (.A(_03194_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _19410_ (.A0(\rbzero.spi_registers.new_texadd1[19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03173_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _19411_ (.A(_03195_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _19412_ (.A0(\rbzero.spi_registers.new_texadd1[20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03173_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _19413_ (.A(_03196_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _19414_ (.A0(\rbzero.spi_registers.new_texadd1[21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03173_),
    .X(_03197_));
 sky130_fd_sc_hd__clkbuf_1 _19415_ (.A(_03197_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _19416_ (.A0(\rbzero.spi_registers.new_texadd1[22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03173_),
    .X(_03198_));
 sky130_fd_sc_hd__clkbuf_1 _19417_ (.A(_03198_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _19418_ (.A0(\rbzero.spi_registers.new_texadd1[23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03173_),
    .X(_03199_));
 sky130_fd_sc_hd__clkbuf_1 _19419_ (.A(_03199_),
    .X(_00923_));
 sky130_fd_sc_hd__a31o_1 _19420_ (.A1(\rbzero.spi_registers.got_new_texadd1 ),
    .A2(_08246_),
    .A3(_03083_),
    .B1(_03174_),
    .X(_00924_));
 sky130_fd_sc_hd__nor3b_4 _19421_ (.A(_03085_),
    .B(_02487_),
    .C_N(_02488_),
    .Y(_03200_));
 sky130_fd_sc_hd__buf_4 _19422_ (.A(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _19423_ (.A0(\rbzero.spi_registers.new_texadd2[0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__clkbuf_1 _19424_ (.A(_03202_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _19425_ (.A0(\rbzero.spi_registers.new_texadd2[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_03201_),
    .X(_03203_));
 sky130_fd_sc_hd__clkbuf_1 _19426_ (.A(_03203_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _19427_ (.A0(\rbzero.spi_registers.new_texadd2[2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_03201_),
    .X(_03204_));
 sky130_fd_sc_hd__clkbuf_1 _19428_ (.A(_03204_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19429_ (.A0(\rbzero.spi_registers.new_texadd2[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_03201_),
    .X(_03205_));
 sky130_fd_sc_hd__clkbuf_1 _19430_ (.A(_03205_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _19431_ (.A0(\rbzero.spi_registers.new_texadd2[4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_03201_),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_1 _19432_ (.A(_03206_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19433_ (.A0(\rbzero.spi_registers.new_texadd2[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_03201_),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_1 _19434_ (.A(_03207_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _19435_ (.A0(\rbzero.spi_registers.new_texadd2[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03201_),
    .X(_03208_));
 sky130_fd_sc_hd__clkbuf_1 _19436_ (.A(_03208_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _19437_ (.A0(\rbzero.spi_registers.new_texadd2[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03201_),
    .X(_03209_));
 sky130_fd_sc_hd__clkbuf_1 _19438_ (.A(_03209_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _19439_ (.A0(\rbzero.spi_registers.new_texadd2[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03201_),
    .X(_03210_));
 sky130_fd_sc_hd__clkbuf_1 _19440_ (.A(_03210_),
    .X(_00933_));
 sky130_fd_sc_hd__buf_4 _19441_ (.A(_03200_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _19442_ (.A0(\rbzero.spi_registers.new_texadd2[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_1 _19443_ (.A(_03212_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _19444_ (.A0(\rbzero.spi_registers.new_texadd2[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03211_),
    .X(_03213_));
 sky130_fd_sc_hd__clkbuf_1 _19445_ (.A(_03213_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _19446_ (.A0(\rbzero.spi_registers.new_texadd2[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03211_),
    .X(_03214_));
 sky130_fd_sc_hd__clkbuf_1 _19447_ (.A(_03214_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _19448_ (.A0(\rbzero.spi_registers.new_texadd2[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03211_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_1 _19449_ (.A(_03215_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _19450_ (.A0(\rbzero.spi_registers.new_texadd2[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03211_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_1 _19451_ (.A(_03216_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _19452_ (.A0(\rbzero.spi_registers.new_texadd2[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03211_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_1 _19453_ (.A(_03217_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _19454_ (.A0(\rbzero.spi_registers.new_texadd2[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03211_),
    .X(_03218_));
 sky130_fd_sc_hd__clkbuf_1 _19455_ (.A(_03218_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _19456_ (.A0(\rbzero.spi_registers.new_texadd2[16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03211_),
    .X(_03219_));
 sky130_fd_sc_hd__clkbuf_1 _19457_ (.A(_03219_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _19458_ (.A0(\rbzero.spi_registers.new_texadd2[17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03211_),
    .X(_03220_));
 sky130_fd_sc_hd__clkbuf_1 _19459_ (.A(_03220_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _19460_ (.A0(\rbzero.spi_registers.new_texadd2[18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03211_),
    .X(_03221_));
 sky130_fd_sc_hd__clkbuf_1 _19461_ (.A(_03221_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _19462_ (.A0(\rbzero.spi_registers.new_texadd2[19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03200_),
    .X(_03222_));
 sky130_fd_sc_hd__clkbuf_1 _19463_ (.A(_03222_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _19464_ (.A0(\rbzero.spi_registers.new_texadd2[20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03200_),
    .X(_03223_));
 sky130_fd_sc_hd__clkbuf_1 _19465_ (.A(_03223_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _19466_ (.A0(\rbzero.spi_registers.new_texadd2[21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03200_),
    .X(_03224_));
 sky130_fd_sc_hd__clkbuf_1 _19467_ (.A(_03224_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _19468_ (.A0(\rbzero.spi_registers.new_texadd2[22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03200_),
    .X(_03225_));
 sky130_fd_sc_hd__clkbuf_1 _19469_ (.A(_03225_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _19470_ (.A0(\rbzero.spi_registers.new_texadd2[23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03200_),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_1 _19471_ (.A(_03226_),
    .X(_00948_));
 sky130_fd_sc_hd__a31o_1 _19472_ (.A1(\rbzero.spi_registers.got_new_texadd2 ),
    .A2(_08246_),
    .A3(_03083_),
    .B1(_03201_),
    .X(_00949_));
 sky130_fd_sc_hd__and2_1 _19473_ (.A(net54),
    .B(_02850_),
    .X(_03227_));
 sky130_fd_sc_hd__clkbuf_1 _19474_ (.A(_03227_),
    .X(_00950_));
 sky130_fd_sc_hd__and2_1 _19475_ (.A(\rbzero.pov.ss_buffer[0] ),
    .B(_02850_),
    .X(_03228_));
 sky130_fd_sc_hd__clkbuf_1 _19476_ (.A(_03228_),
    .X(_00951_));
 sky130_fd_sc_hd__nor2_1 _19477_ (.A(_05226_),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _19478_ (.A(_05226_),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_03230_));
 sky130_fd_sc_hd__and2b_1 _19479_ (.A_N(_03229_),
    .B(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_4 _19480_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_03232_));
 sky130_fd_sc_hd__nor2_1 _19481_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_03233_));
 sky130_fd_sc_hd__nand2_1 _19482_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .Y(_03234_));
 sky130_fd_sc_hd__nor2_1 _19483_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_03235_));
 sky130_fd_sc_hd__and2_1 _19484_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_03236_));
 sky130_fd_sc_hd__o21ba_1 _19485_ (.A1(_03234_),
    .A2(_03235_),
    .B1_N(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__nand2_1 _19486_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_03238_));
 sky130_fd_sc_hd__o21ai_1 _19487_ (.A1(_03233_),
    .A2(_03237_),
    .B1(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__a21o_1 _19488_ (.A1(_03232_),
    .A2(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B1(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__o21ai_1 _19489_ (.A1(_03232_),
    .A2(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B1(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__xnor2_1 _19490_ (.A(_03231_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__a22o_1 _19491_ (.A1(\rbzero.debug_overlay.vplaneY[-9] ),
    .A2(_02539_),
    .B1(_09886_),
    .B2(\rbzero.wall_tracer.rayAddendY[-5] ),
    .X(_03243_));
 sky130_fd_sc_hd__a21o_1 _19492_ (.A1(_09885_),
    .A2(_03242_),
    .B1(_03243_),
    .X(_00952_));
 sky130_fd_sc_hd__nor2_1 _19493_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .Y(_03244_));
 sky130_fd_sc_hd__and2_1 _19494_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_03245_));
 sky130_fd_sc_hd__o21ai_1 _19495_ (.A1(_03229_),
    .A2(_03241_),
    .B1(_03230_),
    .Y(_03246_));
 sky130_fd_sc_hd__or3_1 _19496_ (.A(_03244_),
    .B(_03245_),
    .C(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__o21ai_1 _19497_ (.A1(_03244_),
    .A2(_03245_),
    .B1(_03246_),
    .Y(_03248_));
 sky130_fd_sc_hd__a21oi_1 _19498_ (.A1(_03247_),
    .A2(_03248_),
    .B1(_08262_),
    .Y(_03249_));
 sky130_fd_sc_hd__nand2_1 _19499_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_03250_));
 sky130_fd_sc_hd__or2_1 _19500_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_03251_));
 sky130_fd_sc_hd__a31o_1 _19501_ (.A1(_02544_),
    .A2(_03250_),
    .A3(_03251_),
    .B1(_09881_),
    .X(_03252_));
 sky130_fd_sc_hd__o22a_1 _19502_ (.A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_02551_),
    .B1(_03249_),
    .B2(_03252_),
    .X(_00953_));
 sky130_fd_sc_hd__nor2_1 _19503_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_03253_));
 sky130_fd_sc_hd__and2_1 _19504_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .X(_03254_));
 sky130_fd_sc_hd__or2_1 _19505_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_03255_));
 sky130_fd_sc_hd__a21oi_1 _19506_ (.A1(_03255_),
    .A2(_03246_),
    .B1(_03245_),
    .Y(_03256_));
 sky130_fd_sc_hd__o21ai_1 _19507_ (.A1(_03253_),
    .A2(_03254_),
    .B1(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__o311a_1 _19508_ (.A1(_03253_),
    .A2(_03254_),
    .A3(_03256_),
    .B1(_03257_),
    .C1(_04576_),
    .X(_03258_));
 sky130_fd_sc_hd__or2_1 _19509_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03251_),
    .X(_03259_));
 sky130_fd_sc_hd__nand2_1 _19510_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03251_),
    .Y(_03260_));
 sky130_fd_sc_hd__a31o_1 _19511_ (.A1(_02544_),
    .A2(_03259_),
    .A3(_03260_),
    .B1(_09881_),
    .X(_03261_));
 sky130_fd_sc_hd__o22a_1 _19512_ (.A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A2(_02551_),
    .B1(_03258_),
    .B2(_03261_),
    .X(_00954_));
 sky130_fd_sc_hd__buf_2 _19513_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_03262_));
 sky130_fd_sc_hd__nor2_1 _19514_ (.A(_03262_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_03263_));
 sky130_fd_sc_hd__and2_1 _19515_ (.A(_03262_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_03264_));
 sky130_fd_sc_hd__nand2_1 _19516_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_03265_));
 sky130_fd_sc_hd__o21ai_1 _19517_ (.A1(_03253_),
    .A2(_03256_),
    .B1(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__or3_1 _19518_ (.A(_03263_),
    .B(_03264_),
    .C(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__o21ai_1 _19519_ (.A1(_03263_),
    .A2(_03264_),
    .B1(_03266_),
    .Y(_03268_));
 sky130_fd_sc_hd__a21oi_1 _19520_ (.A1(_03267_),
    .A2(_03268_),
    .B1(_08262_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand2_1 _19521_ (.A(_03232_),
    .B(_03259_),
    .Y(_03270_));
 sky130_fd_sc_hd__or2_1 _19522_ (.A(_03232_),
    .B(_03259_),
    .X(_03271_));
 sky130_fd_sc_hd__a31o_1 _19523_ (.A1(_02544_),
    .A2(_03270_),
    .A3(_03271_),
    .B1(_09880_),
    .X(_03272_));
 sky130_fd_sc_hd__o22a_1 _19524_ (.A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A2(_02551_),
    .B1(_03269_),
    .B2(_03272_),
    .X(_00955_));
 sky130_fd_sc_hd__or2_1 _19525_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_03273_));
 sky130_fd_sc_hd__nand2_1 _19526_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_03274_));
 sky130_fd_sc_hd__or2_1 _19527_ (.A(_03262_),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_03275_));
 sky130_fd_sc_hd__a21o_1 _19528_ (.A1(_03275_),
    .A2(_03266_),
    .B1(_03264_),
    .X(_03276_));
 sky130_fd_sc_hd__nand3_1 _19529_ (.A(_03273_),
    .B(_03274_),
    .C(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__a21o_1 _19530_ (.A1(_03273_),
    .A2(_03274_),
    .B1(_03276_),
    .X(_03278_));
 sky130_fd_sc_hd__inv_2 _19531_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_03279_));
 sky130_fd_sc_hd__o31a_1 _19532_ (.A1(_03232_),
    .A2(\rbzero.debug_overlay.vplaneY[-7] ),
    .A3(\rbzero.debug_overlay.vplaneY[-8] ),
    .B1(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__xor2_1 _19533_ (.A(_05226_),
    .B(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__a22o_1 _19534_ (.A1(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A2(_09880_),
    .B1(_03281_),
    .B2(_02539_),
    .X(_03282_));
 sky130_fd_sc_hd__a31o_1 _19535_ (.A1(_09888_),
    .A2(_03277_),
    .A3(_03278_),
    .B1(_03282_),
    .X(_00956_));
 sky130_fd_sc_hd__a21bo_1 _19536_ (.A1(_03273_),
    .A2(_03276_),
    .B1_N(_03274_),
    .X(_03283_));
 sky130_fd_sc_hd__clkbuf_4 _19537_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_03284_));
 sky130_fd_sc_hd__nor2_1 _19538_ (.A(_03284_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_03285_));
 sky130_fd_sc_hd__and2_1 _19539_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_03286_));
 sky130_fd_sc_hd__or2_1 _19540_ (.A(_03285_),
    .B(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__xnor2_1 _19541_ (.A(_03283_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__or2_1 _19542_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_03289_));
 sky130_fd_sc_hd__nand2_1 _19543_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_03290_));
 sky130_fd_sc_hd__nand2_1 _19544_ (.A(_03289_),
    .B(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__nor2_1 _19545_ (.A(_05226_),
    .B(_03271_),
    .Y(_03292_));
 sky130_fd_sc_hd__a21oi_1 _19546_ (.A1(_05226_),
    .A2(\rbzero.debug_overlay.vplaneY[-9] ),
    .B1(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__xnor2_1 _19547_ (.A(_03291_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__mux2_1 _19548_ (.A0(_03288_),
    .A1(_03294_),
    .S(_04566_),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _19549_ (.A0(\rbzero.wall_tracer.rayAddendY[0] ),
    .A1(_03295_),
    .S(_02550_),
    .X(_03296_));
 sky130_fd_sc_hd__clkbuf_1 _19550_ (.A(_03296_),
    .X(_00957_));
 sky130_fd_sc_hd__nand2_1 _19551_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_03297_));
 sky130_fd_sc_hd__or2_1 _19552_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_03298_));
 sky130_fd_sc_hd__o21a_1 _19553_ (.A1(_03284_),
    .A2(\rbzero.wall_tracer.rayAddendY[0] ),
    .B1(_03283_),
    .X(_03299_));
 sky130_fd_sc_hd__a211o_1 _19554_ (.A1(_03297_),
    .A2(_03298_),
    .B1(_03299_),
    .C1(_03286_),
    .X(_03300_));
 sky130_fd_sc_hd__o211ai_2 _19555_ (.A1(_03286_),
    .A2(_03299_),
    .B1(_03298_),
    .C1(_03297_),
    .Y(_03301_));
 sky130_fd_sc_hd__a21oi_1 _19556_ (.A1(_05226_),
    .A2(\rbzero.debug_overlay.vplaneY[-9] ),
    .B1(_03291_),
    .Y(_03302_));
 sky130_fd_sc_hd__nor2_1 _19557_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_03303_));
 sky130_fd_sc_hd__and2_1 _19558_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(_03304_));
 sky130_fd_sc_hd__nor2_1 _19559_ (.A(_03303_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__xnor2_1 _19560_ (.A(_03289_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__o21a_1 _19561_ (.A1(_03292_),
    .A2(_03302_),
    .B1(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__inv_2 _19562_ (.A(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__or3_1 _19563_ (.A(_03292_),
    .B(_03306_),
    .C(_03302_),
    .X(_03309_));
 sky130_fd_sc_hd__a32o_1 _19564_ (.A1(_02544_),
    .A2(_03308_),
    .A3(_03309_),
    .B1(_09886_),
    .B2(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_03310_));
 sky130_fd_sc_hd__a31o_1 _19565_ (.A1(_09888_),
    .A2(_03300_),
    .A3(_03301_),
    .B1(_03310_),
    .X(_00958_));
 sky130_fd_sc_hd__buf_2 _19566_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_03311_));
 sky130_fd_sc_hd__buf_2 _19567_ (.A(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_4 _19568_ (.A(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__xnor2_1 _19569_ (.A(_03313_),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_03314_));
 sky130_fd_sc_hd__a21oi_1 _19570_ (.A1(_03297_),
    .A2(_03301_),
    .B1(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__a311oi_1 _19571_ (.A1(_03297_),
    .A2(_03301_),
    .A3(_03314_),
    .B1(_03315_),
    .C1(_08262_),
    .Y(_03316_));
 sky130_fd_sc_hd__xor2_1 _19572_ (.A(_03262_),
    .B(_03232_),
    .X(_03317_));
 sky130_fd_sc_hd__o31ai_1 _19573_ (.A1(_03289_),
    .A2(_03303_),
    .A3(_03304_),
    .B1(_03308_),
    .Y(_03318_));
 sky130_fd_sc_hd__xnor2_1 _19574_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__xnor2_1 _19575_ (.A(_03303_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__a21o_1 _19576_ (.A1(_08262_),
    .A2(_03320_),
    .B1(_09886_),
    .X(_03321_));
 sky130_fd_sc_hd__o22a_1 _19577_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(_02551_),
    .B1(_03316_),
    .B2(_03321_),
    .X(_00959_));
 sky130_fd_sc_hd__and2_1 _19578_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_03322_));
 sky130_fd_sc_hd__nor2_1 _19579_ (.A(_03311_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_03323_));
 sky130_fd_sc_hd__o21ai_1 _19580_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(_03311_),
    .Y(_03324_));
 sky130_fd_sc_hd__o21bai_1 _19581_ (.A1(_03311_),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1_N(_03301_),
    .Y(_03325_));
 sky130_fd_sc_hd__o211ai_1 _19582_ (.A1(_03322_),
    .A2(_03323_),
    .B1(_03324_),
    .C1(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__a211o_1 _19583_ (.A1(_03324_),
    .A2(_03325_),
    .B1(_03322_),
    .C1(_03323_),
    .X(_03327_));
 sky130_fd_sc_hd__or2_1 _19584_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_05226_),
    .X(_03328_));
 sky130_fd_sc_hd__nand2_1 _19585_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_05226_),
    .Y(_03329_));
 sky130_fd_sc_hd__and4bb_1 _19586_ (.A_N(_03262_),
    .B_N(_03232_),
    .C(_03328_),
    .D(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__a2bb2o_1 _19587_ (.A1_N(_03262_),
    .A2_N(_03232_),
    .B1(_03328_),
    .B2(_03329_),
    .X(_03331_));
 sky130_fd_sc_hd__and2b_1 _19588_ (.A_N(_03330_),
    .B(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__o21a_1 _19589_ (.A1(_03307_),
    .A2(_03317_),
    .B1(_03303_),
    .X(_03333_));
 sky130_fd_sc_hd__a21o_1 _19590_ (.A1(_03317_),
    .A2(_03318_),
    .B1(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__and2_1 _19591_ (.A(_03332_),
    .B(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__o21ai_1 _19592_ (.A1(_03332_),
    .A2(_03334_),
    .B1(_08261_),
    .Y(_03336_));
 sky130_fd_sc_hd__a2bb2o_1 _19593_ (.A1_N(_03335_),
    .A2_N(_03336_),
    .B1(\rbzero.wall_tracer.rayAddendY[3] ),
    .B2(_09880_),
    .X(_03337_));
 sky130_fd_sc_hd__a31o_1 _19594_ (.A1(_09888_),
    .A2(_03326_),
    .A3(_03327_),
    .B1(_03337_),
    .X(_00960_));
 sky130_fd_sc_hd__nand2_1 _19595_ (.A(_03313_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_03338_));
 sky130_fd_sc_hd__xor2_1 _19596_ (.A(_03311_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_03339_));
 sky130_fd_sc_hd__a21oi_1 _19597_ (.A1(_03338_),
    .A2(_03327_),
    .B1(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__a31o_1 _19598_ (.A1(_03338_),
    .A2(_03327_),
    .A3(_03339_),
    .B1(_04566_),
    .X(_03341_));
 sky130_fd_sc_hd__xor2_1 _19599_ (.A(_03284_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_03342_));
 sky130_fd_sc_hd__o21ai_1 _19600_ (.A1(_03330_),
    .A2(_03335_),
    .B1(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__or3_1 _19601_ (.A(_03330_),
    .B(_03335_),
    .C(_03342_),
    .X(_03344_));
 sky130_fd_sc_hd__and2_1 _19602_ (.A(_03343_),
    .B(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__xnor2_1 _19603_ (.A(_03328_),
    .B(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__o22a_1 _19604_ (.A1(_03340_),
    .A2(_03341_),
    .B1(_03346_),
    .B2(_04568_),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _19605_ (.A0(\rbzero.wall_tracer.rayAddendY[4] ),
    .A1(_03347_),
    .S(_02550_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _19606_ (.A(_03348_),
    .X(_00961_));
 sky130_fd_sc_hd__nor2_1 _19607_ (.A(_03311_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .Y(_03349_));
 sky130_fd_sc_hd__and2_1 _19608_ (.A(_03311_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_03350_));
 sky130_fd_sc_hd__o22a_1 _19609_ (.A1(_03284_),
    .A2(\rbzero.debug_overlay.vplaneY[-4] ),
    .B1(_03349_),
    .B2(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__nor4_1 _19610_ (.A(_03284_),
    .B(\rbzero.debug_overlay.vplaneY[-4] ),
    .C(_03349_),
    .D(_03350_),
    .Y(_03352_));
 sky130_fd_sc_hd__nor2_1 _19611_ (.A(_03351_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__a2bb2o_1 _19612_ (.A1_N(_03335_),
    .A2_N(_03342_),
    .B1(_03343_),
    .B2(_03328_),
    .X(_03354_));
 sky130_fd_sc_hd__xnor2_1 _19613_ (.A(_03353_),
    .B(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__a22o_1 _19614_ (.A1(\rbzero.wall_tracer.rayAddendY[5] ),
    .A2(_09879_),
    .B1(_03355_),
    .B2(_08261_),
    .X(_03356_));
 sky130_fd_sc_hd__or2b_1 _19615_ (.A(_03327_),
    .B_N(_03339_),
    .X(_03357_));
 sky130_fd_sc_hd__o21ai_1 _19616_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_03313_),
    .Y(_03358_));
 sky130_fd_sc_hd__and2_1 _19617_ (.A(_03311_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_03359_));
 sky130_fd_sc_hd__nor2_1 _19618_ (.A(_03311_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_03360_));
 sky130_fd_sc_hd__or2_1 _19619_ (.A(_03359_),
    .B(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__a21oi_1 _19620_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__and3_1 _19621_ (.A(_03361_),
    .B(_03357_),
    .C(_03358_),
    .X(_03363_));
 sky130_fd_sc_hd__or3b_1 _19622_ (.A(_03362_),
    .B(_03363_),
    .C_N(_09883_),
    .X(_03364_));
 sky130_fd_sc_hd__or2b_1 _19623_ (.A(_03356_),
    .B_N(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_1 _19624_ (.A(_03365_),
    .X(_00962_));
 sky130_fd_sc_hd__xor2_1 _19625_ (.A(_03312_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_03366_));
 sky130_fd_sc_hd__o21ai_1 _19626_ (.A1(_03359_),
    .A2(_03362_),
    .B1(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__o31a_1 _19627_ (.A1(_03359_),
    .A2(_03362_),
    .A3(_03366_),
    .B1(_04568_),
    .X(_03368_));
 sky130_fd_sc_hd__or2_1 _19628_ (.A(_03311_),
    .B(_03262_),
    .X(_03369_));
 sky130_fd_sc_hd__nand2_1 _19629_ (.A(_03312_),
    .B(_03262_),
    .Y(_03370_));
 sky130_fd_sc_hd__a21o_1 _19630_ (.A1(_03369_),
    .A2(_03370_),
    .B1(_03349_),
    .X(_03371_));
 sky130_fd_sc_hd__nand2_1 _19631_ (.A(_03262_),
    .B(_03349_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand2_1 _19632_ (.A(_03371_),
    .B(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__o21bai_1 _19633_ (.A1(_03351_),
    .A2(_03354_),
    .B1_N(_03352_),
    .Y(_03374_));
 sky130_fd_sc_hd__xnor2_1 _19634_ (.A(_03373_),
    .B(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__a22o_1 _19635_ (.A1(_03367_),
    .A2(_03368_),
    .B1(_03375_),
    .B2(_08261_),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _19636_ (.A0(\rbzero.wall_tracer.rayAddendY[6] ),
    .A1(_03376_),
    .S(_02550_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_1 _19637_ (.A(_03377_),
    .X(_00963_));
 sky130_fd_sc_hd__nand2_1 _19638_ (.A(_03312_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_03378_));
 sky130_fd_sc_hd__or2_1 _19639_ (.A(_03312_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_03379_));
 sky130_fd_sc_hd__nor3b_1 _19640_ (.A(_03361_),
    .B(_03357_),
    .C_N(_03366_),
    .Y(_03380_));
 sky130_fd_sc_hd__o41a_1 _19641_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .A3(\rbzero.wall_tracer.rayAddendY[4] ),
    .A4(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_03312_),
    .X(_03381_));
 sky130_fd_sc_hd__a211o_1 _19642_ (.A1(_03378_),
    .A2(_03379_),
    .B1(_03380_),
    .C1(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__o211ai_2 _19643_ (.A1(_03380_),
    .A2(_03381_),
    .B1(_03378_),
    .C1(_03379_),
    .Y(_03383_));
 sky130_fd_sc_hd__inv_2 _19644_ (.A(_03372_),
    .Y(_03384_));
 sky130_fd_sc_hd__and3_1 _19645_ (.A(_03371_),
    .B(_03372_),
    .C(_03374_),
    .X(_03385_));
 sky130_fd_sc_hd__nor2_1 _19646_ (.A(_03312_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .Y(_03386_));
 sky130_fd_sc_hd__and2_1 _19647_ (.A(_03312_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_03387_));
 sky130_fd_sc_hd__o21ai_1 _19648_ (.A1(_03386_),
    .A2(_03387_),
    .B1(_03369_),
    .Y(_03388_));
 sky130_fd_sc_hd__or3_1 _19649_ (.A(_03369_),
    .B(_03386_),
    .C(_03387_),
    .X(_03389_));
 sky130_fd_sc_hd__o211ai_2 _19650_ (.A1(_03384_),
    .A2(_03385_),
    .B1(_03388_),
    .C1(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__a211o_1 _19651_ (.A1(_03388_),
    .A2(_03389_),
    .B1(_03384_),
    .C1(_03385_),
    .X(_03391_));
 sky130_fd_sc_hd__a32o_1 _19652_ (.A1(_02544_),
    .A2(_03390_),
    .A3(_03391_),
    .B1(_09886_),
    .B2(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_03392_));
 sky130_fd_sc_hd__a31o_1 _19653_ (.A1(_09888_),
    .A2(_03382_),
    .A3(_03383_),
    .B1(_03392_),
    .X(_00964_));
 sky130_fd_sc_hd__xnor2_1 _19654_ (.A(_03312_),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_03393_));
 sky130_fd_sc_hd__a21oi_1 _19655_ (.A1(_03378_),
    .A2(_03383_),
    .B1(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__a31o_1 _19656_ (.A1(_03378_),
    .A2(_03383_),
    .A3(_03393_),
    .B1(_08261_),
    .X(_03395_));
 sky130_fd_sc_hd__nor2_1 _19657_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__inv_2 _19658_ (.A(_03284_),
    .Y(_03397_));
 sky130_fd_sc_hd__a21oi_1 _19659_ (.A1(_03284_),
    .A2(\rbzero.debug_overlay.vplaneY[-1] ),
    .B1(_03312_),
    .Y(_03398_));
 sky130_fd_sc_hd__a21oi_1 _19660_ (.A1(_03313_),
    .A2(_03284_),
    .B1(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__a21oi_1 _19661_ (.A1(_03397_),
    .A2(_03386_),
    .B1(_03399_),
    .Y(_03400_));
 sky130_fd_sc_hd__a21o_1 _19662_ (.A1(_03389_),
    .A2(_03390_),
    .B1(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__nand3_1 _19663_ (.A(_03389_),
    .B(_03390_),
    .C(_03400_),
    .Y(_03402_));
 sky130_fd_sc_hd__a31o_1 _19664_ (.A1(_02544_),
    .A2(_03401_),
    .A3(_03402_),
    .B1(_09880_),
    .X(_03403_));
 sky130_fd_sc_hd__o22a_1 _19665_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(_02551_),
    .B1(_03396_),
    .B2(_03403_),
    .X(_00965_));
 sky130_fd_sc_hd__or2_1 _19666_ (.A(_03313_),
    .B(_03284_),
    .X(_03404_));
 sky130_fd_sc_hd__mux2_1 _19667_ (.A0(_03404_),
    .A1(_03398_),
    .S(_03401_),
    .X(_03405_));
 sky130_fd_sc_hd__or2_1 _19668_ (.A(_03313_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_03406_));
 sky130_fd_sc_hd__nand2_1 _19669_ (.A(_03313_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _19670_ (.A(_03406_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__o21ai_1 _19671_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(\rbzero.wall_tracer.rayAddendY[7] ),
    .B1(_03313_),
    .Y(_03409_));
 sky130_fd_sc_hd__o21ai_1 _19672_ (.A1(_03383_),
    .A2(_03393_),
    .B1(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__xor2_1 _19673_ (.A(_03408_),
    .B(_03410_),
    .X(_03411_));
 sky130_fd_sc_hd__o2bb2a_1 _19674_ (.A1_N(_02633_),
    .A2_N(_03411_),
    .B1(\rbzero.wall_tracer.rayAddendY[9] ),
    .B2(_02550_),
    .X(_03412_));
 sky130_fd_sc_hd__o21a_1 _19675_ (.A1(_04576_),
    .A2(_03405_),
    .B1(_03412_),
    .X(_00966_));
 sky130_fd_sc_hd__a21bo_1 _19676_ (.A1(_03406_),
    .A2(_03410_),
    .B1_N(_03407_),
    .X(_03413_));
 sky130_fd_sc_hd__xnor2_1 _19677_ (.A(_03313_),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_1 _19678_ (.A(_03413_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__inv_2 _19679_ (.A(_03313_),
    .Y(_03416_));
 sky130_fd_sc_hd__o211a_1 _19680_ (.A1(_03284_),
    .A2(_03401_),
    .B1(_08261_),
    .C1(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__o22a_1 _19681_ (.A1(_02539_),
    .A2(_03415_),
    .B1(_03417_),
    .B2(_09888_),
    .X(_03418_));
 sky130_fd_sc_hd__a21o_1 _19682_ (.A1(\rbzero.wall_tracer.rayAddendY[10] ),
    .A2(_09882_),
    .B1(_03418_),
    .X(_00967_));
 sky130_fd_sc_hd__nor2_2 _19683_ (.A(net41),
    .B(net40),
    .Y(_03419_));
 sky130_fd_sc_hd__and2_4 _19684_ (.A(\rbzero.pov.ready ),
    .B(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__o21ai_4 _19685_ (.A1(net40),
    .A2(_03420_),
    .B1(_02859_),
    .Y(_03421_));
 sky130_fd_sc_hd__buf_2 _19686_ (.A(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__inv_2 _19687_ (.A(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_03423_));
 sky130_fd_sc_hd__nor2_4 _19688_ (.A(_02881_),
    .B(_03419_),
    .Y(_03424_));
 sky130_fd_sc_hd__mux2_1 _19689_ (.A0(\rbzero.pov.ready_buffer[59] ),
    .A1(_03423_),
    .S(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__nand2_1 _19690_ (.A(_03423_),
    .B(_03422_),
    .Y(_03426_));
 sky130_fd_sc_hd__o211a_1 _19691_ (.A1(_03422_),
    .A2(_03425_),
    .B1(_03426_),
    .C1(_03069_),
    .X(_00968_));
 sky130_fd_sc_hd__or2_2 _19692_ (.A(net41),
    .B(net40),
    .X(_03427_));
 sky130_fd_sc_hd__nand2_1 _19693_ (.A(_02859_),
    .B(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__clkbuf_4 _19694_ (.A(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__buf_2 _19695_ (.A(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nand2_1 _19696_ (.A(\rbzero.pov.ready_buffer[60] ),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__o21ai_1 _19697_ (.A1(_08275_),
    .A2(_03430_),
    .B1(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__o21a_1 _19698_ (.A1(net40),
    .A2(_03420_),
    .B1(_02859_),
    .X(_03433_));
 sky130_fd_sc_hd__buf_2 _19699_ (.A(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__or2_1 _19700_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__o211a_1 _19701_ (.A1(_03422_),
    .A2(_03432_),
    .B1(_03435_),
    .C1(_03069_),
    .X(_00969_));
 sky130_fd_sc_hd__clkbuf_4 _19702_ (.A(_03428_),
    .X(_03436_));
 sky130_fd_sc_hd__nor2_1 _19703_ (.A(_08309_),
    .B(_03429_),
    .Y(_03437_));
 sky130_fd_sc_hd__a211o_1 _19704_ (.A1(\rbzero.pov.ready_buffer[61] ),
    .A2(_03436_),
    .B1(_03437_),
    .C1(_03421_),
    .X(_03438_));
 sky130_fd_sc_hd__o211a_1 _19705_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_03434_),
    .B1(_03438_),
    .C1(_03069_),
    .X(_00970_));
 sky130_fd_sc_hd__nor2_1 _19706_ (.A(_08333_),
    .B(_03429_),
    .Y(_03439_));
 sky130_fd_sc_hd__a211o_1 _19707_ (.A1(\rbzero.pov.ready_buffer[62] ),
    .A2(_03436_),
    .B1(_03439_),
    .C1(_03421_),
    .X(_03440_));
 sky130_fd_sc_hd__o211a_1 _19708_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_03434_),
    .B1(_03440_),
    .C1(_03069_),
    .X(_00971_));
 sky130_fd_sc_hd__nand2_1 _19709_ (.A(\rbzero.pov.ready_buffer[63] ),
    .B(_03430_),
    .Y(_03441_));
 sky130_fd_sc_hd__o21ai_1 _19710_ (.A1(_08445_),
    .A2(_03430_),
    .B1(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__or2_1 _19711_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_03434_),
    .X(_03443_));
 sky130_fd_sc_hd__o211a_1 _19712_ (.A1(_03422_),
    .A2(_03442_),
    .B1(_03443_),
    .C1(_03069_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _19713_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(_08455_),
    .S(_03424_),
    .X(_03444_));
 sky130_fd_sc_hd__nand2_1 _19714_ (.A(_08456_),
    .B(_03422_),
    .Y(_03445_));
 sky130_fd_sc_hd__o211a_1 _19715_ (.A1(_03422_),
    .A2(_03444_),
    .B1(_03445_),
    .C1(_03069_),
    .X(_00973_));
 sky130_fd_sc_hd__nor2_1 _19716_ (.A(_08476_),
    .B(_03429_),
    .Y(_03446_));
 sky130_fd_sc_hd__a211o_1 _19717_ (.A1(\rbzero.pov.ready_buffer[65] ),
    .A2(_03436_),
    .B1(_03446_),
    .C1(_03421_),
    .X(_03447_));
 sky130_fd_sc_hd__o211a_1 _19718_ (.A1(\rbzero.debug_overlay.playerX[-3] ),
    .A2(_03434_),
    .B1(_03447_),
    .C1(_03069_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _19719_ (.A0(\rbzero.pov.ready_buffer[66] ),
    .A1(_08584_),
    .S(_03424_),
    .X(_03448_));
 sky130_fd_sc_hd__or2_1 _19720_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_03434_),
    .X(_03449_));
 sky130_fd_sc_hd__buf_2 _19721_ (.A(_02973_),
    .X(_03450_));
 sky130_fd_sc_hd__o211a_1 _19722_ (.A1(_03422_),
    .A2(_03448_),
    .B1(_03449_),
    .C1(_03450_),
    .X(_00975_));
 sky130_fd_sc_hd__a21o_1 _19723_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_03421_),
    .B1(_04544_),
    .X(_03451_));
 sky130_fd_sc_hd__o221a_1 _19724_ (.A1(\rbzero.pov.ready_buffer[67] ),
    .A2(_03427_),
    .B1(_03429_),
    .B2(_08572_),
    .C1(_03433_),
    .X(_03452_));
 sky130_fd_sc_hd__or2_1 _19725_ (.A(_03451_),
    .B(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _19726_ (.A(_03453_),
    .X(_00976_));
 sky130_fd_sc_hd__clkbuf_4 _19727_ (.A(_03424_),
    .X(_03454_));
 sky130_fd_sc_hd__or2_1 _19728_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_08570_),
    .X(_03455_));
 sky130_fd_sc_hd__inv_2 _19729_ (.A(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__a21o_1 _19730_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_08570_),
    .B1(_03428_),
    .X(_03457_));
 sky130_fd_sc_hd__o221a_1 _19731_ (.A1(\rbzero.pov.ready_buffer[68] ),
    .A2(_03454_),
    .B1(_03456_),
    .B2(_03457_),
    .C1(_03434_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_4 _19732_ (.A(_04545_),
    .X(_03459_));
 sky130_fd_sc_hd__a211o_1 _19733_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03422_),
    .B1(_03458_),
    .C1(_03459_),
    .X(_00977_));
 sky130_fd_sc_hd__nor2_1 _19734_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03455_),
    .Y(_03460_));
 sky130_fd_sc_hd__a21o_1 _19735_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03455_),
    .B1(_03428_),
    .X(_03461_));
 sky130_fd_sc_hd__o221a_1 _19736_ (.A1(\rbzero.pov.ready_buffer[69] ),
    .A2(_03454_),
    .B1(_03460_),
    .B2(_03461_),
    .C1(_03434_),
    .X(_03462_));
 sky130_fd_sc_hd__a211o_1 _19737_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03422_),
    .B1(_03462_),
    .C1(_03459_),
    .X(_00978_));
 sky130_fd_sc_hd__nand2_1 _19738_ (.A(_04804_),
    .B(_03460_),
    .Y(_03463_));
 sky130_fd_sc_hd__or2_1 _19739_ (.A(_04804_),
    .B(_03460_),
    .X(_03464_));
 sky130_fd_sc_hd__a21oi_1 _19740_ (.A1(_03463_),
    .A2(_03464_),
    .B1(_03429_),
    .Y(_03465_));
 sky130_fd_sc_hd__a211o_1 _19741_ (.A1(\rbzero.pov.ready_buffer[70] ),
    .A2(_03436_),
    .B1(_03465_),
    .C1(_03421_),
    .X(_03466_));
 sky130_fd_sc_hd__o211a_1 _19742_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_03434_),
    .B1(_03466_),
    .C1(_03450_),
    .X(_00979_));
 sky130_fd_sc_hd__or2_1 _19743_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_03463_),
    .X(_03467_));
 sky130_fd_sc_hd__and2_1 _19744_ (.A(_03427_),
    .B(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__inv_2 _19745_ (.A(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hd__a21o_1 _19746_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03463_),
    .B1(_02881_),
    .X(_03470_));
 sky130_fd_sc_hd__o221a_1 _19747_ (.A1(\rbzero.pov.ready_buffer[71] ),
    .A2(_03454_),
    .B1(_03469_),
    .B2(_03470_),
    .C1(_03434_),
    .X(_03471_));
 sky130_fd_sc_hd__a211o_1 _19748_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03422_),
    .B1(_03471_),
    .C1(_03459_),
    .X(_00980_));
 sky130_fd_sc_hd__o21a_1 _19749_ (.A1(_03421_),
    .A2(_03468_),
    .B1(\rbzero.debug_overlay.playerX[4] ),
    .X(_03472_));
 sky130_fd_sc_hd__nor2_1 _19750_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_03467_),
    .Y(_03473_));
 sky130_fd_sc_hd__o21ai_1 _19751_ (.A1(_03419_),
    .A2(_03473_),
    .B1(_03433_),
    .Y(_03474_));
 sky130_fd_sc_hd__o21ba_1 _19752_ (.A1(\rbzero.pov.ready_buffer[72] ),
    .A2(_03454_),
    .B1_N(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__o21a_1 _19753_ (.A1(_03472_),
    .A2(_03475_),
    .B1(_02868_),
    .X(_00981_));
 sky130_fd_sc_hd__o31ai_1 _19754_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(\rbzero.debug_overlay.playerX[4] ),
    .A3(_03467_),
    .B1(_03424_),
    .Y(_03476_));
 sky130_fd_sc_hd__o211a_1 _19755_ (.A1(\rbzero.pov.ready_buffer[73] ),
    .A2(_03424_),
    .B1(_03476_),
    .C1(_03433_),
    .X(_03477_));
 sky130_fd_sc_hd__a21oi_1 _19756_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_03474_),
    .B1(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__nor2_1 _19757_ (.A(_03459_),
    .B(_03478_),
    .Y(_00982_));
 sky130_fd_sc_hd__o21ai_4 _19758_ (.A1(net41),
    .A2(_03420_),
    .B1(_02859_),
    .Y(_03479_));
 sky130_fd_sc_hd__clkbuf_4 _19759_ (.A(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _19760_ (.A0(\rbzero.pov.ready_buffer[44] ),
    .A1(_08363_),
    .S(_03424_),
    .X(_03481_));
 sky130_fd_sc_hd__nand2_1 _19761_ (.A(_08363_),
    .B(_03480_),
    .Y(_03482_));
 sky130_fd_sc_hd__o211a_1 _19762_ (.A1(_03480_),
    .A2(_03481_),
    .B1(_03482_),
    .C1(_03450_),
    .X(_00983_));
 sky130_fd_sc_hd__nand2_1 _19763_ (.A(\rbzero.pov.ready_buffer[45] ),
    .B(_03430_),
    .Y(_03483_));
 sky130_fd_sc_hd__o21ai_1 _19764_ (.A1(_08283_),
    .A2(_03430_),
    .B1(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__o21a_1 _19765_ (.A1(net41),
    .A2(_03420_),
    .B1(_02859_),
    .X(_03485_));
 sky130_fd_sc_hd__or2_1 _19766_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__o211a_1 _19767_ (.A1(_03480_),
    .A2(_03484_),
    .B1(_03486_),
    .C1(_03450_),
    .X(_00984_));
 sky130_fd_sc_hd__buf_2 _19768_ (.A(_03485_),
    .X(_03487_));
 sky130_fd_sc_hd__nor2_1 _19769_ (.A(_08313_),
    .B(_03436_),
    .Y(_03488_));
 sky130_fd_sc_hd__a211o_1 _19770_ (.A1(\rbzero.pov.ready_buffer[46] ),
    .A2(_03436_),
    .B1(_03479_),
    .C1(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__o211a_1 _19771_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_03487_),
    .B1(_03489_),
    .C1(_03450_),
    .X(_00985_));
 sky130_fd_sc_hd__nor2_1 _19772_ (.A(_08338_),
    .B(_03429_),
    .Y(_03490_));
 sky130_fd_sc_hd__a211o_1 _19773_ (.A1(\rbzero.pov.ready_buffer[47] ),
    .A2(_03436_),
    .B1(_03479_),
    .C1(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__o211a_1 _19774_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_03487_),
    .B1(_03491_),
    .C1(_03450_),
    .X(_00986_));
 sky130_fd_sc_hd__nand2_1 _19775_ (.A(\rbzero.pov.ready_buffer[48] ),
    .B(_03430_),
    .Y(_03492_));
 sky130_fd_sc_hd__o21ai_1 _19776_ (.A1(_08447_),
    .A2(_03430_),
    .B1(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__or2_1 _19777_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_03485_),
    .X(_03494_));
 sky130_fd_sc_hd__o211a_1 _19778_ (.A1(_03480_),
    .A2(_03493_),
    .B1(_03494_),
    .C1(_03450_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _19779_ (.A0(\rbzero.pov.ready_buffer[49] ),
    .A1(_08460_),
    .S(_03424_),
    .X(_03495_));
 sky130_fd_sc_hd__nand2_1 _19780_ (.A(_08461_),
    .B(_03480_),
    .Y(_03496_));
 sky130_fd_sc_hd__o211a_1 _19781_ (.A1(_03480_),
    .A2(_03495_),
    .B1(_03496_),
    .C1(_03450_),
    .X(_00988_));
 sky130_fd_sc_hd__nor2_1 _19782_ (.A(_08480_),
    .B(_03429_),
    .Y(_03497_));
 sky130_fd_sc_hd__a211o_1 _19783_ (.A1(\rbzero.pov.ready_buffer[50] ),
    .A2(_03436_),
    .B1(_03479_),
    .C1(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__o211a_1 _19784_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_03487_),
    .B1(_03498_),
    .C1(_03450_),
    .X(_00989_));
 sky130_fd_sc_hd__nand2_1 _19785_ (.A(\rbzero.pov.ready_buffer[51] ),
    .B(_03436_),
    .Y(_03499_));
 sky130_fd_sc_hd__o211ai_1 _19786_ (.A1(_08581_),
    .A2(_03430_),
    .B1(_03487_),
    .C1(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__o211a_1 _19787_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_03487_),
    .B1(_03500_),
    .C1(_03450_),
    .X(_00990_));
 sky130_fd_sc_hd__o21ai_1 _19788_ (.A1(\rbzero.pov.ready_buffer[52] ),
    .A2(_03427_),
    .B1(_03485_),
    .Y(_03501_));
 sky130_fd_sc_hd__a21oi_1 _19789_ (.A1(_08576_),
    .A2(_03454_),
    .B1(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__a211o_1 _19790_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_03480_),
    .B1(_03502_),
    .C1(_03459_),
    .X(_00991_));
 sky130_fd_sc_hd__or2_1 _19791_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08574_),
    .X(_03503_));
 sky130_fd_sc_hd__nand2_1 _19792_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08574_),
    .Y(_03504_));
 sky130_fd_sc_hd__a21oi_1 _19793_ (.A1(_03503_),
    .A2(_03504_),
    .B1(_03429_),
    .Y(_03505_));
 sky130_fd_sc_hd__a211o_1 _19794_ (.A1(\rbzero.pov.ready_buffer[53] ),
    .A2(_03436_),
    .B1(_03479_),
    .C1(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_4 _19795_ (.A(_02973_),
    .X(_03507_));
 sky130_fd_sc_hd__o211a_1 _19796_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_03487_),
    .B1(_03506_),
    .C1(_03507_),
    .X(_00992_));
 sky130_fd_sc_hd__and2_1 _19797_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(_03503_),
    .X(_03508_));
 sky130_fd_sc_hd__o21ai_1 _19798_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03503_),
    .B1(_03424_),
    .Y(_03509_));
 sky130_fd_sc_hd__o221a_1 _19799_ (.A1(\rbzero.pov.ready_buffer[54] ),
    .A2(_03454_),
    .B1(_03508_),
    .B2(_03509_),
    .C1(_03487_),
    .X(_03510_));
 sky130_fd_sc_hd__a211o_1 _19800_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03480_),
    .B1(_03510_),
    .C1(_03459_),
    .X(_00993_));
 sky130_fd_sc_hd__a21o_1 _19801_ (.A1(_03487_),
    .A2(_03509_),
    .B1(_06182_),
    .X(_03511_));
 sky130_fd_sc_hd__or3_1 _19802_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .C(_03503_),
    .X(_03512_));
 sky130_fd_sc_hd__nor2_1 _19803_ (.A(\rbzero.pov.ready_buffer[55] ),
    .B(_03424_),
    .Y(_03513_));
 sky130_fd_sc_hd__a211o_1 _19804_ (.A1(_03454_),
    .A2(_03512_),
    .B1(_03513_),
    .C1(_03479_),
    .X(_03514_));
 sky130_fd_sc_hd__a21oi_1 _19805_ (.A1(_03511_),
    .A2(_03514_),
    .B1(_03459_),
    .Y(_00994_));
 sky130_fd_sc_hd__o21a_1 _19806_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03512_),
    .B1(_03427_),
    .X(_03515_));
 sky130_fd_sc_hd__inv_2 _19807_ (.A(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__a21o_1 _19808_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03512_),
    .B1(_02881_),
    .X(_03517_));
 sky130_fd_sc_hd__o221a_1 _19809_ (.A1(\rbzero.pov.ready_buffer[56] ),
    .A2(_03454_),
    .B1(_03516_),
    .B2(_03517_),
    .C1(_03487_),
    .X(_03518_));
 sky130_fd_sc_hd__a211o_1 _19810_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03480_),
    .B1(_03518_),
    .C1(_03459_),
    .X(_00995_));
 sky130_fd_sc_hd__o21a_1 _19811_ (.A1(_03480_),
    .A2(_03515_),
    .B1(\rbzero.debug_overlay.playerY[4] ),
    .X(_03519_));
 sky130_fd_sc_hd__and3b_1 _19812_ (.A_N(_03512_),
    .B(_04809_),
    .C(_04803_),
    .X(_03520_));
 sky130_fd_sc_hd__o21a_1 _19813_ (.A1(_03419_),
    .A2(_03520_),
    .B1(_03485_),
    .X(_03521_));
 sky130_fd_sc_hd__o21a_1 _19814_ (.A1(\rbzero.pov.ready_buffer[57] ),
    .A2(_03454_),
    .B1(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__o21a_1 _19815_ (.A1(_03519_),
    .A2(_03522_),
    .B1(_02868_),
    .X(_00996_));
 sky130_fd_sc_hd__nor2_1 _19816_ (.A(_06185_),
    .B(_03521_),
    .Y(_03523_));
 sky130_fd_sc_hd__a21o_1 _19817_ (.A1(_06185_),
    .A2(_03520_),
    .B1(_03429_),
    .X(_03524_));
 sky130_fd_sc_hd__o211a_1 _19818_ (.A1(\rbzero.pov.ready_buffer[58] ),
    .A2(_03454_),
    .B1(_03487_),
    .C1(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__o21a_1 _19819_ (.A1(_03523_),
    .A2(_03525_),
    .B1(_02868_),
    .X(_00997_));
 sky130_fd_sc_hd__nand2_1 _19820_ (.A(_02859_),
    .B(_03420_),
    .Y(_03526_));
 sky130_fd_sc_hd__buf_2 _19821_ (.A(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__buf_2 _19822_ (.A(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__and2_1 _19823_ (.A(_02859_),
    .B(_03420_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_2 _19824_ (.A(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__or2_1 _19825_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__o211a_1 _19826_ (.A1(\rbzero.pov.ready_buffer[33] ),
    .A2(_03528_),
    .B1(_03531_),
    .C1(_03507_),
    .X(_00998_));
 sky130_fd_sc_hd__or2_1 _19827_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(_03530_),
    .X(_03532_));
 sky130_fd_sc_hd__o211a_1 _19828_ (.A1(\rbzero.pov.ready_buffer[34] ),
    .A2(_03528_),
    .B1(_03532_),
    .C1(_03507_),
    .X(_00999_));
 sky130_fd_sc_hd__or2_1 _19829_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(_03530_),
    .X(_03533_));
 sky130_fd_sc_hd__o211a_1 _19830_ (.A1(\rbzero.pov.ready_buffer[35] ),
    .A2(_03528_),
    .B1(_03533_),
    .C1(_03507_),
    .X(_01000_));
 sky130_fd_sc_hd__or2_1 _19831_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(_03530_),
    .X(_03534_));
 sky130_fd_sc_hd__o211a_1 _19832_ (.A1(\rbzero.pov.ready_buffer[36] ),
    .A2(_03528_),
    .B1(_03534_),
    .C1(_03507_),
    .X(_01001_));
 sky130_fd_sc_hd__buf_4 _19833_ (.A(_03526_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_2 _19834_ (.A(_03420_),
    .X(_03536_));
 sky130_fd_sc_hd__clkbuf_2 _19835_ (.A(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__and3_1 _19836_ (.A(\rbzero.pov.ready_buffer[37] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03538_));
 sky130_fd_sc_hd__a211o_1 _19837_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_03535_),
    .B1(_03538_),
    .C1(_03459_),
    .X(_01002_));
 sky130_fd_sc_hd__and3_1 _19838_ (.A(\rbzero.pov.ready_buffer[38] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03539_));
 sky130_fd_sc_hd__a211o_1 _19839_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_03535_),
    .B1(_03539_),
    .C1(_03459_),
    .X(_01003_));
 sky130_fd_sc_hd__and3_1 _19840_ (.A(\rbzero.pov.ready_buffer[39] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_4 _19841_ (.A(_04545_),
    .X(_03541_));
 sky130_fd_sc_hd__a211o_1 _19842_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_03535_),
    .B1(_03540_),
    .C1(_03541_),
    .X(_01004_));
 sky130_fd_sc_hd__or2_1 _19843_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(_03530_),
    .X(_03542_));
 sky130_fd_sc_hd__o211a_1 _19844_ (.A1(\rbzero.pov.ready_buffer[40] ),
    .A2(_03528_),
    .B1(_03542_),
    .C1(_03507_),
    .X(_01005_));
 sky130_fd_sc_hd__and3_1 _19845_ (.A(\rbzero.pov.ready_buffer[41] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03543_));
 sky130_fd_sc_hd__a211o_1 _19846_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(_03535_),
    .B1(_03543_),
    .C1(_03541_),
    .X(_01006_));
 sky130_fd_sc_hd__or2_1 _19847_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(_03530_),
    .X(_03544_));
 sky130_fd_sc_hd__o211a_1 _19848_ (.A1(\rbzero.pov.ready_buffer[42] ),
    .A2(_03528_),
    .B1(_03544_),
    .C1(_03507_),
    .X(_01007_));
 sky130_fd_sc_hd__or2_1 _19849_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(_03530_),
    .X(_03545_));
 sky130_fd_sc_hd__o211a_1 _19850_ (.A1(\rbzero.pov.ready_buffer[43] ),
    .A2(_03528_),
    .B1(_03545_),
    .C1(_03507_),
    .X(_01008_));
 sky130_fd_sc_hd__and3_1 _19851_ (.A(\rbzero.pov.ready_buffer[22] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03546_));
 sky130_fd_sc_hd__a211o_1 _19852_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(_03535_),
    .B1(_03546_),
    .C1(_03541_),
    .X(_01009_));
 sky130_fd_sc_hd__or2_1 _19853_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_03530_),
    .X(_03547_));
 sky130_fd_sc_hd__o211a_1 _19854_ (.A1(\rbzero.pov.ready_buffer[23] ),
    .A2(_03528_),
    .B1(_03547_),
    .C1(_03507_),
    .X(_01010_));
 sky130_fd_sc_hd__buf_2 _19855_ (.A(_03526_),
    .X(_03548_));
 sky130_fd_sc_hd__and3_1 _19856_ (.A(\rbzero.pov.ready_buffer[24] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03549_));
 sky130_fd_sc_hd__a211o_1 _19857_ (.A1(\rbzero.debug_overlay.facingY[-7] ),
    .A2(_03548_),
    .B1(_03549_),
    .C1(_03541_),
    .X(_01011_));
 sky130_fd_sc_hd__and3_1 _19858_ (.A(\rbzero.pov.ready_buffer[25] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03550_));
 sky130_fd_sc_hd__a211o_1 _19859_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_03548_),
    .B1(_03550_),
    .C1(_03541_),
    .X(_01012_));
 sky130_fd_sc_hd__and3_1 _19860_ (.A(\rbzero.pov.ready_buffer[26] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03551_));
 sky130_fd_sc_hd__a211o_1 _19861_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_03548_),
    .B1(_03551_),
    .C1(_03541_),
    .X(_01013_));
 sky130_fd_sc_hd__or2_1 _19862_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(_03530_),
    .X(_03552_));
 sky130_fd_sc_hd__o211a_1 _19863_ (.A1(\rbzero.pov.ready_buffer[27] ),
    .A2(_03528_),
    .B1(_03552_),
    .C1(_03507_),
    .X(_01014_));
 sky130_fd_sc_hd__or2_1 _19864_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(_03530_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_4 _19865_ (.A(_02867_),
    .X(_03554_));
 sky130_fd_sc_hd__o211a_1 _19866_ (.A1(\rbzero.pov.ready_buffer[28] ),
    .A2(_03528_),
    .B1(_03553_),
    .C1(_03554_),
    .X(_01015_));
 sky130_fd_sc_hd__and3_1 _19867_ (.A(\rbzero.pov.ready_buffer[29] ),
    .B(_02923_),
    .C(_03537_),
    .X(_03555_));
 sky130_fd_sc_hd__a211o_1 _19868_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(_03548_),
    .B1(_03555_),
    .C1(_03541_),
    .X(_01016_));
 sky130_fd_sc_hd__clkbuf_4 _19869_ (.A(_03526_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_2 _19870_ (.A(_03529_),
    .X(_03557_));
 sky130_fd_sc_hd__or2_1 _19871_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__o211a_1 _19872_ (.A1(\rbzero.pov.ready_buffer[30] ),
    .A2(_03556_),
    .B1(_03558_),
    .C1(_03554_),
    .X(_01017_));
 sky130_fd_sc_hd__clkbuf_2 _19873_ (.A(_02860_),
    .X(_03559_));
 sky130_fd_sc_hd__and3_1 _19874_ (.A(\rbzero.pov.ready_buffer[31] ),
    .B(_03559_),
    .C(_03537_),
    .X(_03560_));
 sky130_fd_sc_hd__a211o_1 _19875_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_03548_),
    .B1(_03560_),
    .C1(_03541_),
    .X(_01018_));
 sky130_fd_sc_hd__and3_1 _19876_ (.A(\rbzero.pov.ready_buffer[32] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03561_));
 sky130_fd_sc_hd__a211o_1 _19877_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_03548_),
    .B1(_03561_),
    .C1(_03541_),
    .X(_01019_));
 sky130_fd_sc_hd__and3_1 _19878_ (.A(\rbzero.pov.ready_buffer[11] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03562_));
 sky130_fd_sc_hd__a211o_1 _19879_ (.A1(_02538_),
    .A2(_03548_),
    .B1(_03562_),
    .C1(_03541_),
    .X(_01020_));
 sky130_fd_sc_hd__or2_1 _19880_ (.A(_05246_),
    .B(_03557_),
    .X(_03563_));
 sky130_fd_sc_hd__o211a_1 _19881_ (.A1(\rbzero.pov.ready_buffer[12] ),
    .A2(_03556_),
    .B1(_03563_),
    .C1(_03554_),
    .X(_01021_));
 sky130_fd_sc_hd__or2_1 _19882_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_03557_),
    .X(_03564_));
 sky130_fd_sc_hd__o211a_1 _19883_ (.A1(\rbzero.pov.ready_buffer[13] ),
    .A2(_03556_),
    .B1(_03564_),
    .C1(_03554_),
    .X(_01022_));
 sky130_fd_sc_hd__or2_1 _19884_ (.A(_02526_),
    .B(_03557_),
    .X(_03565_));
 sky130_fd_sc_hd__o211a_1 _19885_ (.A1(\rbzero.pov.ready_buffer[14] ),
    .A2(_03556_),
    .B1(_03565_),
    .C1(_03554_),
    .X(_01023_));
 sky130_fd_sc_hd__and3_1 _19886_ (.A(\rbzero.pov.ready_buffer[15] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_4 _19887_ (.A(_04545_),
    .X(_03567_));
 sky130_fd_sc_hd__a211o_1 _19888_ (.A1(_05249_),
    .A2(_03548_),
    .B1(_03566_),
    .C1(_03567_),
    .X(_01024_));
 sky130_fd_sc_hd__and3_1 _19889_ (.A(\rbzero.pov.ready_buffer[16] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03568_));
 sky130_fd_sc_hd__a211o_1 _19890_ (.A1(\rbzero.debug_overlay.vplaneX[-4] ),
    .A2(_03548_),
    .B1(_03568_),
    .C1(_03567_),
    .X(_01025_));
 sky130_fd_sc_hd__or2_1 _19891_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(_03557_),
    .X(_03569_));
 sky130_fd_sc_hd__o211a_1 _19892_ (.A1(\rbzero.pov.ready_buffer[17] ),
    .A2(_03556_),
    .B1(_03569_),
    .C1(_03554_),
    .X(_01026_));
 sky130_fd_sc_hd__and3_1 _19893_ (.A(\rbzero.pov.ready_buffer[18] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03570_));
 sky130_fd_sc_hd__a211o_1 _19894_ (.A1(\rbzero.debug_overlay.vplaneX[-2] ),
    .A2(_03548_),
    .B1(_03570_),
    .C1(_03567_),
    .X(_01027_));
 sky130_fd_sc_hd__or2_1 _19895_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_03557_),
    .X(_03571_));
 sky130_fd_sc_hd__o211a_1 _19896_ (.A1(\rbzero.pov.ready_buffer[19] ),
    .A2(_03556_),
    .B1(_03571_),
    .C1(_03554_),
    .X(_01028_));
 sky130_fd_sc_hd__nand2_1 _19897_ (.A(_02704_),
    .B(_03527_),
    .Y(_03572_));
 sky130_fd_sc_hd__o211a_1 _19898_ (.A1(\rbzero.pov.ready_buffer[20] ),
    .A2(_03556_),
    .B1(_03572_),
    .C1(_03554_),
    .X(_01029_));
 sky130_fd_sc_hd__nand2_1 _19899_ (.A(_02723_),
    .B(_03527_),
    .Y(_03573_));
 sky130_fd_sc_hd__o211a_1 _19900_ (.A1(\rbzero.pov.ready_buffer[21] ),
    .A2(_03556_),
    .B1(_03573_),
    .C1(_03554_),
    .X(_01030_));
 sky130_fd_sc_hd__nand2_1 _19901_ (.A(_03279_),
    .B(_03527_),
    .Y(_03574_));
 sky130_fd_sc_hd__o211a_1 _19902_ (.A1(\rbzero.pov.ready_buffer[0] ),
    .A2(_03556_),
    .B1(_03574_),
    .C1(_03554_),
    .X(_01031_));
 sky130_fd_sc_hd__or2_1 _19903_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_03557_),
    .X(_03575_));
 sky130_fd_sc_hd__buf_2 _19904_ (.A(_02867_),
    .X(_03576_));
 sky130_fd_sc_hd__o211a_1 _19905_ (.A1(\rbzero.pov.ready_buffer[1] ),
    .A2(_03556_),
    .B1(_03575_),
    .C1(_03576_),
    .X(_01032_));
 sky130_fd_sc_hd__or2_1 _19906_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03557_),
    .X(_03577_));
 sky130_fd_sc_hd__o211a_1 _19907_ (.A1(\rbzero.pov.ready_buffer[2] ),
    .A2(_03535_),
    .B1(_03577_),
    .C1(_03576_),
    .X(_01033_));
 sky130_fd_sc_hd__and3_1 _19908_ (.A(\rbzero.pov.ready_buffer[3] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03578_));
 sky130_fd_sc_hd__a211o_1 _19909_ (.A1(_03232_),
    .A2(_03527_),
    .B1(_03578_),
    .C1(_03567_),
    .X(_01034_));
 sky130_fd_sc_hd__and3_1 _19910_ (.A(\rbzero.pov.ready_buffer[4] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03579_));
 sky130_fd_sc_hd__a211o_1 _19911_ (.A1(_05226_),
    .A2(_03527_),
    .B1(_03579_),
    .C1(_03567_),
    .X(_01035_));
 sky130_fd_sc_hd__and3_1 _19912_ (.A(\rbzero.pov.ready_buffer[5] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03580_));
 sky130_fd_sc_hd__a211o_1 _19913_ (.A1(\rbzero.debug_overlay.vplaneY[-4] ),
    .A2(_03527_),
    .B1(_03580_),
    .C1(_03567_),
    .X(_01036_));
 sky130_fd_sc_hd__or2_1 _19914_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(_03557_),
    .X(_03581_));
 sky130_fd_sc_hd__o211a_1 _19915_ (.A1(\rbzero.pov.ready_buffer[6] ),
    .A2(_03535_),
    .B1(_03581_),
    .C1(_03576_),
    .X(_01037_));
 sky130_fd_sc_hd__and3_1 _19916_ (.A(\rbzero.pov.ready_buffer[7] ),
    .B(_03559_),
    .C(_03536_),
    .X(_03582_));
 sky130_fd_sc_hd__a211o_1 _19917_ (.A1(_03262_),
    .A2(_03527_),
    .B1(_03582_),
    .C1(_03567_),
    .X(_01038_));
 sky130_fd_sc_hd__or2_1 _19918_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_03557_),
    .X(_03583_));
 sky130_fd_sc_hd__o211a_1 _19919_ (.A1(\rbzero.pov.ready_buffer[8] ),
    .A2(_03535_),
    .B1(_03583_),
    .C1(_03576_),
    .X(_01039_));
 sky130_fd_sc_hd__nand2_1 _19920_ (.A(_03397_),
    .B(_03527_),
    .Y(_03584_));
 sky130_fd_sc_hd__o211a_1 _19921_ (.A1(\rbzero.pov.ready_buffer[9] ),
    .A2(_03535_),
    .B1(_03584_),
    .C1(_03576_),
    .X(_01040_));
 sky130_fd_sc_hd__nand2_1 _19922_ (.A(_03416_),
    .B(_03527_),
    .Y(_03585_));
 sky130_fd_sc_hd__o211a_1 _19923_ (.A1(\rbzero.pov.ready_buffer[10] ),
    .A2(_03535_),
    .B1(_03585_),
    .C1(_03576_),
    .X(_01041_));
 sky130_fd_sc_hd__and2b_1 _19924_ (.A_N(\rbzero.pov.sclk_buffer[2] ),
    .B(\rbzero.pov.sclk_buffer[1] ),
    .X(_03586_));
 sky130_fd_sc_hd__and2_1 _19925_ (.A(\rbzero.pov.spi_counter[0] ),
    .B(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__nor2_2 _19926_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(_04544_),
    .Y(_03588_));
 sky130_fd_sc_hd__o21ai_1 _19927_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03586_),
    .B1(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__nor2_1 _19928_ (.A(_03587_),
    .B(_03589_),
    .Y(_01042_));
 sky130_fd_sc_hd__and3_1 _19929_ (.A(\rbzero.pov.spi_counter[1] ),
    .B(\rbzero.pov.spi_counter[0] ),
    .C(_03586_),
    .X(_03590_));
 sky130_fd_sc_hd__clkinv_2 _19930_ (.A(\rbzero.pov.spi_counter[6] ),
    .Y(_03591_));
 sky130_fd_sc_hd__or4b_1 _19931_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[2] ),
    .C(\rbzero.pov.spi_counter[1] ),
    .D_N(\rbzero.pov.spi_counter[3] ),
    .X(_03592_));
 sky130_fd_sc_hd__or4b_1 _19932_ (.A(_03591_),
    .B(_03592_),
    .C(\rbzero.pov.spi_counter[5] ),
    .D_N(_03587_),
    .X(_03593_));
 sky130_fd_sc_hd__and2_1 _19933_ (.A(_03588_),
    .B(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__o21ai_1 _19934_ (.A1(\rbzero.pov.spi_counter[1] ),
    .A2(_03587_),
    .B1(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__nor2_1 _19935_ (.A(_03590_),
    .B(_03595_),
    .Y(_01043_));
 sky130_fd_sc_hd__and3_1 _19936_ (.A(\rbzero.pov.spi_counter[2] ),
    .B(\rbzero.pov.spi_counter[1] ),
    .C(_03587_),
    .X(_03596_));
 sky130_fd_sc_hd__o21ai_1 _19937_ (.A1(\rbzero.pov.spi_counter[2] ),
    .A2(_03590_),
    .B1(_03588_),
    .Y(_03597_));
 sky130_fd_sc_hd__nor2_1 _19938_ (.A(_03596_),
    .B(_03597_),
    .Y(_01044_));
 sky130_fd_sc_hd__nand2_1 _19939_ (.A(\rbzero.pov.spi_counter[3] ),
    .B(_03596_),
    .Y(_03598_));
 sky130_fd_sc_hd__o211a_1 _19940_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_03596_),
    .B1(_03598_),
    .C1(_03594_),
    .X(_01045_));
 sky130_fd_sc_hd__and3_1 _19941_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[3] ),
    .C(_03596_),
    .X(_03599_));
 sky130_fd_sc_hd__a21o_1 _19942_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_03596_),
    .B1(\rbzero.pov.spi_counter[4] ),
    .X(_03600_));
 sky130_fd_sc_hd__and3b_1 _19943_ (.A_N(_03599_),
    .B(_03588_),
    .C(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__clkbuf_1 _19944_ (.A(_03601_),
    .X(_01046_));
 sky130_fd_sc_hd__and2_1 _19945_ (.A(\rbzero.pov.spi_counter[5] ),
    .B(_03599_),
    .X(_03602_));
 sky130_fd_sc_hd__o21ai_1 _19946_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_03599_),
    .B1(_03588_),
    .Y(_03603_));
 sky130_fd_sc_hd__nor2_1 _19947_ (.A(_03602_),
    .B(_03603_),
    .Y(_01047_));
 sky130_fd_sc_hd__a21boi_1 _19948_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03602_),
    .B1_N(_03594_),
    .Y(_03604_));
 sky130_fd_sc_hd__o21a_1 _19949_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03602_),
    .B1(_03604_),
    .X(_01048_));
 sky130_fd_sc_hd__and2b_1 _19950_ (.A_N(\rbzero.pov.ss_buffer[1] ),
    .B(_03586_),
    .X(_03605_));
 sky130_fd_sc_hd__buf_4 _19951_ (.A(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__buf_2 _19952_ (.A(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__or3b_1 _19953_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(\rbzero.pov.sclk_buffer[2] ),
    .C_N(\rbzero.pov.sclk_buffer[1] ),
    .X(_03608_));
 sky130_fd_sc_hd__buf_4 _19954_ (.A(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__buf_2 _19955_ (.A(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__or2_1 _19956_ (.A(\rbzero.pov.mosi ),
    .B(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__o211a_1 _19957_ (.A1(\rbzero.pov.spi_buffer[0] ),
    .A2(_03607_),
    .B1(_03611_),
    .C1(_03576_),
    .X(_01049_));
 sky130_fd_sc_hd__or2_1 _19958_ (.A(\rbzero.pov.spi_buffer[0] ),
    .B(_03610_),
    .X(_03612_));
 sky130_fd_sc_hd__o211a_1 _19959_ (.A1(\rbzero.pov.spi_buffer[1] ),
    .A2(_03607_),
    .B1(_03612_),
    .C1(_03576_),
    .X(_01050_));
 sky130_fd_sc_hd__or2_1 _19960_ (.A(\rbzero.pov.spi_buffer[1] ),
    .B(_03610_),
    .X(_03613_));
 sky130_fd_sc_hd__o211a_1 _19961_ (.A1(\rbzero.pov.spi_buffer[2] ),
    .A2(_03607_),
    .B1(_03613_),
    .C1(_03576_),
    .X(_01051_));
 sky130_fd_sc_hd__or2_1 _19962_ (.A(\rbzero.pov.spi_buffer[2] ),
    .B(_03610_),
    .X(_03614_));
 sky130_fd_sc_hd__o211a_1 _19963_ (.A1(\rbzero.pov.spi_buffer[3] ),
    .A2(_03607_),
    .B1(_03614_),
    .C1(_03576_),
    .X(_01052_));
 sky130_fd_sc_hd__or2_1 _19964_ (.A(\rbzero.pov.spi_buffer[3] ),
    .B(_03610_),
    .X(_03615_));
 sky130_fd_sc_hd__buf_2 _19965_ (.A(_02867_),
    .X(_03616_));
 sky130_fd_sc_hd__o211a_1 _19966_ (.A1(\rbzero.pov.spi_buffer[4] ),
    .A2(_03607_),
    .B1(_03615_),
    .C1(_03616_),
    .X(_01053_));
 sky130_fd_sc_hd__or2_1 _19967_ (.A(\rbzero.pov.spi_buffer[4] ),
    .B(_03610_),
    .X(_03617_));
 sky130_fd_sc_hd__o211a_1 _19968_ (.A1(\rbzero.pov.spi_buffer[5] ),
    .A2(_03607_),
    .B1(_03617_),
    .C1(_03616_),
    .X(_01054_));
 sky130_fd_sc_hd__or2_1 _19969_ (.A(\rbzero.pov.spi_buffer[5] ),
    .B(_03610_),
    .X(_03618_));
 sky130_fd_sc_hd__o211a_1 _19970_ (.A1(\rbzero.pov.spi_buffer[6] ),
    .A2(_03607_),
    .B1(_03618_),
    .C1(_03616_),
    .X(_01055_));
 sky130_fd_sc_hd__or2_1 _19971_ (.A(\rbzero.pov.spi_buffer[6] ),
    .B(_03610_),
    .X(_03619_));
 sky130_fd_sc_hd__o211a_1 _19972_ (.A1(\rbzero.pov.spi_buffer[7] ),
    .A2(_03607_),
    .B1(_03619_),
    .C1(_03616_),
    .X(_01056_));
 sky130_fd_sc_hd__or2_1 _19973_ (.A(\rbzero.pov.spi_buffer[7] ),
    .B(_03610_),
    .X(_03620_));
 sky130_fd_sc_hd__o211a_1 _19974_ (.A1(\rbzero.pov.spi_buffer[8] ),
    .A2(_03607_),
    .B1(_03620_),
    .C1(_03616_),
    .X(_01057_));
 sky130_fd_sc_hd__or2_1 _19975_ (.A(\rbzero.pov.spi_buffer[8] ),
    .B(_03610_),
    .X(_03621_));
 sky130_fd_sc_hd__o211a_1 _19976_ (.A1(\rbzero.pov.spi_buffer[9] ),
    .A2(_03607_),
    .B1(_03621_),
    .C1(_03616_),
    .X(_01058_));
 sky130_fd_sc_hd__buf_2 _19977_ (.A(_03606_),
    .X(_03622_));
 sky130_fd_sc_hd__clkbuf_2 _19978_ (.A(_03609_),
    .X(_03623_));
 sky130_fd_sc_hd__or2_1 _19979_ (.A(\rbzero.pov.spi_buffer[9] ),
    .B(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__o211a_1 _19980_ (.A1(\rbzero.pov.spi_buffer[10] ),
    .A2(_03622_),
    .B1(_03624_),
    .C1(_03616_),
    .X(_01059_));
 sky130_fd_sc_hd__or2_1 _19981_ (.A(\rbzero.pov.spi_buffer[10] ),
    .B(_03623_),
    .X(_03625_));
 sky130_fd_sc_hd__o211a_1 _19982_ (.A1(\rbzero.pov.spi_buffer[11] ),
    .A2(_03622_),
    .B1(_03625_),
    .C1(_03616_),
    .X(_01060_));
 sky130_fd_sc_hd__or2_1 _19983_ (.A(\rbzero.pov.spi_buffer[11] ),
    .B(_03623_),
    .X(_03626_));
 sky130_fd_sc_hd__o211a_1 _19984_ (.A1(\rbzero.pov.spi_buffer[12] ),
    .A2(_03622_),
    .B1(_03626_),
    .C1(_03616_),
    .X(_01061_));
 sky130_fd_sc_hd__or2_1 _19985_ (.A(\rbzero.pov.spi_buffer[12] ),
    .B(_03623_),
    .X(_03627_));
 sky130_fd_sc_hd__o211a_1 _19986_ (.A1(\rbzero.pov.spi_buffer[13] ),
    .A2(_03622_),
    .B1(_03627_),
    .C1(_03616_),
    .X(_01062_));
 sky130_fd_sc_hd__or2_1 _19987_ (.A(\rbzero.pov.spi_buffer[13] ),
    .B(_03623_),
    .X(_03628_));
 sky130_fd_sc_hd__buf_2 _19988_ (.A(_02867_),
    .X(_03629_));
 sky130_fd_sc_hd__o211a_1 _19989_ (.A1(\rbzero.pov.spi_buffer[14] ),
    .A2(_03622_),
    .B1(_03628_),
    .C1(_03629_),
    .X(_01063_));
 sky130_fd_sc_hd__or2_1 _19990_ (.A(\rbzero.pov.spi_buffer[14] ),
    .B(_03623_),
    .X(_03630_));
 sky130_fd_sc_hd__o211a_1 _19991_ (.A1(\rbzero.pov.spi_buffer[15] ),
    .A2(_03622_),
    .B1(_03630_),
    .C1(_03629_),
    .X(_01064_));
 sky130_fd_sc_hd__or2_1 _19992_ (.A(\rbzero.pov.spi_buffer[15] ),
    .B(_03623_),
    .X(_03631_));
 sky130_fd_sc_hd__o211a_1 _19993_ (.A1(\rbzero.pov.spi_buffer[16] ),
    .A2(_03622_),
    .B1(_03631_),
    .C1(_03629_),
    .X(_01065_));
 sky130_fd_sc_hd__or2_1 _19994_ (.A(\rbzero.pov.spi_buffer[16] ),
    .B(_03623_),
    .X(_03632_));
 sky130_fd_sc_hd__o211a_1 _19995_ (.A1(\rbzero.pov.spi_buffer[17] ),
    .A2(_03622_),
    .B1(_03632_),
    .C1(_03629_),
    .X(_01066_));
 sky130_fd_sc_hd__or2_1 _19996_ (.A(\rbzero.pov.spi_buffer[17] ),
    .B(_03623_),
    .X(_03633_));
 sky130_fd_sc_hd__o211a_1 _19997_ (.A1(\rbzero.pov.spi_buffer[18] ),
    .A2(_03622_),
    .B1(_03633_),
    .C1(_03629_),
    .X(_01067_));
 sky130_fd_sc_hd__or2_1 _19998_ (.A(\rbzero.pov.spi_buffer[18] ),
    .B(_03623_),
    .X(_03634_));
 sky130_fd_sc_hd__o211a_1 _19999_ (.A1(\rbzero.pov.spi_buffer[19] ),
    .A2(_03622_),
    .B1(_03634_),
    .C1(_03629_),
    .X(_01068_));
 sky130_fd_sc_hd__buf_2 _20000_ (.A(_03606_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_2 _20001_ (.A(_03609_),
    .X(_03636_));
 sky130_fd_sc_hd__or2_1 _20002_ (.A(\rbzero.pov.spi_buffer[19] ),
    .B(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__o211a_1 _20003_ (.A1(\rbzero.pov.spi_buffer[20] ),
    .A2(_03635_),
    .B1(_03637_),
    .C1(_03629_),
    .X(_01069_));
 sky130_fd_sc_hd__or2_1 _20004_ (.A(\rbzero.pov.spi_buffer[20] ),
    .B(_03636_),
    .X(_03638_));
 sky130_fd_sc_hd__o211a_1 _20005_ (.A1(\rbzero.pov.spi_buffer[21] ),
    .A2(_03635_),
    .B1(_03638_),
    .C1(_03629_),
    .X(_01070_));
 sky130_fd_sc_hd__or2_1 _20006_ (.A(\rbzero.pov.spi_buffer[21] ),
    .B(_03636_),
    .X(_03639_));
 sky130_fd_sc_hd__o211a_1 _20007_ (.A1(\rbzero.pov.spi_buffer[22] ),
    .A2(_03635_),
    .B1(_03639_),
    .C1(_03629_),
    .X(_01071_));
 sky130_fd_sc_hd__or2_1 _20008_ (.A(\rbzero.pov.spi_buffer[22] ),
    .B(_03636_),
    .X(_03640_));
 sky130_fd_sc_hd__o211a_1 _20009_ (.A1(\rbzero.pov.spi_buffer[23] ),
    .A2(_03635_),
    .B1(_03640_),
    .C1(_03629_),
    .X(_01072_));
 sky130_fd_sc_hd__or2_1 _20010_ (.A(\rbzero.pov.spi_buffer[23] ),
    .B(_03636_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_2 _20011_ (.A(_02867_),
    .X(_03642_));
 sky130_fd_sc_hd__o211a_1 _20012_ (.A1(\rbzero.pov.spi_buffer[24] ),
    .A2(_03635_),
    .B1(_03641_),
    .C1(_03642_),
    .X(_01073_));
 sky130_fd_sc_hd__or2_1 _20013_ (.A(\rbzero.pov.spi_buffer[24] ),
    .B(_03636_),
    .X(_03643_));
 sky130_fd_sc_hd__o211a_1 _20014_ (.A1(\rbzero.pov.spi_buffer[25] ),
    .A2(_03635_),
    .B1(_03643_),
    .C1(_03642_),
    .X(_01074_));
 sky130_fd_sc_hd__or2_1 _20015_ (.A(\rbzero.pov.spi_buffer[25] ),
    .B(_03636_),
    .X(_03644_));
 sky130_fd_sc_hd__o211a_1 _20016_ (.A1(\rbzero.pov.spi_buffer[26] ),
    .A2(_03635_),
    .B1(_03644_),
    .C1(_03642_),
    .X(_01075_));
 sky130_fd_sc_hd__or2_1 _20017_ (.A(\rbzero.pov.spi_buffer[26] ),
    .B(_03636_),
    .X(_03645_));
 sky130_fd_sc_hd__o211a_1 _20018_ (.A1(\rbzero.pov.spi_buffer[27] ),
    .A2(_03635_),
    .B1(_03645_),
    .C1(_03642_),
    .X(_01076_));
 sky130_fd_sc_hd__or2_1 _20019_ (.A(\rbzero.pov.spi_buffer[27] ),
    .B(_03636_),
    .X(_03646_));
 sky130_fd_sc_hd__o211a_1 _20020_ (.A1(\rbzero.pov.spi_buffer[28] ),
    .A2(_03635_),
    .B1(_03646_),
    .C1(_03642_),
    .X(_01077_));
 sky130_fd_sc_hd__or2_1 _20021_ (.A(\rbzero.pov.spi_buffer[28] ),
    .B(_03636_),
    .X(_03647_));
 sky130_fd_sc_hd__o211a_1 _20022_ (.A1(\rbzero.pov.spi_buffer[29] ),
    .A2(_03635_),
    .B1(_03647_),
    .C1(_03642_),
    .X(_01078_));
 sky130_fd_sc_hd__buf_2 _20023_ (.A(_03606_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_2 _20024_ (.A(_03609_),
    .X(_03649_));
 sky130_fd_sc_hd__or2_1 _20025_ (.A(\rbzero.pov.spi_buffer[29] ),
    .B(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__o211a_1 _20026_ (.A1(\rbzero.pov.spi_buffer[30] ),
    .A2(_03648_),
    .B1(_03650_),
    .C1(_03642_),
    .X(_01079_));
 sky130_fd_sc_hd__or2_1 _20027_ (.A(\rbzero.pov.spi_buffer[30] ),
    .B(_03649_),
    .X(_03651_));
 sky130_fd_sc_hd__o211a_1 _20028_ (.A1(\rbzero.pov.spi_buffer[31] ),
    .A2(_03648_),
    .B1(_03651_),
    .C1(_03642_),
    .X(_01080_));
 sky130_fd_sc_hd__or2_1 _20029_ (.A(\rbzero.pov.spi_buffer[31] ),
    .B(_03649_),
    .X(_03652_));
 sky130_fd_sc_hd__o211a_1 _20030_ (.A1(\rbzero.pov.spi_buffer[32] ),
    .A2(_03648_),
    .B1(_03652_),
    .C1(_03642_),
    .X(_01081_));
 sky130_fd_sc_hd__or2_1 _20031_ (.A(\rbzero.pov.spi_buffer[32] ),
    .B(_03649_),
    .X(_03653_));
 sky130_fd_sc_hd__o211a_1 _20032_ (.A1(\rbzero.pov.spi_buffer[33] ),
    .A2(_03648_),
    .B1(_03653_),
    .C1(_03642_),
    .X(_01082_));
 sky130_fd_sc_hd__or2_1 _20033_ (.A(\rbzero.pov.spi_buffer[33] ),
    .B(_03649_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_2 _20034_ (.A(_02867_),
    .X(_03655_));
 sky130_fd_sc_hd__o211a_1 _20035_ (.A1(\rbzero.pov.spi_buffer[34] ),
    .A2(_03648_),
    .B1(_03654_),
    .C1(_03655_),
    .X(_01083_));
 sky130_fd_sc_hd__or2_1 _20036_ (.A(\rbzero.pov.spi_buffer[34] ),
    .B(_03649_),
    .X(_03656_));
 sky130_fd_sc_hd__o211a_1 _20037_ (.A1(\rbzero.pov.spi_buffer[35] ),
    .A2(_03648_),
    .B1(_03656_),
    .C1(_03655_),
    .X(_01084_));
 sky130_fd_sc_hd__or2_1 _20038_ (.A(\rbzero.pov.spi_buffer[35] ),
    .B(_03649_),
    .X(_03657_));
 sky130_fd_sc_hd__o211a_1 _20039_ (.A1(\rbzero.pov.spi_buffer[36] ),
    .A2(_03648_),
    .B1(_03657_),
    .C1(_03655_),
    .X(_01085_));
 sky130_fd_sc_hd__or2_1 _20040_ (.A(\rbzero.pov.spi_buffer[36] ),
    .B(_03649_),
    .X(_03658_));
 sky130_fd_sc_hd__o211a_1 _20041_ (.A1(\rbzero.pov.spi_buffer[37] ),
    .A2(_03648_),
    .B1(_03658_),
    .C1(_03655_),
    .X(_01086_));
 sky130_fd_sc_hd__or2_1 _20042_ (.A(\rbzero.pov.spi_buffer[37] ),
    .B(_03649_),
    .X(_03659_));
 sky130_fd_sc_hd__o211a_1 _20043_ (.A1(\rbzero.pov.spi_buffer[38] ),
    .A2(_03648_),
    .B1(_03659_),
    .C1(_03655_),
    .X(_01087_));
 sky130_fd_sc_hd__or2_1 _20044_ (.A(\rbzero.pov.spi_buffer[38] ),
    .B(_03649_),
    .X(_03660_));
 sky130_fd_sc_hd__o211a_1 _20045_ (.A1(\rbzero.pov.spi_buffer[39] ),
    .A2(_03648_),
    .B1(_03660_),
    .C1(_03655_),
    .X(_01088_));
 sky130_fd_sc_hd__buf_2 _20046_ (.A(_03606_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_2 _20047_ (.A(_03609_),
    .X(_03662_));
 sky130_fd_sc_hd__or2_1 _20048_ (.A(\rbzero.pov.spi_buffer[39] ),
    .B(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__o211a_1 _20049_ (.A1(\rbzero.pov.spi_buffer[40] ),
    .A2(_03661_),
    .B1(_03663_),
    .C1(_03655_),
    .X(_01089_));
 sky130_fd_sc_hd__or2_1 _20050_ (.A(\rbzero.pov.spi_buffer[40] ),
    .B(_03662_),
    .X(_03664_));
 sky130_fd_sc_hd__o211a_1 _20051_ (.A1(\rbzero.pov.spi_buffer[41] ),
    .A2(_03661_),
    .B1(_03664_),
    .C1(_03655_),
    .X(_01090_));
 sky130_fd_sc_hd__or2_1 _20052_ (.A(\rbzero.pov.spi_buffer[41] ),
    .B(_03662_),
    .X(_03665_));
 sky130_fd_sc_hd__o211a_1 _20053_ (.A1(\rbzero.pov.spi_buffer[42] ),
    .A2(_03661_),
    .B1(_03665_),
    .C1(_03655_),
    .X(_01091_));
 sky130_fd_sc_hd__or2_1 _20054_ (.A(\rbzero.pov.spi_buffer[42] ),
    .B(_03662_),
    .X(_03666_));
 sky130_fd_sc_hd__o211a_1 _20055_ (.A1(\rbzero.pov.spi_buffer[43] ),
    .A2(_03661_),
    .B1(_03666_),
    .C1(_03655_),
    .X(_01092_));
 sky130_fd_sc_hd__or2_1 _20056_ (.A(\rbzero.pov.spi_buffer[43] ),
    .B(_03662_),
    .X(_03667_));
 sky130_fd_sc_hd__buf_2 _20057_ (.A(_02867_),
    .X(_03668_));
 sky130_fd_sc_hd__o211a_1 _20058_ (.A1(\rbzero.pov.spi_buffer[44] ),
    .A2(_03661_),
    .B1(_03667_),
    .C1(_03668_),
    .X(_01093_));
 sky130_fd_sc_hd__or2_1 _20059_ (.A(\rbzero.pov.spi_buffer[44] ),
    .B(_03662_),
    .X(_03669_));
 sky130_fd_sc_hd__o211a_1 _20060_ (.A1(\rbzero.pov.spi_buffer[45] ),
    .A2(_03661_),
    .B1(_03669_),
    .C1(_03668_),
    .X(_01094_));
 sky130_fd_sc_hd__or2_1 _20061_ (.A(\rbzero.pov.spi_buffer[45] ),
    .B(_03662_),
    .X(_03670_));
 sky130_fd_sc_hd__o211a_1 _20062_ (.A1(\rbzero.pov.spi_buffer[46] ),
    .A2(_03661_),
    .B1(_03670_),
    .C1(_03668_),
    .X(_01095_));
 sky130_fd_sc_hd__or2_1 _20063_ (.A(\rbzero.pov.spi_buffer[46] ),
    .B(_03662_),
    .X(_03671_));
 sky130_fd_sc_hd__o211a_1 _20064_ (.A1(\rbzero.pov.spi_buffer[47] ),
    .A2(_03661_),
    .B1(_03671_),
    .C1(_03668_),
    .X(_01096_));
 sky130_fd_sc_hd__or2_1 _20065_ (.A(\rbzero.pov.spi_buffer[47] ),
    .B(_03662_),
    .X(_03672_));
 sky130_fd_sc_hd__o211a_1 _20066_ (.A1(\rbzero.pov.spi_buffer[48] ),
    .A2(_03661_),
    .B1(_03672_),
    .C1(_03668_),
    .X(_01097_));
 sky130_fd_sc_hd__or2_1 _20067_ (.A(\rbzero.pov.spi_buffer[48] ),
    .B(_03662_),
    .X(_03673_));
 sky130_fd_sc_hd__o211a_1 _20068_ (.A1(\rbzero.pov.spi_buffer[49] ),
    .A2(_03661_),
    .B1(_03673_),
    .C1(_03668_),
    .X(_01098_));
 sky130_fd_sc_hd__buf_2 _20069_ (.A(_03606_),
    .X(_03674_));
 sky130_fd_sc_hd__clkbuf_2 _20070_ (.A(_03609_),
    .X(_03675_));
 sky130_fd_sc_hd__or2_1 _20071_ (.A(\rbzero.pov.spi_buffer[49] ),
    .B(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__o211a_1 _20072_ (.A1(\rbzero.pov.spi_buffer[50] ),
    .A2(_03674_),
    .B1(_03676_),
    .C1(_03668_),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _20073_ (.A(\rbzero.pov.spi_buffer[50] ),
    .B(_03675_),
    .X(_03677_));
 sky130_fd_sc_hd__o211a_1 _20074_ (.A1(\rbzero.pov.spi_buffer[51] ),
    .A2(_03674_),
    .B1(_03677_),
    .C1(_03668_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_1 _20075_ (.A(\rbzero.pov.spi_buffer[51] ),
    .B(_03675_),
    .X(_03678_));
 sky130_fd_sc_hd__o211a_1 _20076_ (.A1(\rbzero.pov.spi_buffer[52] ),
    .A2(_03674_),
    .B1(_03678_),
    .C1(_03668_),
    .X(_01101_));
 sky130_fd_sc_hd__or2_1 _20077_ (.A(\rbzero.pov.spi_buffer[52] ),
    .B(_03675_),
    .X(_03679_));
 sky130_fd_sc_hd__o211a_1 _20078_ (.A1(\rbzero.pov.spi_buffer[53] ),
    .A2(_03674_),
    .B1(_03679_),
    .C1(_03668_),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _20079_ (.A(\rbzero.pov.spi_buffer[53] ),
    .B(_03675_),
    .X(_03680_));
 sky130_fd_sc_hd__buf_2 _20080_ (.A(_02867_),
    .X(_03681_));
 sky130_fd_sc_hd__o211a_1 _20081_ (.A1(\rbzero.pov.spi_buffer[54] ),
    .A2(_03674_),
    .B1(_03680_),
    .C1(_03681_),
    .X(_01103_));
 sky130_fd_sc_hd__or2_1 _20082_ (.A(\rbzero.pov.spi_buffer[54] ),
    .B(_03675_),
    .X(_03682_));
 sky130_fd_sc_hd__o211a_1 _20083_ (.A1(\rbzero.pov.spi_buffer[55] ),
    .A2(_03674_),
    .B1(_03682_),
    .C1(_03681_),
    .X(_01104_));
 sky130_fd_sc_hd__or2_1 _20084_ (.A(\rbzero.pov.spi_buffer[55] ),
    .B(_03675_),
    .X(_03683_));
 sky130_fd_sc_hd__o211a_1 _20085_ (.A1(\rbzero.pov.spi_buffer[56] ),
    .A2(_03674_),
    .B1(_03683_),
    .C1(_03681_),
    .X(_01105_));
 sky130_fd_sc_hd__or2_1 _20086_ (.A(\rbzero.pov.spi_buffer[56] ),
    .B(_03675_),
    .X(_03684_));
 sky130_fd_sc_hd__o211a_1 _20087_ (.A1(\rbzero.pov.spi_buffer[57] ),
    .A2(_03674_),
    .B1(_03684_),
    .C1(_03681_),
    .X(_01106_));
 sky130_fd_sc_hd__or2_1 _20088_ (.A(\rbzero.pov.spi_buffer[57] ),
    .B(_03675_),
    .X(_03685_));
 sky130_fd_sc_hd__o211a_1 _20089_ (.A1(\rbzero.pov.spi_buffer[58] ),
    .A2(_03674_),
    .B1(_03685_),
    .C1(_03681_),
    .X(_01107_));
 sky130_fd_sc_hd__or2_1 _20090_ (.A(\rbzero.pov.spi_buffer[58] ),
    .B(_03675_),
    .X(_03686_));
 sky130_fd_sc_hd__o211a_1 _20091_ (.A1(\rbzero.pov.spi_buffer[59] ),
    .A2(_03674_),
    .B1(_03686_),
    .C1(_03681_),
    .X(_01108_));
 sky130_fd_sc_hd__buf_2 _20092_ (.A(_03605_),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_2 _20093_ (.A(_03608_),
    .X(_03688_));
 sky130_fd_sc_hd__or2_1 _20094_ (.A(\rbzero.pov.spi_buffer[59] ),
    .B(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__o211a_1 _20095_ (.A1(\rbzero.pov.spi_buffer[60] ),
    .A2(_03687_),
    .B1(_03689_),
    .C1(_03681_),
    .X(_01109_));
 sky130_fd_sc_hd__or2_1 _20096_ (.A(\rbzero.pov.spi_buffer[60] ),
    .B(_03688_),
    .X(_03690_));
 sky130_fd_sc_hd__o211a_1 _20097_ (.A1(\rbzero.pov.spi_buffer[61] ),
    .A2(_03687_),
    .B1(_03690_),
    .C1(_03681_),
    .X(_01110_));
 sky130_fd_sc_hd__or2_1 _20098_ (.A(\rbzero.pov.spi_buffer[61] ),
    .B(_03688_),
    .X(_03691_));
 sky130_fd_sc_hd__o211a_1 _20099_ (.A1(\rbzero.pov.spi_buffer[62] ),
    .A2(_03687_),
    .B1(_03691_),
    .C1(_03681_),
    .X(_01111_));
 sky130_fd_sc_hd__or2_1 _20100_ (.A(\rbzero.pov.spi_buffer[62] ),
    .B(_03688_),
    .X(_03692_));
 sky130_fd_sc_hd__o211a_1 _20101_ (.A1(\rbzero.pov.spi_buffer[63] ),
    .A2(_03687_),
    .B1(_03692_),
    .C1(_03681_),
    .X(_01112_));
 sky130_fd_sc_hd__or2_1 _20102_ (.A(\rbzero.pov.spi_buffer[63] ),
    .B(_03688_),
    .X(_03693_));
 sky130_fd_sc_hd__buf_2 _20103_ (.A(_02867_),
    .X(_03694_));
 sky130_fd_sc_hd__o211a_1 _20104_ (.A1(\rbzero.pov.spi_buffer[64] ),
    .A2(_03687_),
    .B1(_03693_),
    .C1(_03694_),
    .X(_01113_));
 sky130_fd_sc_hd__or2_1 _20105_ (.A(\rbzero.pov.spi_buffer[64] ),
    .B(_03688_),
    .X(_03695_));
 sky130_fd_sc_hd__o211a_1 _20106_ (.A1(\rbzero.pov.spi_buffer[65] ),
    .A2(_03687_),
    .B1(_03695_),
    .C1(_03694_),
    .X(_01114_));
 sky130_fd_sc_hd__or2_1 _20107_ (.A(\rbzero.pov.spi_buffer[65] ),
    .B(_03688_),
    .X(_03696_));
 sky130_fd_sc_hd__o211a_1 _20108_ (.A1(\rbzero.pov.spi_buffer[66] ),
    .A2(_03687_),
    .B1(_03696_),
    .C1(_03694_),
    .X(_01115_));
 sky130_fd_sc_hd__or2_1 _20109_ (.A(\rbzero.pov.spi_buffer[66] ),
    .B(_03688_),
    .X(_03697_));
 sky130_fd_sc_hd__o211a_1 _20110_ (.A1(\rbzero.pov.spi_buffer[67] ),
    .A2(_03687_),
    .B1(_03697_),
    .C1(_03694_),
    .X(_01116_));
 sky130_fd_sc_hd__or2_1 _20111_ (.A(\rbzero.pov.spi_buffer[67] ),
    .B(_03688_),
    .X(_03698_));
 sky130_fd_sc_hd__o211a_1 _20112_ (.A1(\rbzero.pov.spi_buffer[68] ),
    .A2(_03687_),
    .B1(_03698_),
    .C1(_03694_),
    .X(_01117_));
 sky130_fd_sc_hd__or2_1 _20113_ (.A(\rbzero.pov.spi_buffer[68] ),
    .B(_03688_),
    .X(_03699_));
 sky130_fd_sc_hd__o211a_1 _20114_ (.A1(\rbzero.pov.spi_buffer[69] ),
    .A2(_03687_),
    .B1(_03699_),
    .C1(_03694_),
    .X(_01118_));
 sky130_fd_sc_hd__or2_1 _20115_ (.A(\rbzero.pov.spi_buffer[69] ),
    .B(_03609_),
    .X(_03700_));
 sky130_fd_sc_hd__o211a_1 _20116_ (.A1(\rbzero.pov.spi_buffer[70] ),
    .A2(_03606_),
    .B1(_03700_),
    .C1(_03694_),
    .X(_01119_));
 sky130_fd_sc_hd__or2_1 _20117_ (.A(\rbzero.pov.spi_buffer[70] ),
    .B(_03609_),
    .X(_03701_));
 sky130_fd_sc_hd__o211a_1 _20118_ (.A1(\rbzero.pov.spi_buffer[71] ),
    .A2(_03606_),
    .B1(_03701_),
    .C1(_03694_),
    .X(_01120_));
 sky130_fd_sc_hd__or2_1 _20119_ (.A(\rbzero.pov.spi_buffer[71] ),
    .B(_03609_),
    .X(_03702_));
 sky130_fd_sc_hd__o211a_1 _20120_ (.A1(\rbzero.pov.spi_buffer[72] ),
    .A2(_03606_),
    .B1(_03702_),
    .C1(_03694_),
    .X(_01121_));
 sky130_fd_sc_hd__or2_1 _20121_ (.A(\rbzero.pov.spi_buffer[72] ),
    .B(_03609_),
    .X(_03703_));
 sky130_fd_sc_hd__o211a_1 _20122_ (.A1(\rbzero.pov.spi_buffer[73] ),
    .A2(_03606_),
    .B1(_03703_),
    .C1(_03694_),
    .X(_01122_));
 sky130_fd_sc_hd__buf_1 _20123_ (.A(clknet_1_1__leaf__04767_),
    .X(_03704_));
 sky130_fd_sc_hd__buf_1 _20124_ (.A(clknet_1_0__leaf__03704_),
    .X(_03705_));
 sky130_fd_sc_hd__inv_2 _20126__29 (.A(clknet_1_1__leaf__03705_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _20127__30 (.A(clknet_1_1__leaf__03705_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _20128__31 (.A(clknet_1_1__leaf__03705_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _20129__32 (.A(clknet_1_1__leaf__03705_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _20130__33 (.A(clknet_1_0__leaf__03705_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _20131__34 (.A(clknet_1_0__leaf__03705_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _20132__35 (.A(clknet_1_0__leaf__03705_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _20133__36 (.A(clknet_1_0__leaf__03705_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _20134__37 (.A(clknet_1_0__leaf__03705_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _20136__38 (.A(clknet_1_0__leaf__03706_),
    .Y(net163));
 sky130_fd_sc_hd__buf_1 _20135_ (.A(clknet_1_1__leaf__03704_),
    .X(_03706_));
 sky130_fd_sc_hd__inv_2 _20137__39 (.A(clknet_1_0__leaf__03706_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _20138__40 (.A(clknet_1_0__leaf__03706_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _20139__41 (.A(clknet_1_1__leaf__03706_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _20140__42 (.A(clknet_1_0__leaf__03706_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _20141__43 (.A(clknet_1_1__leaf__03706_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _20142__44 (.A(clknet_1_1__leaf__03706_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _20143__45 (.A(clknet_1_1__leaf__03706_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _20144__46 (.A(clknet_1_1__leaf__03706_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _20145__47 (.A(clknet_1_1__leaf__03706_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _20147__48 (.A(clknet_1_1__leaf__03707_),
    .Y(net173));
 sky130_fd_sc_hd__buf_1 _20146_ (.A(clknet_1_1__leaf__03704_),
    .X(_03707_));
 sky130_fd_sc_hd__inv_2 _20148__49 (.A(clknet_1_1__leaf__03707_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _20149__50 (.A(clknet_1_1__leaf__03707_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _20150__51 (.A(clknet_1_1__leaf__03707_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _20151__52 (.A(clknet_1_1__leaf__03707_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _20152__53 (.A(clknet_1_1__leaf__03707_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _20153__54 (.A(clknet_1_0__leaf__03707_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _20154__55 (.A(clknet_1_0__leaf__03707_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _20155__56 (.A(clknet_1_0__leaf__03707_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _20156__57 (.A(clknet_1_0__leaf__03707_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _20158__58 (.A(clknet_1_1__leaf__03708_),
    .Y(net183));
 sky130_fd_sc_hd__buf_1 _20157_ (.A(clknet_1_0__leaf__03704_),
    .X(_03708_));
 sky130_fd_sc_hd__inv_2 _20159__59 (.A(clknet_1_1__leaf__03708_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _20160__60 (.A(clknet_1_1__leaf__03708_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _20161__61 (.A(clknet_1_1__leaf__03708_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _20162__62 (.A(clknet_1_1__leaf__03708_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _20163__63 (.A(clknet_1_0__leaf__03708_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _20164__64 (.A(clknet_1_0__leaf__03708_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _20165__65 (.A(clknet_1_0__leaf__03708_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _20166__66 (.A(clknet_1_0__leaf__03708_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _20167__67 (.A(clknet_1_0__leaf__03708_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _20169__68 (.A(clknet_1_0__leaf__03709_),
    .Y(net193));
 sky130_fd_sc_hd__buf_1 _20168_ (.A(clknet_1_0__leaf__03704_),
    .X(_03709_));
 sky130_fd_sc_hd__inv_2 _20170__69 (.A(clknet_1_0__leaf__03709_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _20171__70 (.A(clknet_1_0__leaf__03709_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _20172__71 (.A(clknet_1_0__leaf__03709_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _20173__72 (.A(clknet_1_0__leaf__03709_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _20174__73 (.A(clknet_1_1__leaf__03709_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _20175__74 (.A(clknet_1_1__leaf__03709_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _20176__75 (.A(clknet_1_1__leaf__03709_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _20177__76 (.A(clknet_1_1__leaf__03709_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _20178__77 (.A(clknet_1_1__leaf__03709_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _20180__78 (.A(clknet_1_1__leaf__03710_),
    .Y(net203));
 sky130_fd_sc_hd__buf_1 _20179_ (.A(clknet_1_0__leaf__03704_),
    .X(_03710_));
 sky130_fd_sc_hd__inv_2 _20181__79 (.A(clknet_1_1__leaf__03710_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _20182__80 (.A(clknet_1_1__leaf__03710_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _20183__81 (.A(clknet_1_1__leaf__03710_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _20184__82 (.A(clknet_1_0__leaf__03710_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _20185__83 (.A(clknet_1_0__leaf__03710_),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _20186__84 (.A(clknet_1_0__leaf__03710_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _20187__85 (.A(clknet_1_0__leaf__03710_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _20188__86 (.A(clknet_1_0__leaf__03710_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _20189__87 (.A(clknet_1_0__leaf__03710_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _20192__88 (.A(clknet_1_0__leaf__03712_),
    .Y(net213));
 sky130_fd_sc_hd__buf_1 _20190_ (.A(clknet_1_1__leaf__04767_),
    .X(_03711_));
 sky130_fd_sc_hd__buf_1 _20191_ (.A(clknet_1_1__leaf__03711_),
    .X(_03712_));
 sky130_fd_sc_hd__inv_2 _20193__89 (.A(clknet_1_0__leaf__03712_),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _20194__90 (.A(clknet_1_0__leaf__03712_),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _20195__91 (.A(clknet_1_0__leaf__03712_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _20486__92 (.A(clknet_1_1__leaf__03712_),
    .Y(net217));
 sky130_fd_sc_hd__buf_4 _20196_ (.A(\rbzero.pov.spi_done ),
    .X(_03713_));
 sky130_fd_sc_hd__o211a_1 _20197_ (.A1(_03713_),
    .A2(\rbzero.pov.ready ),
    .B1(_02883_),
    .C1(_03430_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _20198_ (.A0(\rbzero.pov.ready_buffer[0] ),
    .A1(\rbzero.pov.spi_buffer[0] ),
    .S(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__and2_1 _20199_ (.A(_08249_),
    .B(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_1 _20200_ (.A(_03715_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _20201_ (.A0(\rbzero.pov.ready_buffer[1] ),
    .A1(\rbzero.pov.spi_buffer[1] ),
    .S(_03713_),
    .X(_03716_));
 sky130_fd_sc_hd__and2_1 _20202_ (.A(_08249_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_1 _20203_ (.A(_03717_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _20204_ (.A0(\rbzero.pov.ready_buffer[2] ),
    .A1(\rbzero.pov.spi_buffer[2] ),
    .S(_03713_),
    .X(_03718_));
 sky130_fd_sc_hd__and2_1 _20205_ (.A(_08249_),
    .B(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_1 _20206_ (.A(_03719_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _20207_ (.A0(\rbzero.pov.ready_buffer[3] ),
    .A1(\rbzero.pov.spi_buffer[3] ),
    .S(_03713_),
    .X(_03720_));
 sky130_fd_sc_hd__and2_1 _20208_ (.A(_08249_),
    .B(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_1 _20209_ (.A(_03721_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _20210_ (.A0(\rbzero.pov.ready_buffer[4] ),
    .A1(\rbzero.pov.spi_buffer[4] ),
    .S(_03713_),
    .X(_03722_));
 sky130_fd_sc_hd__and2_1 _20211_ (.A(_08249_),
    .B(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_1 _20212_ (.A(_03723_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _20213_ (.A0(\rbzero.pov.ready_buffer[5] ),
    .A1(\rbzero.pov.spi_buffer[5] ),
    .S(_03713_),
    .X(_03724_));
 sky130_fd_sc_hd__and2_1 _20214_ (.A(_08249_),
    .B(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_1 _20215_ (.A(_03725_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _20216_ (.A0(\rbzero.pov.ready_buffer[6] ),
    .A1(\rbzero.pov.spi_buffer[6] ),
    .S(_03713_),
    .X(_03726_));
 sky130_fd_sc_hd__and2_1 _20217_ (.A(_08249_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _20218_ (.A(_03727_),
    .X(_01194_));
 sky130_fd_sc_hd__clkbuf_2 _20219_ (.A(_08245_),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_1 _20220_ (.A0(\rbzero.pov.ready_buffer[7] ),
    .A1(\rbzero.pov.spi_buffer[7] ),
    .S(_03713_),
    .X(_03729_));
 sky130_fd_sc_hd__and2_1 _20221_ (.A(_03728_),
    .B(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__clkbuf_1 _20222_ (.A(_03730_),
    .X(_01195_));
 sky130_fd_sc_hd__buf_4 _20223_ (.A(\rbzero.pov.spi_done ),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_4 _20224_ (.A(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__mux2_1 _20225_ (.A0(\rbzero.pov.ready_buffer[8] ),
    .A1(\rbzero.pov.spi_buffer[8] ),
    .S(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__and2_1 _20226_ (.A(_03728_),
    .B(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__clkbuf_1 _20227_ (.A(_03734_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _20228_ (.A0(\rbzero.pov.ready_buffer[9] ),
    .A1(\rbzero.pov.spi_buffer[9] ),
    .S(_03732_),
    .X(_03735_));
 sky130_fd_sc_hd__and2_1 _20229_ (.A(_03728_),
    .B(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_1 _20230_ (.A(_03736_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _20231_ (.A0(\rbzero.pov.ready_buffer[10] ),
    .A1(\rbzero.pov.spi_buffer[10] ),
    .S(_03732_),
    .X(_03737_));
 sky130_fd_sc_hd__and2_1 _20232_ (.A(_03728_),
    .B(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__clkbuf_1 _20233_ (.A(_03738_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _20234_ (.A0(\rbzero.pov.ready_buffer[11] ),
    .A1(\rbzero.pov.spi_buffer[11] ),
    .S(_03732_),
    .X(_03739_));
 sky130_fd_sc_hd__and2_1 _20235_ (.A(_03728_),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__clkbuf_1 _20236_ (.A(_03740_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _20237_ (.A0(\rbzero.pov.ready_buffer[12] ),
    .A1(\rbzero.pov.spi_buffer[12] ),
    .S(_03732_),
    .X(_03741_));
 sky130_fd_sc_hd__and2_1 _20238_ (.A(_03728_),
    .B(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _20239_ (.A(_03742_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _20240_ (.A0(\rbzero.pov.ready_buffer[13] ),
    .A1(\rbzero.pov.spi_buffer[13] ),
    .S(_03732_),
    .X(_03743_));
 sky130_fd_sc_hd__and2_1 _20241_ (.A(_03728_),
    .B(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_1 _20242_ (.A(_03744_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _20243_ (.A0(\rbzero.pov.ready_buffer[14] ),
    .A1(\rbzero.pov.spi_buffer[14] ),
    .S(_03732_),
    .X(_03745_));
 sky130_fd_sc_hd__and2_1 _20244_ (.A(_03728_),
    .B(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _20245_ (.A(_03746_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _20246_ (.A0(\rbzero.pov.ready_buffer[15] ),
    .A1(\rbzero.pov.spi_buffer[15] ),
    .S(_03732_),
    .X(_03747_));
 sky130_fd_sc_hd__and2_1 _20247_ (.A(_03728_),
    .B(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__clkbuf_1 _20248_ (.A(_03748_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _20249_ (.A0(\rbzero.pov.ready_buffer[16] ),
    .A1(\rbzero.pov.spi_buffer[16] ),
    .S(_03732_),
    .X(_03749_));
 sky130_fd_sc_hd__and2_1 _20250_ (.A(_03728_),
    .B(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__clkbuf_1 _20251_ (.A(_03750_),
    .X(_01204_));
 sky130_fd_sc_hd__clkbuf_2 _20252_ (.A(_08245_),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_1 _20253_ (.A0(\rbzero.pov.ready_buffer[17] ),
    .A1(\rbzero.pov.spi_buffer[17] ),
    .S(_03732_),
    .X(_03752_));
 sky130_fd_sc_hd__and2_1 _20254_ (.A(_03751_),
    .B(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__clkbuf_1 _20255_ (.A(_03753_),
    .X(_01205_));
 sky130_fd_sc_hd__clkbuf_4 _20256_ (.A(_03731_),
    .X(_03754_));
 sky130_fd_sc_hd__mux2_1 _20257_ (.A0(\rbzero.pov.ready_buffer[18] ),
    .A1(\rbzero.pov.spi_buffer[18] ),
    .S(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__and2_1 _20258_ (.A(_03751_),
    .B(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _20259_ (.A(_03756_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _20260_ (.A0(\rbzero.pov.ready_buffer[19] ),
    .A1(\rbzero.pov.spi_buffer[19] ),
    .S(_03754_),
    .X(_03757_));
 sky130_fd_sc_hd__and2_1 _20261_ (.A(_03751_),
    .B(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _20262_ (.A(_03758_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _20263_ (.A0(\rbzero.pov.ready_buffer[20] ),
    .A1(\rbzero.pov.spi_buffer[20] ),
    .S(_03754_),
    .X(_03759_));
 sky130_fd_sc_hd__and2_1 _20264_ (.A(_03751_),
    .B(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_1 _20265_ (.A(_03760_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _20266_ (.A0(\rbzero.pov.ready_buffer[21] ),
    .A1(\rbzero.pov.spi_buffer[21] ),
    .S(_03754_),
    .X(_03761_));
 sky130_fd_sc_hd__and2_1 _20267_ (.A(_03751_),
    .B(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _20268_ (.A(_03762_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _20269_ (.A0(\rbzero.pov.ready_buffer[22] ),
    .A1(\rbzero.pov.spi_buffer[22] ),
    .S(_03754_),
    .X(_03763_));
 sky130_fd_sc_hd__and2_1 _20270_ (.A(_03751_),
    .B(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _20271_ (.A(_03764_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _20272_ (.A0(\rbzero.pov.ready_buffer[23] ),
    .A1(\rbzero.pov.spi_buffer[23] ),
    .S(_03754_),
    .X(_03765_));
 sky130_fd_sc_hd__and2_1 _20273_ (.A(_03751_),
    .B(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _20274_ (.A(_03766_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _20275_ (.A0(\rbzero.pov.ready_buffer[24] ),
    .A1(\rbzero.pov.spi_buffer[24] ),
    .S(_03754_),
    .X(_03767_));
 sky130_fd_sc_hd__and2_1 _20276_ (.A(_03751_),
    .B(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_1 _20277_ (.A(_03768_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _20278_ (.A0(\rbzero.pov.ready_buffer[25] ),
    .A1(\rbzero.pov.spi_buffer[25] ),
    .S(_03754_),
    .X(_03769_));
 sky130_fd_sc_hd__and2_1 _20279_ (.A(_03751_),
    .B(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _20280_ (.A(_03770_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _20281_ (.A0(\rbzero.pov.ready_buffer[26] ),
    .A1(\rbzero.pov.spi_buffer[26] ),
    .S(_03754_),
    .X(_03771_));
 sky130_fd_sc_hd__and2_1 _20282_ (.A(_03751_),
    .B(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _20283_ (.A(_03772_),
    .X(_01214_));
 sky130_fd_sc_hd__clkbuf_2 _20284_ (.A(_08245_),
    .X(_03773_));
 sky130_fd_sc_hd__mux2_1 _20285_ (.A0(\rbzero.pov.ready_buffer[27] ),
    .A1(\rbzero.pov.spi_buffer[27] ),
    .S(_03754_),
    .X(_03774_));
 sky130_fd_sc_hd__and2_1 _20286_ (.A(_03773_),
    .B(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__clkbuf_1 _20287_ (.A(_03775_),
    .X(_01215_));
 sky130_fd_sc_hd__clkbuf_4 _20288_ (.A(_03731_),
    .X(_03776_));
 sky130_fd_sc_hd__mux2_1 _20289_ (.A0(\rbzero.pov.ready_buffer[28] ),
    .A1(\rbzero.pov.spi_buffer[28] ),
    .S(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__and2_1 _20290_ (.A(_03773_),
    .B(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__clkbuf_1 _20291_ (.A(_03778_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _20292_ (.A0(\rbzero.pov.ready_buffer[29] ),
    .A1(\rbzero.pov.spi_buffer[29] ),
    .S(_03776_),
    .X(_03779_));
 sky130_fd_sc_hd__and2_1 _20293_ (.A(_03773_),
    .B(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_1 _20294_ (.A(_03780_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _20295_ (.A0(\rbzero.pov.ready_buffer[30] ),
    .A1(\rbzero.pov.spi_buffer[30] ),
    .S(_03776_),
    .X(_03781_));
 sky130_fd_sc_hd__and2_1 _20296_ (.A(_03773_),
    .B(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_1 _20297_ (.A(_03782_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _20298_ (.A0(\rbzero.pov.ready_buffer[31] ),
    .A1(\rbzero.pov.spi_buffer[31] ),
    .S(_03776_),
    .X(_03783_));
 sky130_fd_sc_hd__and2_1 _20299_ (.A(_03773_),
    .B(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__clkbuf_1 _20300_ (.A(_03784_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _20301_ (.A0(\rbzero.pov.ready_buffer[32] ),
    .A1(\rbzero.pov.spi_buffer[32] ),
    .S(_03776_),
    .X(_03785_));
 sky130_fd_sc_hd__and2_1 _20302_ (.A(_03773_),
    .B(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__clkbuf_1 _20303_ (.A(_03786_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _20304_ (.A0(\rbzero.pov.ready_buffer[33] ),
    .A1(\rbzero.pov.spi_buffer[33] ),
    .S(_03776_),
    .X(_03787_));
 sky130_fd_sc_hd__and2_1 _20305_ (.A(_03773_),
    .B(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__clkbuf_1 _20306_ (.A(_03788_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _20307_ (.A0(\rbzero.pov.ready_buffer[34] ),
    .A1(\rbzero.pov.spi_buffer[34] ),
    .S(_03776_),
    .X(_03789_));
 sky130_fd_sc_hd__and2_1 _20308_ (.A(_03773_),
    .B(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__clkbuf_1 _20309_ (.A(_03790_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _20310_ (.A0(\rbzero.pov.ready_buffer[35] ),
    .A1(\rbzero.pov.spi_buffer[35] ),
    .S(_03776_),
    .X(_03791_));
 sky130_fd_sc_hd__and2_1 _20311_ (.A(_03773_),
    .B(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__clkbuf_1 _20312_ (.A(_03792_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _20313_ (.A0(\rbzero.pov.ready_buffer[36] ),
    .A1(\rbzero.pov.spi_buffer[36] ),
    .S(_03776_),
    .X(_03793_));
 sky130_fd_sc_hd__and2_1 _20314_ (.A(_03773_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__clkbuf_1 _20315_ (.A(_03794_),
    .X(_01224_));
 sky130_fd_sc_hd__clkbuf_2 _20316_ (.A(_08245_),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _20317_ (.A0(\rbzero.pov.ready_buffer[37] ),
    .A1(\rbzero.pov.spi_buffer[37] ),
    .S(_03776_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _20318_ (.A(_03795_),
    .B(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__clkbuf_1 _20319_ (.A(_03797_),
    .X(_01225_));
 sky130_fd_sc_hd__clkbuf_4 _20320_ (.A(_03731_),
    .X(_03798_));
 sky130_fd_sc_hd__mux2_1 _20321_ (.A0(\rbzero.pov.ready_buffer[38] ),
    .A1(\rbzero.pov.spi_buffer[38] ),
    .S(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_1 _20322_ (.A(_03795_),
    .B(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__clkbuf_1 _20323_ (.A(_03800_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _20324_ (.A0(\rbzero.pov.ready_buffer[39] ),
    .A1(\rbzero.pov.spi_buffer[39] ),
    .S(_03798_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_1 _20325_ (.A(_03795_),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__clkbuf_1 _20326_ (.A(_03802_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _20327_ (.A0(\rbzero.pov.ready_buffer[40] ),
    .A1(\rbzero.pov.spi_buffer[40] ),
    .S(_03798_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_1 _20328_ (.A(_03795_),
    .B(_03803_),
    .X(_03804_));
 sky130_fd_sc_hd__clkbuf_1 _20329_ (.A(_03804_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _20330_ (.A0(\rbzero.pov.ready_buffer[41] ),
    .A1(\rbzero.pov.spi_buffer[41] ),
    .S(_03798_),
    .X(_03805_));
 sky130_fd_sc_hd__and2_1 _20331_ (.A(_03795_),
    .B(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_1 _20332_ (.A(_03806_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _20333_ (.A0(\rbzero.pov.ready_buffer[42] ),
    .A1(\rbzero.pov.spi_buffer[42] ),
    .S(_03798_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_1 _20334_ (.A(_03795_),
    .B(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__clkbuf_1 _20335_ (.A(_03808_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _20336_ (.A0(\rbzero.pov.ready_buffer[43] ),
    .A1(\rbzero.pov.spi_buffer[43] ),
    .S(_03798_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_1 _20337_ (.A(_03795_),
    .B(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _20338_ (.A(_03810_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _20339_ (.A0(\rbzero.pov.ready_buffer[44] ),
    .A1(\rbzero.pov.spi_buffer[44] ),
    .S(_03798_),
    .X(_03811_));
 sky130_fd_sc_hd__and2_1 _20340_ (.A(_03795_),
    .B(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_1 _20341_ (.A(_03812_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _20342_ (.A0(\rbzero.pov.ready_buffer[45] ),
    .A1(\rbzero.pov.spi_buffer[45] ),
    .S(_03798_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_1 _20343_ (.A(_03795_),
    .B(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_1 _20344_ (.A(_03814_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _20345_ (.A0(\rbzero.pov.ready_buffer[46] ),
    .A1(\rbzero.pov.spi_buffer[46] ),
    .S(_03798_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _20346_ (.A(_03795_),
    .B(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _20347_ (.A(_03816_),
    .X(_01234_));
 sky130_fd_sc_hd__clkbuf_2 _20348_ (.A(_08245_),
    .X(_03817_));
 sky130_fd_sc_hd__mux2_1 _20349_ (.A0(\rbzero.pov.ready_buffer[47] ),
    .A1(\rbzero.pov.spi_buffer[47] ),
    .S(_03798_),
    .X(_03818_));
 sky130_fd_sc_hd__and2_1 _20350_ (.A(_03817_),
    .B(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_1 _20351_ (.A(_03819_),
    .X(_01235_));
 sky130_fd_sc_hd__clkbuf_4 _20352_ (.A(\rbzero.pov.spi_done ),
    .X(_03820_));
 sky130_fd_sc_hd__mux2_1 _20353_ (.A0(\rbzero.pov.ready_buffer[48] ),
    .A1(\rbzero.pov.spi_buffer[48] ),
    .S(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_1 _20354_ (.A(_03817_),
    .B(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _20355_ (.A(_03822_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _20356_ (.A0(\rbzero.pov.ready_buffer[49] ),
    .A1(\rbzero.pov.spi_buffer[49] ),
    .S(_03820_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_1 _20357_ (.A(_03817_),
    .B(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _20358_ (.A(_03824_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _20359_ (.A0(\rbzero.pov.ready_buffer[50] ),
    .A1(\rbzero.pov.spi_buffer[50] ),
    .S(_03820_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_1 _20360_ (.A(_03817_),
    .B(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__clkbuf_1 _20361_ (.A(_03826_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _20362_ (.A0(\rbzero.pov.ready_buffer[51] ),
    .A1(\rbzero.pov.spi_buffer[51] ),
    .S(_03820_),
    .X(_03827_));
 sky130_fd_sc_hd__and2_1 _20363_ (.A(_03817_),
    .B(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_1 _20364_ (.A(_03828_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _20365_ (.A0(\rbzero.pov.ready_buffer[52] ),
    .A1(\rbzero.pov.spi_buffer[52] ),
    .S(_03820_),
    .X(_03829_));
 sky130_fd_sc_hd__and2_1 _20366_ (.A(_03817_),
    .B(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__clkbuf_1 _20367_ (.A(_03830_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _20368_ (.A0(\rbzero.pov.ready_buffer[53] ),
    .A1(\rbzero.pov.spi_buffer[53] ),
    .S(_03820_),
    .X(_03831_));
 sky130_fd_sc_hd__and2_1 _20369_ (.A(_03817_),
    .B(_03831_),
    .X(_03832_));
 sky130_fd_sc_hd__clkbuf_1 _20370_ (.A(_03832_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _20371_ (.A0(\rbzero.pov.ready_buffer[54] ),
    .A1(\rbzero.pov.spi_buffer[54] ),
    .S(_03820_),
    .X(_03833_));
 sky130_fd_sc_hd__and2_1 _20372_ (.A(_03817_),
    .B(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _20373_ (.A(_03834_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _20374_ (.A0(\rbzero.pov.ready_buffer[55] ),
    .A1(\rbzero.pov.spi_buffer[55] ),
    .S(_03820_),
    .X(_03835_));
 sky130_fd_sc_hd__and2_1 _20375_ (.A(_03817_),
    .B(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__clkbuf_1 _20376_ (.A(_03836_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _20377_ (.A0(\rbzero.pov.ready_buffer[56] ),
    .A1(\rbzero.pov.spi_buffer[56] ),
    .S(_03820_),
    .X(_03837_));
 sky130_fd_sc_hd__and2_1 _20378_ (.A(_03817_),
    .B(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__clkbuf_1 _20379_ (.A(_03838_),
    .X(_01244_));
 sky130_fd_sc_hd__clkbuf_2 _20380_ (.A(_08244_),
    .X(_03839_));
 sky130_fd_sc_hd__mux2_1 _20381_ (.A0(\rbzero.pov.ready_buffer[57] ),
    .A1(\rbzero.pov.spi_buffer[57] ),
    .S(_03820_),
    .X(_03840_));
 sky130_fd_sc_hd__and2_1 _20382_ (.A(_03839_),
    .B(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__clkbuf_1 _20383_ (.A(_03841_),
    .X(_01245_));
 sky130_fd_sc_hd__clkbuf_4 _20384_ (.A(\rbzero.pov.spi_done ),
    .X(_03842_));
 sky130_fd_sc_hd__mux2_1 _20385_ (.A0(\rbzero.pov.ready_buffer[58] ),
    .A1(\rbzero.pov.spi_buffer[58] ),
    .S(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__and2_1 _20386_ (.A(_03839_),
    .B(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__clkbuf_1 _20387_ (.A(_03844_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _20388_ (.A0(\rbzero.pov.ready_buffer[59] ),
    .A1(\rbzero.pov.spi_buffer[59] ),
    .S(_03842_),
    .X(_03845_));
 sky130_fd_sc_hd__and2_1 _20389_ (.A(_03839_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_1 _20390_ (.A(_03846_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _20391_ (.A0(\rbzero.pov.ready_buffer[60] ),
    .A1(\rbzero.pov.spi_buffer[60] ),
    .S(_03842_),
    .X(_03847_));
 sky130_fd_sc_hd__and2_1 _20392_ (.A(_03839_),
    .B(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__clkbuf_1 _20393_ (.A(_03848_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _20394_ (.A0(\rbzero.pov.ready_buffer[61] ),
    .A1(\rbzero.pov.spi_buffer[61] ),
    .S(_03842_),
    .X(_03849_));
 sky130_fd_sc_hd__and2_1 _20395_ (.A(_03839_),
    .B(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__clkbuf_1 _20396_ (.A(_03850_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _20397_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(\rbzero.pov.spi_buffer[62] ),
    .S(_03842_),
    .X(_03851_));
 sky130_fd_sc_hd__and2_1 _20398_ (.A(_03839_),
    .B(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__clkbuf_1 _20399_ (.A(_03852_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _20400_ (.A0(\rbzero.pov.ready_buffer[63] ),
    .A1(\rbzero.pov.spi_buffer[63] ),
    .S(_03842_),
    .X(_03853_));
 sky130_fd_sc_hd__and2_1 _20401_ (.A(_03839_),
    .B(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__clkbuf_1 _20402_ (.A(_03854_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _20403_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(\rbzero.pov.spi_buffer[64] ),
    .S(_03842_),
    .X(_03855_));
 sky130_fd_sc_hd__and2_1 _20404_ (.A(_03839_),
    .B(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__clkbuf_1 _20405_ (.A(_03856_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _20406_ (.A0(\rbzero.pov.ready_buffer[65] ),
    .A1(\rbzero.pov.spi_buffer[65] ),
    .S(_03842_),
    .X(_03857_));
 sky130_fd_sc_hd__and2_1 _20407_ (.A(_03839_),
    .B(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_1 _20408_ (.A(_03858_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _20409_ (.A0(\rbzero.pov.ready_buffer[66] ),
    .A1(\rbzero.pov.spi_buffer[66] ),
    .S(_03842_),
    .X(_03859_));
 sky130_fd_sc_hd__and2_1 _20410_ (.A(_03839_),
    .B(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_1 _20411_ (.A(_03860_),
    .X(_01254_));
 sky130_fd_sc_hd__clkbuf_4 _20412_ (.A(_08244_),
    .X(_03861_));
 sky130_fd_sc_hd__mux2_1 _20413_ (.A0(\rbzero.pov.ready_buffer[67] ),
    .A1(\rbzero.pov.spi_buffer[67] ),
    .S(_03842_),
    .X(_03862_));
 sky130_fd_sc_hd__and2_1 _20414_ (.A(_03861_),
    .B(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__clkbuf_1 _20415_ (.A(_03863_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _20416_ (.A0(\rbzero.pov.ready_buffer[68] ),
    .A1(\rbzero.pov.spi_buffer[68] ),
    .S(_03731_),
    .X(_03864_));
 sky130_fd_sc_hd__and2_1 _20417_ (.A(_03861_),
    .B(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__clkbuf_1 _20418_ (.A(_03865_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _20419_ (.A0(\rbzero.pov.ready_buffer[69] ),
    .A1(\rbzero.pov.spi_buffer[69] ),
    .S(_03731_),
    .X(_03866_));
 sky130_fd_sc_hd__and2_1 _20420_ (.A(_03861_),
    .B(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__clkbuf_1 _20421_ (.A(_03867_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _20422_ (.A0(\rbzero.pov.ready_buffer[70] ),
    .A1(\rbzero.pov.spi_buffer[70] ),
    .S(_03731_),
    .X(_03868_));
 sky130_fd_sc_hd__and2_1 _20423_ (.A(_03861_),
    .B(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__clkbuf_1 _20424_ (.A(_03869_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _20425_ (.A0(\rbzero.pov.ready_buffer[71] ),
    .A1(\rbzero.pov.spi_buffer[71] ),
    .S(_03731_),
    .X(_03870_));
 sky130_fd_sc_hd__and2_1 _20426_ (.A(_03861_),
    .B(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _20427_ (.A(_03871_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _20428_ (.A0(\rbzero.pov.ready_buffer[72] ),
    .A1(\rbzero.pov.spi_buffer[72] ),
    .S(_03731_),
    .X(_03872_));
 sky130_fd_sc_hd__and2_1 _20429_ (.A(_03861_),
    .B(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_1 _20430_ (.A(_03873_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _20431_ (.A0(\rbzero.pov.ready_buffer[73] ),
    .A1(\rbzero.pov.spi_buffer[73] ),
    .S(_03731_),
    .X(_03874_));
 sky130_fd_sc_hd__and2_1 _20432_ (.A(_03861_),
    .B(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_1 _20433_ (.A(_03875_),
    .X(_01261_));
 sky130_fd_sc_hd__nor3b_1 _20434_ (.A(_03593_),
    .B(_03713_),
    .C_N(_03588_),
    .Y(_01262_));
 sky130_fd_sc_hd__and2_1 _20435_ (.A(_05772_),
    .B(_02850_),
    .X(_03876_));
 sky130_fd_sc_hd__clkbuf_1 _20436_ (.A(_03876_),
    .X(_01263_));
 sky130_fd_sc_hd__and2_1 _20437_ (.A(\rbzero.pov.mosi_buffer[0] ),
    .B(_02850_),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_1 _20438_ (.A(_03877_),
    .X(_01264_));
 sky130_fd_sc_hd__nand2_1 _20439_ (.A(_05261_),
    .B(_02855_),
    .Y(_03878_));
 sky130_fd_sc_hd__inv_2 _20440_ (.A(\gpout0.vpos[2] ),
    .Y(_03879_));
 sky130_fd_sc_hd__or4_1 _20441_ (.A(_04822_),
    .B(_03879_),
    .C(_05745_),
    .D(_05744_),
    .X(_03880_));
 sky130_fd_sc_hd__and3_1 _20442_ (.A(_05745_),
    .B(_05261_),
    .C(_02855_),
    .X(_03881_));
 sky130_fd_sc_hd__a41o_1 _20443_ (.A1(_05739_),
    .A2(_03879_),
    .A3(_04859_),
    .A4(_03881_),
    .B1(\rbzero.vga_sync.vsync ),
    .X(_03882_));
 sky130_fd_sc_hd__o211a_1 _20444_ (.A1(_03878_),
    .A2(_03880_),
    .B1(_03882_),
    .C1(_02883_),
    .X(_01265_));
 sky130_fd_sc_hd__and3b_1 _20445_ (.A_N(_04813_),
    .B(_04548_),
    .C(_04112_),
    .X(_03883_));
 sky130_fd_sc_hd__a31o_1 _20446_ (.A1(_04588_),
    .A2(_05392_),
    .A3(_03883_),
    .B1(_04544_),
    .X(_03884_));
 sky130_fd_sc_hd__a31o_1 _20447_ (.A1(_04107_),
    .A2(_09865_),
    .A3(_03883_),
    .B1(\rbzero.hsync ),
    .X(_03885_));
 sky130_fd_sc_hd__and2b_1 _20448_ (.A_N(_03884_),
    .B(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__clkbuf_1 _20449_ (.A(_03886_),
    .X(_01266_));
 sky130_fd_sc_hd__or4b_1 _20450_ (.A(_05177_),
    .B(_04866_),
    .C(_03880_),
    .D_N(_05746_),
    .X(_03887_));
 sky130_fd_sc_hd__and2_1 _20451_ (.A(_09867_),
    .B(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__nand2_1 _20452_ (.A(_05744_),
    .B(_09867_),
    .Y(_03889_));
 sky130_fd_sc_hd__o211a_1 _20453_ (.A1(_05744_),
    .A2(_03888_),
    .B1(_03889_),
    .C1(_02883_),
    .X(_01267_));
 sky130_fd_sc_hd__nand3_1 _20454_ (.A(_05745_),
    .B(_05744_),
    .C(_09867_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21o_1 _20455_ (.A1(_05744_),
    .A2(_09867_),
    .B1(_05745_),
    .X(_03891_));
 sky130_fd_sc_hd__and3_1 _20456_ (.A(_02850_),
    .B(_03890_),
    .C(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__clkbuf_1 _20457_ (.A(_03892_),
    .X(_01268_));
 sky130_fd_sc_hd__a21o_1 _20458_ (.A1(_08244_),
    .A2(_03887_),
    .B1(_09870_),
    .X(_03893_));
 sky130_fd_sc_hd__a21bo_1 _20459_ (.A1(_09867_),
    .A2(_02856_),
    .B1_N(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__a21oi_1 _20460_ (.A1(_03879_),
    .A2(_03890_),
    .B1(_03894_),
    .Y(_01269_));
 sky130_fd_sc_hd__clkbuf_8 _20461_ (.A(_09870_),
    .X(_03895_));
 sky130_fd_sc_hd__a21oi_1 _20462_ (.A1(_05739_),
    .A2(_02856_),
    .B1(_04544_),
    .Y(_03896_));
 sky130_fd_sc_hd__o21a_1 _20463_ (.A1(_05739_),
    .A2(_02856_),
    .B1(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__a22o_1 _20464_ (.A1(_05739_),
    .A2(_03895_),
    .B1(_03888_),
    .B2(_03897_),
    .X(_01270_));
 sky130_fd_sc_hd__and2_1 _20465_ (.A(_05742_),
    .B(_02857_),
    .X(_03898_));
 sky130_fd_sc_hd__inv_2 _20466_ (.A(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__o211a_1 _20467_ (.A1(_05742_),
    .A2(_02863_),
    .B1(_03899_),
    .C1(_02883_),
    .X(_01271_));
 sky130_fd_sc_hd__and3_1 _20468_ (.A(_04787_),
    .B(_05742_),
    .C(_02863_),
    .X(_03900_));
 sky130_fd_sc_hd__inv_2 _20469_ (.A(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__o211a_1 _20470_ (.A1(_04787_),
    .A2(_03898_),
    .B1(_03901_),
    .C1(_02883_),
    .X(_01272_));
 sky130_fd_sc_hd__nor2_1 _20471_ (.A(_04802_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__or2_1 _20472_ (.A(_04782_),
    .B(_03900_),
    .X(_03903_));
 sky130_fd_sc_hd__and3b_1 _20473_ (.A_N(_03902_),
    .B(_08245_),
    .C(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__clkbuf_1 _20474_ (.A(_03904_),
    .X(_01273_));
 sky130_fd_sc_hd__o21ai_1 _20475_ (.A1(_04775_),
    .A2(_03902_),
    .B1(_08246_),
    .Y(_03905_));
 sky130_fd_sc_hd__a21oi_1 _20476_ (.A1(_05178_),
    .A2(_03898_),
    .B1(_03905_),
    .Y(_01274_));
 sky130_fd_sc_hd__and3_1 _20477_ (.A(_04787_),
    .B(_02854_),
    .C(_03898_),
    .X(_03906_));
 sky130_fd_sc_hd__a31o_1 _20478_ (.A1(_05742_),
    .A2(_05178_),
    .A3(_02857_),
    .B1(_05177_),
    .X(_03907_));
 sky130_fd_sc_hd__and3b_1 _20479_ (.A_N(_03906_),
    .B(_08245_),
    .C(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__clkbuf_1 _20480_ (.A(_03908_),
    .X(_01275_));
 sky130_fd_sc_hd__or2_1 _20481_ (.A(_05746_),
    .B(_03906_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_1 _20482_ (.A(_05746_),
    .B(_03906_),
    .Y(_03910_));
 sky130_fd_sc_hd__and3_1 _20483_ (.A(_03893_),
    .B(_03909_),
    .C(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__clkbuf_1 _20484_ (.A(_03911_),
    .X(_01276_));
 sky130_fd_sc_hd__a31o_1 _20485_ (.A1(\rbzero.spi_registers.got_new_texadd3 ),
    .A2(_08246_),
    .A3(_02881_),
    .B1(_02492_),
    .X(_01277_));
 sky130_fd_sc_hd__inv_2 _20487__93 (.A(clknet_1_1__leaf__03712_),
    .Y(net218));
 sky130_fd_sc_hd__inv_2 _20488__94 (.A(clknet_1_1__leaf__03712_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _20489__95 (.A(clknet_1_1__leaf__03712_),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _20490__96 (.A(clknet_1_1__leaf__03712_),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _20491__97 (.A(clknet_1_1__leaf__03712_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _20493__98 (.A(clknet_1_0__leaf__03912_),
    .Y(net223));
 sky130_fd_sc_hd__buf_1 _20492_ (.A(clknet_1_1__leaf__03711_),
    .X(_03912_));
 sky130_fd_sc_hd__inv_2 _20494__99 (.A(clknet_1_0__leaf__03912_),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _20495__100 (.A(clknet_1_1__leaf__03912_),
    .Y(net225));
 sky130_fd_sc_hd__inv_2 _20496__101 (.A(clknet_1_1__leaf__03912_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _20497__102 (.A(clknet_1_1__leaf__03912_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _20498__103 (.A(clknet_1_0__leaf__03912_),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _20499__104 (.A(clknet_1_0__leaf__03912_),
    .Y(net229));
 sky130_fd_sc_hd__inv_2 _20500__105 (.A(clknet_1_0__leaf__03912_),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _20501__106 (.A(clknet_1_1__leaf__03912_),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _20502__107 (.A(clknet_1_1__leaf__03912_),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _20504__108 (.A(clknet_1_1__leaf__03913_),
    .Y(net233));
 sky130_fd_sc_hd__buf_1 _20503_ (.A(clknet_1_1__leaf__03711_),
    .X(_03913_));
 sky130_fd_sc_hd__inv_2 _20505__109 (.A(clknet_1_1__leaf__03913_),
    .Y(net234));
 sky130_fd_sc_hd__inv_2 _20506__110 (.A(clknet_1_1__leaf__03913_),
    .Y(net235));
 sky130_fd_sc_hd__inv_2 _20507__111 (.A(clknet_1_1__leaf__03913_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _20508__112 (.A(clknet_1_1__leaf__03913_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _20509__113 (.A(clknet_1_0__leaf__03913_),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _20510__114 (.A(clknet_1_0__leaf__03913_),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _20511__115 (.A(clknet_1_0__leaf__03913_),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _20512__116 (.A(clknet_1_0__leaf__03913_),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _20513__117 (.A(clknet_1_0__leaf__03913_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _20515__118 (.A(clknet_1_1__leaf__03914_),
    .Y(net243));
 sky130_fd_sc_hd__buf_1 _20514_ (.A(clknet_1_1__leaf__03711_),
    .X(_03914_));
 sky130_fd_sc_hd__inv_2 _20516__119 (.A(clknet_1_1__leaf__03914_),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _20517__120 (.A(clknet_1_1__leaf__03914_),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _20518__121 (.A(clknet_1_0__leaf__03914_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _20519__122 (.A(clknet_1_0__leaf__03914_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _20520__123 (.A(clknet_1_0__leaf__03914_),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _20521__124 (.A(clknet_1_0__leaf__03914_),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _20522__125 (.A(clknet_1_0__leaf__03914_),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _20523__126 (.A(clknet_1_0__leaf__03914_),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _20524__127 (.A(clknet_1_1__leaf__03914_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _20526__128 (.A(clknet_1_0__leaf__03915_),
    .Y(net253));
 sky130_fd_sc_hd__buf_1 _20525_ (.A(clknet_1_0__leaf__03711_),
    .X(_03915_));
 sky130_fd_sc_hd__inv_2 _20527__129 (.A(clknet_1_0__leaf__03915_),
    .Y(net254));
 sky130_fd_sc_hd__inv_2 _20528__130 (.A(clknet_1_0__leaf__03915_),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _20529__131 (.A(clknet_1_1__leaf__03915_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _20530__132 (.A(clknet_1_1__leaf__03915_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _20531__133 (.A(clknet_1_1__leaf__03915_),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _20532__134 (.A(clknet_1_1__leaf__03915_),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _20533__135 (.A(clknet_1_1__leaf__03915_),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _20534__136 (.A(clknet_1_1__leaf__03915_),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _20535__137 (.A(clknet_1_0__leaf__03915_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _20537__138 (.A(clknet_1_1__leaf__03916_),
    .Y(net263));
 sky130_fd_sc_hd__buf_1 _20536_ (.A(clknet_1_0__leaf__03711_),
    .X(_03916_));
 sky130_fd_sc_hd__inv_2 _20538__139 (.A(clknet_1_1__leaf__03916_),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _20539__140 (.A(clknet_1_1__leaf__03916_),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _20540__141 (.A(clknet_1_1__leaf__03916_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _20541__142 (.A(clknet_1_1__leaf__03916_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _20542__143 (.A(clknet_1_0__leaf__03916_),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _20543__144 (.A(clknet_1_0__leaf__03916_),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _20544__145 (.A(clknet_1_0__leaf__03916_),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _20545__146 (.A(clknet_1_0__leaf__03916_),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _20546__147 (.A(clknet_1_0__leaf__03916_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _20548__148 (.A(clknet_1_1__leaf__03917_),
    .Y(net273));
 sky130_fd_sc_hd__buf_1 _20547_ (.A(clknet_1_0__leaf__03711_),
    .X(_03917_));
 sky130_fd_sc_hd__inv_2 _20549__149 (.A(clknet_1_1__leaf__03917_),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _20550__150 (.A(clknet_1_1__leaf__03917_),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _20551__151 (.A(clknet_1_1__leaf__03917_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _20552__152 (.A(clknet_1_1__leaf__03917_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _20553__153 (.A(clknet_1_0__leaf__03917_),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _20554__154 (.A(clknet_1_0__leaf__03917_),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _20555__155 (.A(clknet_1_0__leaf__03917_),
    .Y(net280));
 sky130_fd_sc_hd__inv_2 _20556__156 (.A(clknet_1_0__leaf__03917_),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _20557__157 (.A(clknet_1_0__leaf__03917_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _20559__158 (.A(clknet_1_1__leaf__03918_),
    .Y(net283));
 sky130_fd_sc_hd__buf_1 _20558_ (.A(clknet_1_0__leaf__03711_),
    .X(_03918_));
 sky130_fd_sc_hd__inv_2 _20560__159 (.A(clknet_1_1__leaf__03918_),
    .Y(net284));
 sky130_fd_sc_hd__inv_2 _20561__160 (.A(clknet_1_0__leaf__03918_),
    .Y(net285));
 sky130_fd_sc_hd__inv_2 _20562__161 (.A(clknet_1_0__leaf__03918_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _20563__162 (.A(clknet_1_0__leaf__03918_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _20564__163 (.A(clknet_1_0__leaf__03918_),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _20565__164 (.A(clknet_1_0__leaf__03918_),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _20566__165 (.A(clknet_1_0__leaf__03918_),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _20567__166 (.A(clknet_1_1__leaf__03918_),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _20568__167 (.A(clknet_1_1__leaf__03918_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _20570__168 (.A(clknet_1_0__leaf__03919_),
    .Y(net293));
 sky130_fd_sc_hd__buf_1 _20569_ (.A(clknet_1_0__leaf__03711_),
    .X(_03919_));
 sky130_fd_sc_hd__inv_2 _20571__169 (.A(clknet_1_0__leaf__03919_),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _20572__170 (.A(clknet_1_0__leaf__03919_),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _20573__171 (.A(clknet_1_0__leaf__03919_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _20574__172 (.A(clknet_1_0__leaf__03919_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _20575__173 (.A(clknet_1_1__leaf__03919_),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _20576__174 (.A(clknet_1_1__leaf__03919_),
    .Y(net299));
 sky130_fd_sc_hd__inv_2 _20577__175 (.A(clknet_1_1__leaf__03919_),
    .Y(net300));
 sky130_fd_sc_hd__inv_2 _20578__176 (.A(clknet_1_1__leaf__03919_),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _20579__177 (.A(clknet_1_1__leaf__03919_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _20581__178 (.A(clknet_1_0__leaf__03920_),
    .Y(net303));
 sky130_fd_sc_hd__buf_1 _20580_ (.A(clknet_1_1__leaf__03711_),
    .X(_03920_));
 sky130_fd_sc_hd__inv_2 _20582__179 (.A(clknet_1_0__leaf__03920_),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _20583__180 (.A(clknet_1_0__leaf__03920_),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _20584__181 (.A(clknet_1_0__leaf__03920_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _20585__182 (.A(clknet_1_0__leaf__03920_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _20586__183 (.A(clknet_1_1__leaf__03920_),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _20587__184 (.A(clknet_1_1__leaf__03920_),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _20588__185 (.A(clknet_1_1__leaf__03920_),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 _20589__186 (.A(clknet_1_1__leaf__03920_),
    .Y(net311));
 sky130_fd_sc_hd__inv_2 _20590__187 (.A(clknet_1_1__leaf__03920_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _20593__188 (.A(clknet_1_1__leaf__03922_),
    .Y(net313));
 sky130_fd_sc_hd__buf_1 _20591_ (.A(clknet_1_0__leaf__04767_),
    .X(_03921_));
 sky130_fd_sc_hd__buf_1 _20592_ (.A(clknet_1_1__leaf__03921_),
    .X(_03922_));
 sky130_fd_sc_hd__inv_2 _20594__189 (.A(clknet_1_1__leaf__03922_),
    .Y(net314));
 sky130_fd_sc_hd__inv_2 _20595__190 (.A(clknet_1_1__leaf__03922_),
    .Y(net315));
 sky130_fd_sc_hd__inv_2 _20596__191 (.A(clknet_1_1__leaf__03922_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _20597__192 (.A(clknet_1_1__leaf__03922_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _20598__193 (.A(clknet_1_0__leaf__03922_),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _20599__194 (.A(clknet_1_0__leaf__03922_),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 _20600__195 (.A(clknet_1_0__leaf__03922_),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _20601__196 (.A(clknet_1_0__leaf__03922_),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _20602__197 (.A(clknet_1_0__leaf__03922_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _20604__198 (.A(clknet_1_1__leaf__03923_),
    .Y(net323));
 sky130_fd_sc_hd__buf_1 _20603_ (.A(clknet_1_0__leaf__03921_),
    .X(_03923_));
 sky130_fd_sc_hd__inv_2 _20605__199 (.A(clknet_1_1__leaf__03923_),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _20606__200 (.A(clknet_1_0__leaf__03923_),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _20607__201 (.A(clknet_1_0__leaf__03923_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _20608__202 (.A(clknet_1_0__leaf__03923_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _20609__203 (.A(clknet_1_0__leaf__03923_),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _20610__204 (.A(clknet_1_0__leaf__03923_),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _20611__205 (.A(clknet_1_1__leaf__03923_),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _20612__206 (.A(clknet_1_1__leaf__03923_),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _20613__207 (.A(clknet_1_1__leaf__03923_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _20615__208 (.A(clknet_1_0__leaf__03924_),
    .Y(net333));
 sky130_fd_sc_hd__buf_1 _20614_ (.A(clknet_1_1__leaf__03921_),
    .X(_03924_));
 sky130_fd_sc_hd__inv_2 _20616__209 (.A(clknet_1_1__leaf__03924_),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _20617__210 (.A(clknet_1_1__leaf__03924_),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _20618__211 (.A(clknet_1_1__leaf__03924_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _20619__212 (.A(clknet_1_1__leaf__03924_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _20620__213 (.A(clknet_1_1__leaf__03924_),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _20621__214 (.A(clknet_1_0__leaf__03924_),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _20622__215 (.A(clknet_1_0__leaf__03924_),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _20623__216 (.A(clknet_1_0__leaf__03924_),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _20624__217 (.A(clknet_1_0__leaf__03924_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _20626__218 (.A(clknet_1_1__leaf__03925_),
    .Y(net343));
 sky130_fd_sc_hd__buf_1 _20625_ (.A(clknet_1_0__leaf__03921_),
    .X(_03925_));
 sky130_fd_sc_hd__inv_2 _20627__219 (.A(clknet_1_1__leaf__03925_),
    .Y(net344));
 sky130_fd_sc_hd__inv_2 _20628__220 (.A(clknet_1_1__leaf__03925_),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _20629__221 (.A(clknet_1_1__leaf__03925_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _20630__222 (.A(clknet_1_0__leaf__03925_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _20631__223 (.A(clknet_1_0__leaf__03925_),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _20632__224 (.A(clknet_1_0__leaf__03925_),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _20633__225 (.A(clknet_1_0__leaf__03925_),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _20634__226 (.A(clknet_1_0__leaf__03925_),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _20635__227 (.A(clknet_1_0__leaf__03925_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _20637__228 (.A(clknet_1_1__leaf__03926_),
    .Y(net353));
 sky130_fd_sc_hd__buf_1 _20636_ (.A(clknet_1_0__leaf__03921_),
    .X(_03926_));
 sky130_fd_sc_hd__inv_2 _20638__229 (.A(clknet_1_1__leaf__03926_),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _20639__230 (.A(clknet_1_1__leaf__03926_),
    .Y(net355));
 sky130_fd_sc_hd__inv_2 _20640__231 (.A(clknet_1_1__leaf__03926_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _20641__232 (.A(clknet_1_0__leaf__03926_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _20642__233 (.A(clknet_1_0__leaf__03926_),
    .Y(net358));
 sky130_fd_sc_hd__inv_2 _20643__234 (.A(clknet_1_0__leaf__03926_),
    .Y(net359));
 sky130_fd_sc_hd__inv_2 _20644__235 (.A(clknet_1_0__leaf__03926_),
    .Y(net360));
 sky130_fd_sc_hd__inv_2 _20645__236 (.A(clknet_1_0__leaf__03926_),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 _20646__237 (.A(clknet_1_0__leaf__03926_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _20648__238 (.A(clknet_1_0__leaf__03927_),
    .Y(net363));
 sky130_fd_sc_hd__buf_1 _20647_ (.A(clknet_1_0__leaf__03921_),
    .X(_03927_));
 sky130_fd_sc_hd__inv_2 _20649__239 (.A(clknet_1_0__leaf__03927_),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _20650__240 (.A(clknet_1_0__leaf__03927_),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _20651__241 (.A(clknet_1_0__leaf__03927_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _20652__242 (.A(clknet_1_1__leaf__03927_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _20653__243 (.A(clknet_1_1__leaf__03927_),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _20654__244 (.A(clknet_1_1__leaf__03927_),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _20655__245 (.A(clknet_1_1__leaf__03927_),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _20656__246 (.A(clknet_1_1__leaf__03927_),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _20657__247 (.A(clknet_1_1__leaf__03927_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _20659__248 (.A(clknet_1_0__leaf__03928_),
    .Y(net373));
 sky130_fd_sc_hd__buf_1 _20658_ (.A(clknet_1_1__leaf__03921_),
    .X(_03928_));
 sky130_fd_sc_hd__inv_2 _20660__249 (.A(clknet_1_0__leaf__03928_),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _20661__250 (.A(clknet_1_0__leaf__03928_),
    .Y(net375));
 sky130_fd_sc_hd__inv_2 _20662__251 (.A(clknet_1_0__leaf__03928_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _20663__252 (.A(clknet_1_1__leaf__03928_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _20664__253 (.A(clknet_1_1__leaf__03928_),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _20665__254 (.A(clknet_1_1__leaf__03928_),
    .Y(net379));
 sky130_fd_sc_hd__inv_2 _20666__255 (.A(clknet_1_1__leaf__03928_),
    .Y(net380));
 sky130_fd_sc_hd__inv_2 _20667__256 (.A(clknet_1_1__leaf__03928_),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _20668__257 (.A(clknet_1_1__leaf__03928_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _20670__258 (.A(clknet_1_0__leaf__03929_),
    .Y(net383));
 sky130_fd_sc_hd__buf_1 _20669_ (.A(clknet_1_1__leaf__03921_),
    .X(_03929_));
 sky130_fd_sc_hd__inv_2 _20671__259 (.A(clknet_1_0__leaf__03929_),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _20672__260 (.A(clknet_1_0__leaf__03929_),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _20673__261 (.A(clknet_1_0__leaf__03929_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _20674__262 (.A(clknet_1_1__leaf__03929_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _20675__263 (.A(clknet_1_1__leaf__03929_),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _20676__264 (.A(clknet_1_1__leaf__03929_),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _20677__265 (.A(clknet_1_1__leaf__03929_),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _20678__266 (.A(clknet_1_1__leaf__03929_),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _20679__267 (.A(clknet_1_1__leaf__03929_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _20681__268 (.A(clknet_1_1__leaf__03930_),
    .Y(net393));
 sky130_fd_sc_hd__buf_1 _20680_ (.A(clknet_1_1__leaf__03921_),
    .X(_03930_));
 sky130_fd_sc_hd__inv_2 _20682__269 (.A(clknet_1_1__leaf__03930_),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _20683__270 (.A(clknet_1_1__leaf__03930_),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _20684__271 (.A(clknet_1_0__leaf__03930_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _20685__272 (.A(clknet_1_0__leaf__03930_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _20686__273 (.A(clknet_1_0__leaf__03930_),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _20687__274 (.A(clknet_1_0__leaf__03930_),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _20688__275 (.A(clknet_1_0__leaf__03930_),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _20689__276 (.A(clknet_1_1__leaf__03930_),
    .Y(net401));
 sky130_fd_sc_hd__inv_2 _20690__277 (.A(clknet_1_1__leaf__03930_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _20692__278 (.A(clknet_1_0__leaf__03931_),
    .Y(net403));
 sky130_fd_sc_hd__buf_1 _20691_ (.A(clknet_1_1__leaf__03921_),
    .X(_03931_));
 sky130_fd_sc_hd__inv_2 _20693__279 (.A(clknet_1_0__leaf__03931_),
    .Y(net404));
 sky130_fd_sc_hd__inv_2 _20694__280 (.A(clknet_1_0__leaf__03931_),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _20695__281 (.A(clknet_1_0__leaf__03931_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _20696__282 (.A(clknet_1_1__leaf__03931_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _20697__283 (.A(clknet_1_0__leaf__03931_),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _20698__284 (.A(clknet_1_1__leaf__03931_),
    .Y(net409));
 sky130_fd_sc_hd__inv_2 _20699__285 (.A(clknet_1_1__leaf__03931_),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _20700__286 (.A(clknet_1_1__leaf__03931_),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _20701__287 (.A(clknet_1_1__leaf__03931_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _20704__288 (.A(clknet_1_0__leaf__03933_),
    .Y(net413));
 sky130_fd_sc_hd__buf_1 _20702_ (.A(clknet_1_1__leaf__04767_),
    .X(_03932_));
 sky130_fd_sc_hd__buf_1 _20703_ (.A(clknet_1_0__leaf__03932_),
    .X(_03933_));
 sky130_fd_sc_hd__inv_2 _20705__289 (.A(clknet_1_0__leaf__03933_),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _20706__290 (.A(clknet_1_0__leaf__03933_),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _20707__291 (.A(clknet_1_0__leaf__03933_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _20708__292 (.A(clknet_1_1__leaf__03933_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _20709__293 (.A(clknet_1_1__leaf__03933_),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _20710__294 (.A(clknet_1_1__leaf__03933_),
    .Y(net419));
 sky130_fd_sc_hd__inv_2 _20711__295 (.A(clknet_1_1__leaf__03933_),
    .Y(net420));
 sky130_fd_sc_hd__inv_2 _20712__296 (.A(clknet_1_1__leaf__03933_),
    .Y(net421));
 sky130_fd_sc_hd__inv_2 _20713__297 (.A(clknet_1_1__leaf__03933_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _20715__298 (.A(clknet_1_0__leaf__03934_),
    .Y(net423));
 sky130_fd_sc_hd__buf_1 _20714_ (.A(clknet_1_0__leaf__03932_),
    .X(_03934_));
 sky130_fd_sc_hd__inv_2 _20716__299 (.A(clknet_1_0__leaf__03934_),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _20717__300 (.A(clknet_1_1__leaf__03934_),
    .Y(net425));
 sky130_fd_sc_hd__inv_2 _20718__301 (.A(clknet_1_1__leaf__03934_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _20719__302 (.A(clknet_1_1__leaf__03934_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _20720__303 (.A(clknet_1_1__leaf__03934_),
    .Y(net428));
 sky130_fd_sc_hd__inv_2 _20721__304 (.A(clknet_1_1__leaf__03934_),
    .Y(net429));
 sky130_fd_sc_hd__inv_2 _20722__305 (.A(clknet_1_1__leaf__03934_),
    .Y(net430));
 sky130_fd_sc_hd__inv_2 _20723__306 (.A(clknet_1_0__leaf__03934_),
    .Y(net431));
 sky130_fd_sc_hd__inv_2 _20724__307 (.A(clknet_1_0__leaf__03934_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _20726__308 (.A(clknet_1_1__leaf__03935_),
    .Y(net433));
 sky130_fd_sc_hd__buf_1 _20725_ (.A(clknet_1_1__leaf__03932_),
    .X(_03935_));
 sky130_fd_sc_hd__inv_2 _20727__309 (.A(clknet_1_0__leaf__03935_),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _20728__310 (.A(clknet_1_0__leaf__03935_),
    .Y(net435));
 sky130_fd_sc_hd__inv_2 _20729__311 (.A(clknet_1_0__leaf__03935_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _20730__312 (.A(clknet_1_0__leaf__03935_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _20731__313 (.A(clknet_1_0__leaf__03935_),
    .Y(net438));
 sky130_fd_sc_hd__inv_2 _20732__314 (.A(clknet_1_0__leaf__03935_),
    .Y(net439));
 sky130_fd_sc_hd__inv_2 _20733__315 (.A(clknet_1_1__leaf__03935_),
    .Y(net440));
 sky130_fd_sc_hd__inv_2 _20734__316 (.A(clknet_1_1__leaf__03935_),
    .Y(net441));
 sky130_fd_sc_hd__inv_2 _20735__317 (.A(clknet_1_1__leaf__03935_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _20737__318 (.A(clknet_1_1__leaf__03936_),
    .Y(net443));
 sky130_fd_sc_hd__buf_1 _20736_ (.A(clknet_1_1__leaf__03932_),
    .X(_03936_));
 sky130_fd_sc_hd__inv_2 _20738__319 (.A(clknet_1_1__leaf__03936_),
    .Y(net444));
 sky130_fd_sc_hd__inv_2 _20739__320 (.A(clknet_1_1__leaf__03936_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _20740__321 (.A(clknet_1_0__leaf__03936_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _20741__322 (.A(clknet_1_0__leaf__03936_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _20742__323 (.A(clknet_1_0__leaf__03936_),
    .Y(net448));
 sky130_fd_sc_hd__inv_2 _20743__324 (.A(clknet_1_0__leaf__03936_),
    .Y(net449));
 sky130_fd_sc_hd__inv_2 _20744__325 (.A(clknet_1_0__leaf__03936_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _20745__326 (.A(clknet_1_1__leaf__03936_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _20746__327 (.A(clknet_1_1__leaf__03936_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _20748__328 (.A(clknet_1_0__leaf__03937_),
    .Y(net453));
 sky130_fd_sc_hd__buf_1 _20747_ (.A(clknet_1_1__leaf__03932_),
    .X(_03937_));
 sky130_fd_sc_hd__inv_2 _20749__329 (.A(clknet_1_0__leaf__03937_),
    .Y(net454));
 sky130_fd_sc_hd__inv_2 _20750__330 (.A(clknet_1_0__leaf__03937_),
    .Y(net455));
 sky130_fd_sc_hd__inv_2 _20751__331 (.A(clknet_1_1__leaf__03937_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _20752__332 (.A(clknet_1_1__leaf__03937_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _20753__333 (.A(clknet_1_0__leaf__03937_),
    .Y(net458));
 sky130_fd_sc_hd__inv_2 _20754__334 (.A(clknet_1_0__leaf__03937_),
    .Y(net459));
 sky130_fd_sc_hd__inv_2 _20755__335 (.A(clknet_1_1__leaf__03937_),
    .Y(net460));
 sky130_fd_sc_hd__inv_2 _20756__336 (.A(clknet_1_1__leaf__03937_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _20757__337 (.A(clknet_1_1__leaf__03937_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _20759__338 (.A(clknet_1_1__leaf__03938_),
    .Y(net463));
 sky130_fd_sc_hd__buf_1 _20758_ (.A(clknet_1_1__leaf__03932_),
    .X(_03938_));
 sky130_fd_sc_hd__inv_2 _20760__339 (.A(clknet_1_1__leaf__03938_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _20761__340 (.A(clknet_1_1__leaf__03938_),
    .Y(net465));
 sky130_fd_sc_hd__inv_2 _20762__341 (.A(clknet_1_1__leaf__03938_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _20763__342 (.A(clknet_1_1__leaf__03938_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _20764__343 (.A(clknet_1_0__leaf__03938_),
    .Y(net468));
 sky130_fd_sc_hd__inv_2 _20765__344 (.A(clknet_1_0__leaf__03938_),
    .Y(net469));
 sky130_fd_sc_hd__inv_2 _20766__345 (.A(clknet_1_0__leaf__03938_),
    .Y(net470));
 sky130_fd_sc_hd__inv_2 _20767__346 (.A(clknet_1_0__leaf__03938_),
    .Y(net471));
 sky130_fd_sc_hd__inv_2 _20768__347 (.A(clknet_1_0__leaf__03938_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _20770__348 (.A(clknet_1_0__leaf__03939_),
    .Y(net473));
 sky130_fd_sc_hd__buf_1 _20769_ (.A(clknet_1_0__leaf__03932_),
    .X(_03939_));
 sky130_fd_sc_hd__inv_2 _20771__349 (.A(clknet_1_0__leaf__03939_),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _20772__350 (.A(clknet_1_0__leaf__03939_),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _20773__351 (.A(clknet_1_0__leaf__03939_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _20774__352 (.A(clknet_1_0__leaf__03939_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _20775__353 (.A(clknet_1_1__leaf__03939_),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _20776__354 (.A(clknet_1_1__leaf__03939_),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _20777__355 (.A(clknet_1_1__leaf__03939_),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _20778__356 (.A(clknet_1_1__leaf__03939_),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _20779__357 (.A(clknet_1_1__leaf__03939_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _20781__358 (.A(clknet_1_0__leaf__03940_),
    .Y(net483));
 sky130_fd_sc_hd__buf_1 _20780_ (.A(clknet_1_0__leaf__03932_),
    .X(_03940_));
 sky130_fd_sc_hd__inv_2 _20782__359 (.A(clknet_1_0__leaf__03940_),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _20783__360 (.A(clknet_1_0__leaf__03940_),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _20784__361 (.A(clknet_1_0__leaf__03940_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _20785__362 (.A(clknet_1_0__leaf__03940_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _20786__363 (.A(clknet_1_0__leaf__03940_),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _20787__364 (.A(clknet_1_1__leaf__03940_),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _20788__365 (.A(clknet_1_1__leaf__03940_),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _20789__366 (.A(clknet_1_1__leaf__03940_),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _20790__367 (.A(clknet_1_1__leaf__03940_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _20792__368 (.A(clknet_1_0__leaf__03941_),
    .Y(net493));
 sky130_fd_sc_hd__buf_1 _20791_ (.A(clknet_1_0__leaf__03932_),
    .X(_03941_));
 sky130_fd_sc_hd__inv_2 _20793__369 (.A(clknet_1_0__leaf__03941_),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _20794__370 (.A(clknet_1_0__leaf__03941_),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _20795__371 (.A(clknet_1_0__leaf__03941_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _20796__372 (.A(clknet_1_0__leaf__03941_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _20797__373 (.A(clknet_1_0__leaf__03941_),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _20798__374 (.A(clknet_1_1__leaf__03941_),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _20799__375 (.A(clknet_1_1__leaf__03941_),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _20800__376 (.A(clknet_1_1__leaf__03941_),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _20801__377 (.A(clknet_1_1__leaf__03941_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _20803__378 (.A(clknet_1_1__leaf__03942_),
    .Y(net503));
 sky130_fd_sc_hd__buf_1 _20802_ (.A(clknet_1_0__leaf__03932_),
    .X(_03942_));
 sky130_fd_sc_hd__inv_2 _20804__379 (.A(clknet_1_1__leaf__03942_),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _20805__380 (.A(clknet_1_0__leaf__03942_),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _20806__381 (.A(clknet_1_0__leaf__03942_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _20807__382 (.A(clknet_1_0__leaf__03942_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _20808__383 (.A(clknet_1_0__leaf__03942_),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _20809__384 (.A(clknet_1_0__leaf__03942_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _20810__385 (.A(clknet_1_1__leaf__03942_),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _20811__386 (.A(clknet_1_1__leaf__03942_),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _20812__387 (.A(clknet_1_1__leaf__03942_),
    .Y(net512));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__buf_1 _20813_ (.A(clknet_1_1__leaf__04767_),
    .X(_03943_));
 sky130_fd_sc_hd__inv_2 _20815__9 (.A(clknet_1_0__leaf__03943_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _20816__10 (.A(clknet_1_0__leaf__03943_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _20817__11 (.A(clknet_1_0__leaf__03943_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _20818__12 (.A(clknet_1_0__leaf__03943_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _20819__13 (.A(clknet_1_1__leaf__03943_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _20820__14 (.A(clknet_1_1__leaf__03943_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _20821__15 (.A(clknet_1_1__leaf__03943_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _20822__16 (.A(clknet_1_1__leaf__03943_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _20823__17 (.A(clknet_1_1__leaf__03943_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _20825__18 (.A(clknet_1_1__leaf__03944_),
    .Y(net143));
 sky130_fd_sc_hd__buf_1 _20824_ (.A(clknet_1_1__leaf__04767_),
    .X(_03944_));
 sky130_fd_sc_hd__inv_2 _20826__19 (.A(clknet_1_1__leaf__03944_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _20827__20 (.A(clknet_1_1__leaf__03944_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _20828__21 (.A(clknet_1_1__leaf__03944_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _20829__22 (.A(clknet_1_1__leaf__03944_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _20830__23 (.A(clknet_1_0__leaf__03944_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _20831__24 (.A(clknet_1_1__leaf__03944_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _20832__25 (.A(clknet_1_0__leaf__03944_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _20833__26 (.A(clknet_1_0__leaf__03944_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _20834__27 (.A(clknet_1_0__leaf__03944_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _20125__28 (.A(clknet_1_1__leaf__03705_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _20836__5 (.A(clknet_1_1__leaf__03704_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _20837__6 (.A(clknet_1_1__leaf__03704_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _20838__7 (.A(clknet_1_1__leaf__03704_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _20814__8 (.A(clknet_1_0__leaf__03943_),
    .Y(net133));
 sky130_fd_sc_hd__nor2_1 _20839_ (.A(\gpout5.clk_div[0] ),
    .B(net64),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_1 _20840_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .Y(_03945_));
 sky130_fd_sc_hd__or2_1 _20841_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .X(_03946_));
 sky130_fd_sc_hd__and3_1 _20842_ (.A(_02850_),
    .B(_03945_),
    .C(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__clkbuf_1 _20843_ (.A(_03947_),
    .X(_01599_));
 sky130_fd_sc_hd__clkbuf_4 _20844_ (.A(_09870_),
    .X(_03948_));
 sky130_fd_sc_hd__nand2_1 _20845_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .Y(_03949_));
 sky130_fd_sc_hd__or2_1 _20846_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .X(_03950_));
 sky130_fd_sc_hd__clkbuf_4 _20847_ (.A(_04545_),
    .X(_03951_));
 sky130_fd_sc_hd__a32o_1 _20848_ (.A1(_03948_),
    .A2(_03949_),
    .A3(_03950_),
    .B1(_03951_),
    .B2(\rbzero.texV[-11] ),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _20849_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .X(_03952_));
 sky130_fd_sc_hd__nand2_1 _20850_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03953_));
 sky130_fd_sc_hd__nand3b_1 _20851_ (.A_N(_03949_),
    .B(_03952_),
    .C(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__a21bo_1 _20852_ (.A1(_03952_),
    .A2(_03953_),
    .B1_N(_03949_),
    .X(_03955_));
 sky130_fd_sc_hd__a32o_1 _20853_ (.A1(_03948_),
    .A2(_03954_),
    .A3(_03955_),
    .B1(_03951_),
    .B2(\rbzero.texV[-10] ),
    .X(_01601_));
 sky130_fd_sc_hd__and2_1 _20854_ (.A(_03953_),
    .B(_03954_),
    .X(_03956_));
 sky130_fd_sc_hd__nor2_1 _20855_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03957_));
 sky130_fd_sc_hd__nand2_1 _20856_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03958_));
 sky130_fd_sc_hd__and2b_1 _20857_ (.A_N(_03957_),
    .B(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__xnor2_1 _20858_ (.A(_03956_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__a22o_1 _20859_ (.A1(\rbzero.texV[-9] ),
    .A2(_03567_),
    .B1(_03895_),
    .B2(_03960_),
    .X(_01602_));
 sky130_fd_sc_hd__or2_1 _20860_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .X(_03961_));
 sky130_fd_sc_hd__nand2_1 _20861_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_1 _20862_ (.A(_03961_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__o21ai_1 _20863_ (.A1(_03956_),
    .A2(_03957_),
    .B1(_03958_),
    .Y(_03964_));
 sky130_fd_sc_hd__xnor2_1 _20864_ (.A(_03963_),
    .B(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hd__a22o_1 _20865_ (.A1(\rbzero.texV[-8] ),
    .A2(_03567_),
    .B1(_03895_),
    .B2(_03965_),
    .X(_01603_));
 sky130_fd_sc_hd__nor2_1 _20866_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .Y(_03966_));
 sky130_fd_sc_hd__and2_1 _20867_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .X(_03967_));
 sky130_fd_sc_hd__a21boi_1 _20868_ (.A1(_03961_),
    .A2(_03964_),
    .B1_N(_03962_),
    .Y(_03968_));
 sky130_fd_sc_hd__o21ai_1 _20869_ (.A1(_03966_),
    .A2(_03967_),
    .B1(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__or3_1 _20870_ (.A(_03966_),
    .B(_03967_),
    .C(_03968_),
    .X(_03970_));
 sky130_fd_sc_hd__a32o_1 _20871_ (.A1(_03948_),
    .A2(_03969_),
    .A3(_03970_),
    .B1(_03951_),
    .B2(\rbzero.texV[-7] ),
    .X(_01604_));
 sky130_fd_sc_hd__or2_1 _20872_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .X(_03971_));
 sky130_fd_sc_hd__nand2_1 _20873_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_03972_));
 sky130_fd_sc_hd__o21bai_1 _20874_ (.A1(_03966_),
    .A2(_03968_),
    .B1_N(_03967_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand3_1 _20875_ (.A(_03971_),
    .B(_03972_),
    .C(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__a21o_1 _20876_ (.A1(_03971_),
    .A2(_03972_),
    .B1(_03973_),
    .X(_03975_));
 sky130_fd_sc_hd__a32o_1 _20877_ (.A1(_03948_),
    .A2(_03974_),
    .A3(_03975_),
    .B1(_03951_),
    .B2(\rbzero.texV[-6] ),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _20878_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_03976_));
 sky130_fd_sc_hd__and2_1 _20879_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .X(_03977_));
 sky130_fd_sc_hd__a21boi_1 _20880_ (.A1(_03971_),
    .A2(_03973_),
    .B1_N(_03972_),
    .Y(_03978_));
 sky130_fd_sc_hd__or3_1 _20881_ (.A(_03976_),
    .B(_03977_),
    .C(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__o21ai_1 _20882_ (.A1(_03976_),
    .A2(_03977_),
    .B1(_03978_),
    .Y(_03980_));
 sky130_fd_sc_hd__a32o_1 _20883_ (.A1(_03948_),
    .A2(_03979_),
    .A3(_03980_),
    .B1(_02915_),
    .B2(\rbzero.texV[-5] ),
    .X(_01606_));
 sky130_fd_sc_hd__xnor2_1 _20884_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_03981_));
 sky130_fd_sc_hd__o21bai_1 _20885_ (.A1(_03976_),
    .A2(_03978_),
    .B1_N(_03977_),
    .Y(_03982_));
 sky130_fd_sc_hd__xnor2_1 _20886_ (.A(_03981_),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__a22o_1 _20887_ (.A1(\rbzero.texV[-4] ),
    .A2(_03567_),
    .B1(_03895_),
    .B2(_03983_),
    .X(_01607_));
 sky130_fd_sc_hd__nor2_1 _20888_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_1 _20889_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03985_));
 sky130_fd_sc_hd__and2b_1 _20890_ (.A_N(_03984_),
    .B(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__a21o_1 _20891_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_03982_),
    .X(_03987_));
 sky130_fd_sc_hd__o21ai_1 _20892_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__xnor2_1 _20893_ (.A(_03986_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__a22o_1 _20894_ (.A1(\rbzero.texV[-3] ),
    .A2(_03951_),
    .B1(_03895_),
    .B2(_03989_),
    .X(_01608_));
 sky130_fd_sc_hd__or2_1 _20895_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .X(_03990_));
 sky130_fd_sc_hd__nand2_1 _20896_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .Y(_03991_));
 sky130_fd_sc_hd__o21ai_2 _20897_ (.A1(_03984_),
    .A2(_03988_),
    .B1(_03985_),
    .Y(_03992_));
 sky130_fd_sc_hd__a21o_1 _20898_ (.A1(_03990_),
    .A2(_03991_),
    .B1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__nand3_1 _20899_ (.A(_03990_),
    .B(_03991_),
    .C(_03992_),
    .Y(_03994_));
 sky130_fd_sc_hd__a32o_1 _20900_ (.A1(_03948_),
    .A2(_03993_),
    .A3(_03994_),
    .B1(_02915_),
    .B2(\rbzero.texV[-2] ),
    .X(_01609_));
 sky130_fd_sc_hd__nor2_1 _20901_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .Y(_03995_));
 sky130_fd_sc_hd__and2_1 _20902_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .X(_03996_));
 sky130_fd_sc_hd__or2_1 _20903_ (.A(_03995_),
    .B(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__a21boi_1 _20904_ (.A1(_03990_),
    .A2(_03992_),
    .B1_N(_03991_),
    .Y(_03998_));
 sky130_fd_sc_hd__xor2_1 _20905_ (.A(_03997_),
    .B(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__a22o_1 _20906_ (.A1(\rbzero.texV[-1] ),
    .A2(_03951_),
    .B1(_03895_),
    .B2(_03999_),
    .X(_01610_));
 sky130_fd_sc_hd__nor2_1 _20907_ (.A(_03997_),
    .B(_03998_),
    .Y(_04000_));
 sky130_fd_sc_hd__or2_1 _20908_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .X(_04001_));
 sky130_fd_sc_hd__nand2_1 _20909_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .Y(_04002_));
 sky130_fd_sc_hd__o211a_1 _20910_ (.A1(_03996_),
    .A2(_04000_),
    .B1(_04001_),
    .C1(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__inv_2 _20911_ (.A(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__a211o_1 _20912_ (.A1(_04001_),
    .A2(_04002_),
    .B1(_03996_),
    .C1(_04000_),
    .X(_04005_));
 sky130_fd_sc_hd__a32o_1 _20913_ (.A1(_03948_),
    .A2(_04004_),
    .A3(_04005_),
    .B1(_02915_),
    .B2(\rbzero.texV[0] ),
    .X(_01611_));
 sky130_fd_sc_hd__or2_1 _20914_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .X(_04006_));
 sky130_fd_sc_hd__nand2_1 _20915_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .Y(_04007_));
 sky130_fd_sc_hd__nand2_1 _20916_ (.A(_04002_),
    .B(_04004_),
    .Y(_04008_));
 sky130_fd_sc_hd__a21o_1 _20917_ (.A1(_04006_),
    .A2(_04007_),
    .B1(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__and3_1 _20918_ (.A(_04006_),
    .B(_04007_),
    .C(_04008_),
    .X(_04010_));
 sky130_fd_sc_hd__inv_2 _20919_ (.A(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__a32o_1 _20920_ (.A1(_03948_),
    .A2(_04009_),
    .A3(_04011_),
    .B1(_02915_),
    .B2(\rbzero.texV[1] ),
    .X(_01612_));
 sky130_fd_sc_hd__or2_1 _20921_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .X(_04012_));
 sky130_fd_sc_hd__nand2_1 _20922_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .Y(_04013_));
 sky130_fd_sc_hd__nand2_1 _20923_ (.A(_04007_),
    .B(_04011_),
    .Y(_04014_));
 sky130_fd_sc_hd__and3_1 _20924_ (.A(_04012_),
    .B(_04013_),
    .C(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__inv_2 _20925_ (.A(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__a21o_1 _20926_ (.A1(_04012_),
    .A2(_04013_),
    .B1(_04014_),
    .X(_04017_));
 sky130_fd_sc_hd__a32o_1 _20927_ (.A1(_03948_),
    .A2(_04016_),
    .A3(_04017_),
    .B1(_02915_),
    .B2(\rbzero.texV[2] ),
    .X(_01613_));
 sky130_fd_sc_hd__or2_1 _20928_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .X(_04018_));
 sky130_fd_sc_hd__nand2_1 _20929_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .Y(_04019_));
 sky130_fd_sc_hd__nand2_1 _20930_ (.A(_04013_),
    .B(_04016_),
    .Y(_04020_));
 sky130_fd_sc_hd__a21o_1 _20931_ (.A1(_04018_),
    .A2(_04019_),
    .B1(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__and3_1 _20932_ (.A(_04018_),
    .B(_04019_),
    .C(_04020_),
    .X(_04022_));
 sky130_fd_sc_hd__inv_2 _20933_ (.A(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__a32o_1 _20934_ (.A1(_03948_),
    .A2(_04021_),
    .A3(_04023_),
    .B1(_02915_),
    .B2(\rbzero.texV[3] ),
    .X(_01614_));
 sky130_fd_sc_hd__or2_1 _20935_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .X(_04024_));
 sky130_fd_sc_hd__nand2_1 _20936_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_04025_));
 sky130_fd_sc_hd__nand2_1 _20937_ (.A(_04019_),
    .B(_04023_),
    .Y(_04026_));
 sky130_fd_sc_hd__a21o_1 _20938_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__nand3_1 _20939_ (.A(_04024_),
    .B(_04025_),
    .C(_04026_),
    .Y(_04028_));
 sky130_fd_sc_hd__a32o_1 _20940_ (.A1(_09870_),
    .A2(_04027_),
    .A3(_04028_),
    .B1(_02915_),
    .B2(\rbzero.texV[4] ),
    .X(_01615_));
 sky130_fd_sc_hd__a21boi_1 _20941_ (.A1(_04024_),
    .A2(_04026_),
    .B1_N(_04025_),
    .Y(_04029_));
 sky130_fd_sc_hd__nor2_1 _20942_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_1 _20943_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_04031_));
 sky130_fd_sc_hd__and2b_1 _20944_ (.A_N(_04030_),
    .B(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__xnor2_1 _20945_ (.A(_04029_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__a22o_1 _20946_ (.A1(\rbzero.texV[5] ),
    .A2(_03951_),
    .B1(_03895_),
    .B2(_04033_),
    .X(_01616_));
 sky130_fd_sc_hd__or2_1 _20947_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .X(_04034_));
 sky130_fd_sc_hd__nand2_1 _20948_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_1 _20949_ (.A(_04034_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__o21ai_1 _20950_ (.A1(_04029_),
    .A2(_04030_),
    .B1(_04031_),
    .Y(_04037_));
 sky130_fd_sc_hd__xnor2_1 _20951_ (.A(_04036_),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__a22o_1 _20952_ (.A1(\rbzero.texV[6] ),
    .A2(_03951_),
    .B1(_03895_),
    .B2(_04038_),
    .X(_01617_));
 sky130_fd_sc_hd__nor2_1 _20953_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_1 _20954_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_04040_));
 sky130_fd_sc_hd__and2b_1 _20955_ (.A_N(_04039_),
    .B(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__a21boi_1 _20956_ (.A1(_04034_),
    .A2(_04037_),
    .B1_N(_04035_),
    .Y(_04042_));
 sky130_fd_sc_hd__xnor2_1 _20957_ (.A(_04041_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__a22o_1 _20958_ (.A1(\rbzero.texV[7] ),
    .A2(_03951_),
    .B1(_03895_),
    .B2(_04043_),
    .X(_01618_));
 sky130_fd_sc_hd__or2_1 _20959_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .X(_04044_));
 sky130_fd_sc_hd__nand2_1 _20960_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_04045_));
 sky130_fd_sc_hd__o21ai_1 _20961_ (.A1(_04039_),
    .A2(_04042_),
    .B1(_04040_),
    .Y(_04046_));
 sky130_fd_sc_hd__a21o_1 _20962_ (.A1(_04044_),
    .A2(_04045_),
    .B1(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__nand3_1 _20963_ (.A(_04044_),
    .B(_04045_),
    .C(_04046_),
    .Y(_04048_));
 sky130_fd_sc_hd__a32o_1 _20964_ (.A1(_09870_),
    .A2(_04047_),
    .A3(_04048_),
    .B1(_02915_),
    .B2(\rbzero.texV[8] ),
    .X(_01619_));
 sky130_fd_sc_hd__or2_1 _20965_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .X(_04049_));
 sky130_fd_sc_hd__nand2_1 _20966_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_04050_));
 sky130_fd_sc_hd__a21o_1 _20967_ (.A1(\rbzero.traced_texa[8] ),
    .A2(\rbzero.texV[8] ),
    .B1(_04046_),
    .X(_04051_));
 sky130_fd_sc_hd__a22o_1 _20968_ (.A1(_04049_),
    .A2(_04050_),
    .B1(_04051_),
    .B2(_04044_),
    .X(_04052_));
 sky130_fd_sc_hd__nand4_1 _20969_ (.A(_04044_),
    .B(_04049_),
    .C(_04050_),
    .D(_04051_),
    .Y(_04053_));
 sky130_fd_sc_hd__a32o_1 _20970_ (.A1(_09870_),
    .A2(_04052_),
    .A3(_04053_),
    .B1(_02915_),
    .B2(\rbzero.texV[9] ),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_1 _20971_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_04054_));
 sky130_fd_sc_hd__and3_1 _20972_ (.A(_04050_),
    .B(_04053_),
    .C(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__a21oi_1 _20973_ (.A1(_04050_),
    .A2(_04053_),
    .B1(_04054_),
    .Y(_04056_));
 sky130_fd_sc_hd__nor2_1 _20974_ (.A(_04055_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__a22o_1 _20975_ (.A1(\rbzero.texV[10] ),
    .A2(_03951_),
    .B1(_03895_),
    .B2(_04057_),
    .X(_01621_));
 sky130_fd_sc_hd__nand2_1 _20976_ (.A(_04571_),
    .B(_09867_),
    .Y(_04058_));
 sky130_fd_sc_hd__a21o_1 _20977_ (.A1(_05173_),
    .A2(_04058_),
    .B1(_08165_),
    .X(_04059_));
 sky130_fd_sc_hd__inv_2 _20978_ (.A(_04059_),
    .Y(_04060_));
 sky130_fd_sc_hd__o211ai_1 _20979_ (.A1(_04570_),
    .A2(_08266_),
    .B1(_04060_),
    .C1(_04571_),
    .Y(_04061_));
 sky130_fd_sc_hd__o211a_1 _20980_ (.A1(_04571_),
    .A2(_04060_),
    .B1(_04061_),
    .C1(_04576_),
    .X(_01622_));
 sky130_fd_sc_hd__and3_1 _20981_ (.A(_04570_),
    .B(_04571_),
    .C(_04060_),
    .X(_04062_));
 sky130_fd_sc_hd__and3b_1 _20982_ (.A_N(_04062_),
    .B(_04576_),
    .C(_04564_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _20983_ (.A(_04063_),
    .X(_01623_));
 sky130_fd_sc_hd__a21oi_1 _20984_ (.A1(_04563_),
    .A2(_04062_),
    .B1(_08262_),
    .Y(_04064_));
 sky130_fd_sc_hd__o21a_1 _20985_ (.A1(_04563_),
    .A2(_04062_),
    .B1(_04064_),
    .X(_01624_));
 sky130_fd_sc_hd__a21boi_1 _20986_ (.A1(_04563_),
    .A2(_04570_),
    .B1_N(\rbzero.trace_state[3] ),
    .Y(_04065_));
 sky130_fd_sc_hd__o31a_1 _20987_ (.A1(_09069_),
    .A2(_04059_),
    .A3(_04065_),
    .B1(_01633_),
    .X(_01625_));
 sky130_fd_sc_hd__and2_2 _20988_ (.A(_03861_),
    .B(clknet_1_1__leaf__05795_),
    .X(_04066_));
 sky130_fd_sc_hd__buf_1 _20989_ (.A(_04066_),
    .X(_01626_));
 sky130_fd_sc_hd__and2_2 _20990_ (.A(_03861_),
    .B(clknet_1_0__leaf__05854_),
    .X(_04067_));
 sky130_fd_sc_hd__buf_1 _20991_ (.A(_04067_),
    .X(_01627_));
 sky130_fd_sc_hd__and2_2 _20992_ (.A(_03861_),
    .B(clknet_1_0__leaf__05916_),
    .X(_04068_));
 sky130_fd_sc_hd__buf_1 _20993_ (.A(_04068_),
    .X(_01628_));
 sky130_fd_sc_hd__and2_2 _20994_ (.A(_02808_),
    .B(clknet_1_1__leaf__05977_),
    .X(_04069_));
 sky130_fd_sc_hd__buf_1 _20995_ (.A(_04069_),
    .X(_01629_));
 sky130_fd_sc_hd__and2_2 _20996_ (.A(_02808_),
    .B(clknet_1_1__leaf__06036_),
    .X(_04070_));
 sky130_fd_sc_hd__buf_1 _20997_ (.A(_04070_),
    .X(_01630_));
 sky130_fd_sc_hd__and2_2 _20998_ (.A(_02808_),
    .B(clknet_1_0__leaf__06092_),
    .X(_04071_));
 sky130_fd_sc_hd__buf_1 _20999_ (.A(_04071_),
    .X(_01631_));
 sky130_fd_sc_hd__nor2_1 _21000_ (.A(\rbzero.hsync ),
    .B(net64),
    .Y(_01632_));
 sky130_fd_sc_hd__a22o_1 _21001_ (.A1(\rbzero.traced_texVinit[0] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(_09257_),
    .X(_01634_));
 sky130_fd_sc_hd__a22o_1 _21002_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(_09253_),
    .X(_01635_));
 sky130_fd_sc_hd__a22o_1 _21003_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(_09249_),
    .X(_01636_));
 sky130_fd_sc_hd__a22o_1 _21004_ (.A1(\rbzero.traced_texVinit[3] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(_09366_),
    .X(_01637_));
 sky130_fd_sc_hd__a22o_1 _21005_ (.A1(\rbzero.traced_texVinit[4] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(_09487_),
    .X(_01638_));
 sky130_fd_sc_hd__a22o_1 _21006_ (.A1(\rbzero.traced_texVinit[5] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(_10009_),
    .X(_01639_));
 sky130_fd_sc_hd__a22o_1 _21007_ (.A1(\rbzero.traced_texVinit[6] ),
    .A2(_09894_),
    .B1(_09895_),
    .B2(_09738_),
    .X(_01640_));
 sky130_fd_sc_hd__buf_6 _21008_ (.A(_09881_),
    .X(_04072_));
 sky130_fd_sc_hd__a22o_1 _21009_ (.A1(\rbzero.traced_texVinit[7] ),
    .A2(_04072_),
    .B1(_09895_),
    .B2(_09859_),
    .X(_01641_));
 sky130_fd_sc_hd__a22o_1 _21010_ (.A1(\rbzero.traced_texVinit[8] ),
    .A2(_04072_),
    .B1(_09895_),
    .B2(_10152_),
    .X(_01642_));
 sky130_fd_sc_hd__a22o_1 _21011_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_10268_),
    .X(_01643_));
 sky130_fd_sc_hd__a22o_1 _21012_ (.A1(\rbzero.traced_texVinit[10] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_10390_),
    .X(_01644_));
 sky130_fd_sc_hd__nor2_1 _21013_ (.A(\gpout0.clk_div[0] ),
    .B(net64),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _21014_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .Y(_04073_));
 sky130_fd_sc_hd__or2_1 _21015_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .X(_04074_));
 sky130_fd_sc_hd__and3_1 _21016_ (.A(_02850_),
    .B(_04073_),
    .C(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__clkbuf_1 _21017_ (.A(_04075_),
    .X(_01646_));
 sky130_fd_sc_hd__or2_1 _21018_ (.A(_02538_),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_04076_));
 sky130_fd_sc_hd__and3_1 _21019_ (.A(_09884_),
    .B(_02528_),
    .C(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__a21o_1 _21020_ (.A1(\rbzero.wall_tracer.rayAddendX[-9] ),
    .A2(_09882_),
    .B1(_04077_),
    .X(_01647_));
 sky130_fd_sc_hd__xor2_1 _21021_ (.A(_02528_),
    .B(_02531_),
    .X(_04078_));
 sky130_fd_sc_hd__a22o_1 _21022_ (.A1(\rbzero.wall_tracer.rayAddendX[-8] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_04078_),
    .X(_01648_));
 sky130_fd_sc_hd__and2b_1 _21023_ (.A_N(_02527_),
    .B(_02533_),
    .X(_04079_));
 sky130_fd_sc_hd__xnor2_1 _21024_ (.A(_02532_),
    .B(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__a22o_1 _21025_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_04080_),
    .X(_01649_));
 sky130_fd_sc_hd__xnor2_1 _21026_ (.A(_02526_),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .Y(_04081_));
 sky130_fd_sc_hd__xnor2_1 _21027_ (.A(_02534_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__a22o_1 _21028_ (.A1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_04082_),
    .X(_01650_));
 sky130_fd_sc_hd__or2_1 _21029_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_04083_));
 sky130_fd_sc_hd__and3_1 _21030_ (.A(_09884_),
    .B(_03234_),
    .C(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__a21o_1 _21031_ (.A1(\rbzero.wall_tracer.rayAddendY[-9] ),
    .A2(_09882_),
    .B1(_04084_),
    .X(_01651_));
 sky130_fd_sc_hd__nor2_1 _21032_ (.A(_03236_),
    .B(_03235_),
    .Y(_04085_));
 sky130_fd_sc_hd__xnor2_1 _21033_ (.A(_03234_),
    .B(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__a22o_1 _21034_ (.A1(\rbzero.wall_tracer.rayAddendY[-8] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_04086_),
    .X(_01652_));
 sky130_fd_sc_hd__and2b_1 _21035_ (.A_N(_03233_),
    .B(_03238_),
    .X(_04087_));
 sky130_fd_sc_hd__xnor2_1 _21036_ (.A(_03237_),
    .B(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__a22o_1 _21037_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_04088_),
    .X(_01653_));
 sky130_fd_sc_hd__xnor2_1 _21038_ (.A(_03232_),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .Y(_04089_));
 sky130_fd_sc_hd__xnor2_1 _21039_ (.A(_03239_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__a22o_1 _21040_ (.A1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .A2(_04072_),
    .B1(_02571_),
    .B2(_04090_),
    .X(_01654_));
 sky130_fd_sc_hd__nor2_1 _21041_ (.A(\gpout1.clk_div[0] ),
    .B(net64),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_1 _21042_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .Y(_04091_));
 sky130_fd_sc_hd__or2_1 _21043_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .X(_04092_));
 sky130_fd_sc_hd__and3_1 _21044_ (.A(_02876_),
    .B(_04091_),
    .C(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__clkbuf_1 _21045_ (.A(_04093_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_1 _21046_ (.A(\gpout2.clk_div[0] ),
    .B(net64),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _21047_ (.A(\gpout2.clk_div[1] ),
    .B(\gpout2.clk_div[0] ),
    .Y(_04094_));
 sky130_fd_sc_hd__or2_1 _21048_ (.A(\gpout2.clk_div[1] ),
    .B(\gpout2.clk_div[0] ),
    .X(_04095_));
 sky130_fd_sc_hd__and3_1 _21049_ (.A(_02876_),
    .B(_04094_),
    .C(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _21050_ (.A(_04096_),
    .X(_01658_));
 sky130_fd_sc_hd__nor2_1 _21051_ (.A(\gpout3.clk_div[0] ),
    .B(net64),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _21052_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .Y(_04097_));
 sky130_fd_sc_hd__or2_1 _21053_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .X(_04098_));
 sky130_fd_sc_hd__and3_1 _21054_ (.A(_02876_),
    .B(_04097_),
    .C(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__clkbuf_1 _21055_ (.A(_04099_),
    .X(_01660_));
 sky130_fd_sc_hd__nor2_1 _21056_ (.A(\gpout4.clk_div[0] ),
    .B(net64),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _21057_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .Y(_04100_));
 sky130_fd_sc_hd__or2_1 _21058_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .X(_04101_));
 sky130_fd_sc_hd__and3_1 _21059_ (.A(_02876_),
    .B(_04100_),
    .C(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__clkbuf_1 _21060_ (.A(_04102_),
    .X(_01662_));
 sky130_fd_sc_hd__dfxtp_2 _21061_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00000_),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21062_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00001_),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00386_),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00387_),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00388_),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00389_),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00390_),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21068_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00391_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00392_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00393_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21071_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00394_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00395_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21073_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00396_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21074_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00397_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00398_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00399_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00400_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00401_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00402_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21080_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00403_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21081_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00404_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00405_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21088_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00413_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_4 _21091_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00414_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _21092_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00415_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21093_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00416_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00417_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00418_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00419_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21097_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00420_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21098_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00421_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21099_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00422_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21100_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00423_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21101_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00424_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_4 _21102_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00425_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_4 _21103_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00426_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21104_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00427_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_4 _21105_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00428_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_4 _21106_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00429_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21107_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00430_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_4 _21108_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00431_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_4 _21109_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00432_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_4 _21110_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00433_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_4 _21111_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00434_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21112_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21113_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21114_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21115_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21116_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21117_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21118_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21119_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21120_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21122_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21125_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21127_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21128_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21129_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21130_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21131_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21133_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21134_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00457_),
    .Q(\reg_rgb[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21135_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00458_),
    .Q(\reg_rgb[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21136_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00459_),
    .Q(\reg_rgb[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00460_),
    .Q(\reg_rgb[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21138_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00461_),
    .Q(\reg_rgb[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21139_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00462_),
    .Q(\reg_rgb[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21140_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00463_),
    .Q(\rbzero.wall_hot[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21141_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00464_),
    .Q(\rbzero.wall_hot[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21142_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00465_),
    .Q(\rbzero.side_hot ));
 sky130_fd_sc_hd__dfxtp_1 _21143_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00466_),
    .Q(\rbzero.texu_hot[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21144_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00467_),
    .Q(\rbzero.texu_hot[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21145_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00468_),
    .Q(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21146_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00469_),
    .Q(\rbzero.texu_hot[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21147_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00470_),
    .Q(\rbzero.texu_hot[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21148_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00471_),
    .Q(\rbzero.texu_hot[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21149_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00472_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21150_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00473_),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21151_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00474_),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21152_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00475_),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21153_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00476_),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21154_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00477_),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21155_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00478_),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21156_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00479_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21157_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00480_),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_4 _21158_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00481_),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_4 _21159_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00482_),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00483_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00484_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21162_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00485_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21163_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00486_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21164_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00487_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00488_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21166_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00489_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00490_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00491_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00492_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00493_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21171_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00494_),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00495_),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21173_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00496_),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00497_),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21175_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00498_),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21176_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00499_),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21177_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00500_),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00501_),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00502_),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00503_),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00504_),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21182_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00505_),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00506_),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21184_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00507_),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00508_),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00509_),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00510_),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00511_),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21189_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00512_),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00513_),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00514_),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00515_),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00516_),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00517_),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21195_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00518_),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21196_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00519_),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00520_),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21198_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00521_),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00522_),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00523_),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00524_),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00525_),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00526_),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00527_),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21205_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00528_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21206_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00529_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00530_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00531_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21209_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00532_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21210_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00533_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00534_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21212_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00535_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00536_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21214_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00537_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21215_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00538_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21216_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00539_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00540_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21220_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21225_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21226_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21227_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21245_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21247_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21248_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00572_),
    .Q(\rbzero.spi_registers.new_texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00573_),
    .Q(\rbzero.spi_registers.new_texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00574_),
    .Q(\rbzero.spi_registers.new_texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00575_),
    .Q(\rbzero.spi_registers.new_texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00576_),
    .Q(\rbzero.spi_registers.new_texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00577_),
    .Q(\rbzero.spi_registers.new_texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00578_),
    .Q(\rbzero.spi_registers.new_texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00579_),
    .Q(\rbzero.spi_registers.new_texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00580_),
    .Q(\rbzero.spi_registers.new_texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21258_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00581_),
    .Q(\rbzero.spi_registers.new_texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21259_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00582_),
    .Q(\rbzero.spi_registers.new_texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21260_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00583_),
    .Q(\rbzero.spi_registers.new_texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21261_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00584_),
    .Q(\rbzero.spi_registers.new_texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21262_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00585_),
    .Q(\rbzero.spi_registers.new_texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00586_),
    .Q(\rbzero.spi_registers.new_texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21264_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00587_),
    .Q(\rbzero.spi_registers.new_texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00588_),
    .Q(\rbzero.spi_registers.new_texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00589_),
    .Q(\rbzero.spi_registers.new_texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21267_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00590_),
    .Q(\rbzero.spi_registers.new_texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00591_),
    .Q(\rbzero.spi_registers.new_texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21269_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00592_),
    .Q(\rbzero.spi_registers.new_texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00593_),
    .Q(\rbzero.spi_registers.new_texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00594_),
    .Q(\rbzero.spi_registers.new_texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00595_),
    .Q(\rbzero.spi_registers.new_texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00596_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00597_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21275_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00598_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21276_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00599_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21277_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00600_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21278_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00601_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00602_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21280_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00603_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00604_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21282_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00605_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00606_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21284_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00607_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00608_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00609_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00610_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00611_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00612_),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_4 _21290_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00613_),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_2 _21291_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00614_),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_2 _21292_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00615_),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_4 _21293_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00616_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21294_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00617_),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00618_),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00619_),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_1 _21297_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00620_),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00621_),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_4 _21299_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00622_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00623_),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21301_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00624_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00625_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21303_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00626_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00627_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00628_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00629_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00630_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00631_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21309_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00632_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21310_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00633_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00634_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00635_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00636_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00637_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00638_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00639_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21317_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00640_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21318_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00641_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21319_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00642_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21320_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00643_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21321_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00644_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21322_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00645_),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _21323_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00646_),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21324_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00647_),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _21325_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00648_),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _21326_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00649_),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00650_),
    .Q(\rbzero.spi_registers.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00651_),
    .Q(\rbzero.spi_registers.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00652_),
    .Q(\rbzero.spi_registers.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00653_),
    .Q(\rbzero.spi_registers.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00654_),
    .Q(\rbzero.spi_registers.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00655_),
    .Q(\rbzero.spi_registers.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00656_),
    .Q(\rbzero.spi_registers.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00657_),
    .Q(\rbzero.spi_registers.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_2 _21335_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00658_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00659_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00660_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00661_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00662_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00663_),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00664_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00665_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00666_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00667_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00668_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00669_),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00670_),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00671_),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00672_),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00673_),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00674_),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00675_),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00676_),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00677_),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00678_),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21356_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00679_),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00680_),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00681_),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00682_),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00683_),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00684_),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00685_),
    .Q(\rbzero.map_overlay.i_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00686_),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00687_),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00688_),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00689_),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00690_),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00691_),
    .Q(\rbzero.map_overlay.i_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00692_),
    .Q(\rbzero.mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00693_),
    .Q(\rbzero.mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00694_),
    .Q(\rbzero.mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00695_),
    .Q(\rbzero.mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00696_),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00697_),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00698_),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00699_),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00700_),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00701_),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00702_),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00703_),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00704_),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00705_),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00706_),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00707_),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00708_),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00709_),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00710_),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00711_),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00712_),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00713_),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00714_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00715_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00716_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00717_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00718_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00719_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00720_),
    .Q(\rbzero.spi_registers.texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00721_),
    .Q(\rbzero.spi_registers.texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00722_),
    .Q(\rbzero.spi_registers.texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00723_),
    .Q(\rbzero.spi_registers.texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00724_),
    .Q(\rbzero.spi_registers.texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00725_),
    .Q(\rbzero.spi_registers.texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00726_),
    .Q(\rbzero.spi_registers.texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00727_),
    .Q(\rbzero.spi_registers.texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00728_),
    .Q(\rbzero.spi_registers.texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00729_),
    .Q(\rbzero.spi_registers.texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00730_),
    .Q(\rbzero.spi_registers.texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00731_),
    .Q(\rbzero.spi_registers.texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21409_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00732_),
    .Q(\rbzero.spi_registers.texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21410_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00733_),
    .Q(\rbzero.spi_registers.texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21411_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00734_),
    .Q(\rbzero.spi_registers.texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21412_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00735_),
    .Q(\rbzero.spi_registers.texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21413_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00736_),
    .Q(\rbzero.spi_registers.texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00737_),
    .Q(\rbzero.spi_registers.texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00738_),
    .Q(\rbzero.spi_registers.texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21416_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00739_),
    .Q(\rbzero.spi_registers.texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00740_),
    .Q(\rbzero.spi_registers.texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00741_),
    .Q(\rbzero.spi_registers.texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21419_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00742_),
    .Q(\rbzero.spi_registers.texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00743_),
    .Q(\rbzero.spi_registers.texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00744_),
    .Q(\rbzero.spi_registers.texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00745_),
    .Q(\rbzero.spi_registers.texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00746_),
    .Q(\rbzero.spi_registers.texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21424_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00747_),
    .Q(\rbzero.spi_registers.texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21425_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00748_),
    .Q(\rbzero.spi_registers.texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00749_),
    .Q(\rbzero.spi_registers.texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00750_),
    .Q(\rbzero.spi_registers.texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00751_),
    .Q(\rbzero.spi_registers.texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00752_),
    .Q(\rbzero.spi_registers.texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00753_),
    .Q(\rbzero.spi_registers.texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21431_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00754_),
    .Q(\rbzero.spi_registers.texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21432_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00755_),
    .Q(\rbzero.spi_registers.texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21433_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00756_),
    .Q(\rbzero.spi_registers.texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21434_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00757_),
    .Q(\rbzero.spi_registers.texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00758_),
    .Q(\rbzero.spi_registers.texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21436_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00759_),
    .Q(\rbzero.spi_registers.texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21437_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00760_),
    .Q(\rbzero.spi_registers.texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21438_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00761_),
    .Q(\rbzero.spi_registers.texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00762_),
    .Q(\rbzero.spi_registers.texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21440_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00763_),
    .Q(\rbzero.spi_registers.texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21441_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00764_),
    .Q(\rbzero.spi_registers.texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00765_),
    .Q(\rbzero.spi_registers.texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00766_),
    .Q(\rbzero.spi_registers.texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00767_),
    .Q(\rbzero.spi_registers.texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00768_),
    .Q(\rbzero.spi_registers.texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00769_),
    .Q(\rbzero.spi_registers.texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21447_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00770_),
    .Q(\rbzero.spi_registers.texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00771_),
    .Q(\rbzero.spi_registers.texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00772_),
    .Q(\rbzero.spi_registers.texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21450_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00773_),
    .Q(\rbzero.spi_registers.texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00774_),
    .Q(\rbzero.spi_registers.texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00775_),
    .Q(\rbzero.spi_registers.texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00776_),
    .Q(\rbzero.spi_registers.texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00777_),
    .Q(\rbzero.spi_registers.texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00778_),
    .Q(\rbzero.spi_registers.texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00779_),
    .Q(\rbzero.spi_registers.texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00780_),
    .Q(\rbzero.spi_registers.texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00781_),
    .Q(\rbzero.spi_registers.texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00782_),
    .Q(\rbzero.spi_registers.texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21460_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00783_),
    .Q(\rbzero.spi_registers.texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21461_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00784_),
    .Q(\rbzero.spi_registers.texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21462_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00785_),
    .Q(\rbzero.spi_registers.texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21463_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00786_),
    .Q(\rbzero.spi_registers.texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00787_),
    .Q(\rbzero.spi_registers.texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21465_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00788_),
    .Q(\rbzero.spi_registers.texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00789_),
    .Q(\rbzero.spi_registers.texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00790_),
    .Q(\rbzero.spi_registers.texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21468_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00791_),
    .Q(\rbzero.spi_registers.texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21469_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00792_),
    .Q(\rbzero.spi_registers.texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21470_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00793_),
    .Q(\rbzero.spi_registers.texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00794_),
    .Q(\rbzero.spi_registers.texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21472_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00795_),
    .Q(\rbzero.spi_registers.texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21473_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00796_),
    .Q(\rbzero.spi_registers.texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21474_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00797_),
    .Q(\rbzero.spi_registers.texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00798_),
    .Q(\rbzero.spi_registers.texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21476_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00799_),
    .Q(\rbzero.spi_registers.texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00800_),
    .Q(\rbzero.spi_registers.texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00801_),
    .Q(\rbzero.spi_registers.texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00802_),
    .Q(\rbzero.spi_registers.texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00803_),
    .Q(\rbzero.spi_registers.texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00804_),
    .Q(\rbzero.spi_registers.texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00805_),
    .Q(\rbzero.spi_registers.texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21483_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00806_),
    .Q(\rbzero.spi_registers.texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00807_),
    .Q(\rbzero.spi_registers.texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00808_),
    .Q(\rbzero.spi_registers.texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21486_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00809_),
    .Q(\rbzero.spi_registers.texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00810_),
    .Q(\rbzero.spi_registers.texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21488_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00811_),
    .Q(\rbzero.spi_registers.texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21489_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00812_),
    .Q(\rbzero.spi_registers.texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21490_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00813_),
    .Q(\rbzero.spi_registers.texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21491_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00814_),
    .Q(\rbzero.spi_registers.texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21492_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00815_),
    .Q(\rbzero.spi_registers.texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21493_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00816_),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00817_),
    .Q(\rbzero.spi_registers.new_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21495_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00818_),
    .Q(\rbzero.spi_registers.new_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21496_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00819_),
    .Q(\rbzero.spi_registers.new_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21497_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00820_),
    .Q(\rbzero.spi_registers.new_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21498_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00821_),
    .Q(\rbzero.spi_registers.new_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21499_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00822_),
    .Q(\rbzero.spi_registers.new_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21500_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00823_),
    .Q(\rbzero.spi_registers.got_new_sky ));
 sky130_fd_sc_hd__dfxtp_1 _21501_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00824_),
    .Q(\rbzero.spi_registers.new_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21502_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00825_),
    .Q(\rbzero.spi_registers.new_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21503_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00826_),
    .Q(\rbzero.spi_registers.new_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21504_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00827_),
    .Q(\rbzero.spi_registers.new_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00828_),
    .Q(\rbzero.spi_registers.new_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21506_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00829_),
    .Q(\rbzero.spi_registers.new_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00830_),
    .Q(\rbzero.spi_registers.got_new_floor ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00831_),
    .Q(\rbzero.spi_registers.new_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00832_),
    .Q(\rbzero.spi_registers.new_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21510_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00833_),
    .Q(\rbzero.spi_registers.new_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21511_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00834_),
    .Q(\rbzero.spi_registers.new_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21512_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00835_),
    .Q(\rbzero.spi_registers.new_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21513_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00836_),
    .Q(\rbzero.spi_registers.new_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21514_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00837_),
    .Q(\rbzero.spi_registers.got_new_leak ));
 sky130_fd_sc_hd__dfxtp_1 _21515_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00838_),
    .Q(\rbzero.spi_registers.new_other[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21516_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00839_),
    .Q(\rbzero.spi_registers.new_other[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21517_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00840_),
    .Q(\rbzero.spi_registers.new_other[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21518_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00841_),
    .Q(\rbzero.spi_registers.new_other[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00842_),
    .Q(\rbzero.spi_registers.new_other[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00843_),
    .Q(\rbzero.spi_registers.new_other[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21521_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00844_),
    .Q(\rbzero.spi_registers.new_other[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21522_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00845_),
    .Q(\rbzero.spi_registers.new_other[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21523_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00846_),
    .Q(\rbzero.spi_registers.new_other[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21524_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00847_),
    .Q(\rbzero.spi_registers.new_other[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00848_),
    .Q(\rbzero.spi_registers.got_new_other ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00849_),
    .Q(\rbzero.spi_registers.new_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00850_),
    .Q(\rbzero.spi_registers.new_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21528_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00851_),
    .Q(\rbzero.spi_registers.new_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21529_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00852_),
    .Q(\rbzero.spi_registers.new_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00853_),
    .Q(\rbzero.spi_registers.new_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21531_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00854_),
    .Q(\rbzero.spi_registers.new_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21532_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00855_),
    .Q(\rbzero.spi_registers.got_new_vshift ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00856_),
    .Q(\rbzero.spi_registers.new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21534_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00857_),
    .Q(\rbzero.spi_registers.got_new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21535_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00858_),
    .Q(\rbzero.spi_registers.new_mapd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00859_),
    .Q(\rbzero.spi_registers.new_mapd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21537_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00860_),
    .Q(\rbzero.spi_registers.new_mapd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00861_),
    .Q(\rbzero.spi_registers.new_mapd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21539_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00862_),
    .Q(\rbzero.spi_registers.new_mapd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00863_),
    .Q(\rbzero.spi_registers.new_mapd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21541_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00864_),
    .Q(\rbzero.spi_registers.new_mapd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21542_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00865_),
    .Q(\rbzero.spi_registers.new_mapd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21543_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00866_),
    .Q(\rbzero.spi_registers.new_mapd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00867_),
    .Q(\rbzero.spi_registers.new_mapd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21545_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00868_),
    .Q(\rbzero.spi_registers.new_mapd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21546_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00869_),
    .Q(\rbzero.spi_registers.new_mapd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00870_),
    .Q(\rbzero.spi_registers.new_mapd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21548_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00871_),
    .Q(\rbzero.spi_registers.new_mapd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00872_),
    .Q(\rbzero.spi_registers.new_mapd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21550_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00873_),
    .Q(\rbzero.spi_registers.new_mapd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00874_),
    .Q(\rbzero.spi_registers.got_new_mapd ));
 sky130_fd_sc_hd__dfxtp_1 _21552_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00875_),
    .Q(\rbzero.spi_registers.new_texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21553_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00876_),
    .Q(\rbzero.spi_registers.new_texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21554_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00877_),
    .Q(\rbzero.spi_registers.new_texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00878_),
    .Q(\rbzero.spi_registers.new_texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21556_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00879_),
    .Q(\rbzero.spi_registers.new_texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21557_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00880_),
    .Q(\rbzero.spi_registers.new_texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21558_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00881_),
    .Q(\rbzero.spi_registers.new_texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21559_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00882_),
    .Q(\rbzero.spi_registers.new_texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00883_),
    .Q(\rbzero.spi_registers.new_texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00884_),
    .Q(\rbzero.spi_registers.new_texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00885_),
    .Q(\rbzero.spi_registers.new_texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00886_),
    .Q(\rbzero.spi_registers.new_texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00887_),
    .Q(\rbzero.spi_registers.new_texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00888_),
    .Q(\rbzero.spi_registers.new_texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21566_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00889_),
    .Q(\rbzero.spi_registers.new_texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00890_),
    .Q(\rbzero.spi_registers.new_texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21568_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00891_),
    .Q(\rbzero.spi_registers.new_texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00892_),
    .Q(\rbzero.spi_registers.new_texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00893_),
    .Q(\rbzero.spi_registers.new_texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00894_),
    .Q(\rbzero.spi_registers.new_texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21572_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00895_),
    .Q(\rbzero.spi_registers.new_texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00896_),
    .Q(\rbzero.spi_registers.new_texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00897_),
    .Q(\rbzero.spi_registers.new_texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00898_),
    .Q(\rbzero.spi_registers.new_texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00899_),
    .Q(\rbzero.spi_registers.got_new_texadd0 ));
 sky130_fd_sc_hd__dfxtp_1 _21577_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00900_),
    .Q(\rbzero.spi_registers.new_texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21578_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00901_),
    .Q(\rbzero.spi_registers.new_texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21579_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00902_),
    .Q(\rbzero.spi_registers.new_texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00903_),
    .Q(\rbzero.spi_registers.new_texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21581_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00904_),
    .Q(\rbzero.spi_registers.new_texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21582_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00905_),
    .Q(\rbzero.spi_registers.new_texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00906_),
    .Q(\rbzero.spi_registers.new_texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21584_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00907_),
    .Q(\rbzero.spi_registers.new_texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21585_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00908_),
    .Q(\rbzero.spi_registers.new_texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21586_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00909_),
    .Q(\rbzero.spi_registers.new_texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21587_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00910_),
    .Q(\rbzero.spi_registers.new_texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21588_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00911_),
    .Q(\rbzero.spi_registers.new_texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21589_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00912_),
    .Q(\rbzero.spi_registers.new_texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21590_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00913_),
    .Q(\rbzero.spi_registers.new_texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21591_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00914_),
    .Q(\rbzero.spi_registers.new_texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00915_),
    .Q(\rbzero.spi_registers.new_texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21593_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00916_),
    .Q(\rbzero.spi_registers.new_texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21594_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00917_),
    .Q(\rbzero.spi_registers.new_texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00918_),
    .Q(\rbzero.spi_registers.new_texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21596_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00919_),
    .Q(\rbzero.spi_registers.new_texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21597_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00920_),
    .Q(\rbzero.spi_registers.new_texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00921_),
    .Q(\rbzero.spi_registers.new_texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21599_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00922_),
    .Q(\rbzero.spi_registers.new_texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21600_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00923_),
    .Q(\rbzero.spi_registers.new_texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21601_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00924_),
    .Q(\rbzero.spi_registers.got_new_texadd1 ));
 sky130_fd_sc_hd__dfxtp_1 _21602_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00925_),
    .Q(\rbzero.spi_registers.new_texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21603_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00926_),
    .Q(\rbzero.spi_registers.new_texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21604_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00927_),
    .Q(\rbzero.spi_registers.new_texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21605_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00928_),
    .Q(\rbzero.spi_registers.new_texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21606_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00929_),
    .Q(\rbzero.spi_registers.new_texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00930_),
    .Q(\rbzero.spi_registers.new_texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00931_),
    .Q(\rbzero.spi_registers.new_texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21609_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00932_),
    .Q(\rbzero.spi_registers.new_texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00933_),
    .Q(\rbzero.spi_registers.new_texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00934_),
    .Q(\rbzero.spi_registers.new_texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00935_),
    .Q(\rbzero.spi_registers.new_texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00936_),
    .Q(\rbzero.spi_registers.new_texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21614_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00937_),
    .Q(\rbzero.spi_registers.new_texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00938_),
    .Q(\rbzero.spi_registers.new_texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00939_),
    .Q(\rbzero.spi_registers.new_texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00940_),
    .Q(\rbzero.spi_registers.new_texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21618_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00941_),
    .Q(\rbzero.spi_registers.new_texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21619_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00942_),
    .Q(\rbzero.spi_registers.new_texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00943_),
    .Q(\rbzero.spi_registers.new_texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00944_),
    .Q(\rbzero.spi_registers.new_texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00945_),
    .Q(\rbzero.spi_registers.new_texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00946_),
    .Q(\rbzero.spi_registers.new_texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00947_),
    .Q(\rbzero.spi_registers.new_texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00948_),
    .Q(\rbzero.spi_registers.new_texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21626_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00949_),
    .Q(\rbzero.spi_registers.got_new_texadd2 ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00950_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00951_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21629_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00952_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21630_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00953_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21631_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00954_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21632_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00955_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00956_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21634_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00957_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21635_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00958_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21636_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00959_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21637_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00960_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21638_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00961_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00962_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21640_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00963_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21641_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00964_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21642_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00965_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21643_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00966_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00967_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_4 _21645_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00968_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21646_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00969_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21647_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00970_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21648_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00971_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21649_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00972_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21650_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00973_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21651_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00974_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _21652_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00975_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21653_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00976_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_4 _21654_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00977_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_4 _21655_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00978_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21656_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00979_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21657_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00980_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_4 _21658_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00981_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21659_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00982_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00983_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00984_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00985_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00986_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21664_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00987_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00988_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21666_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00989_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_4 _21667_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00990_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21668_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00991_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21669_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00992_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21670_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00993_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21671_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00994_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21672_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00995_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21673_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00996_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21674_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00997_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21675_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00998_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00999_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21677_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01000_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01001_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01002_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01003_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01004_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21682_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01005_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01006_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01007_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21685_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01008_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21686_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01009_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21687_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01010_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01011_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21689_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01012_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21690_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01013_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21691_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01014_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01015_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21693_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01016_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21694_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01017_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21695_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01018_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21696_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01019_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01020_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21698_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01021_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21699_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01022_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01023_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01024_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21702_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01025_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21703_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01026_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21704_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01027_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21705_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01028_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21706_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01029_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21707_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01030_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21708_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01031_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21709_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01032_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21710_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01033_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21711_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01034_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21712_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01035_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_4 _21713_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01036_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21714_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01037_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21715_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01038_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _21716_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01039_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21717_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01040_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21718_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01041_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21719_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01042_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21720_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01043_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21721_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01044_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21722_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01045_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21723_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01046_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21724_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01047_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21725_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01048_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21726_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01049_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21727_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01050_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01051_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01052_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01053_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21731_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01054_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21732_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01055_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21733_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01056_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21734_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01057_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21735_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01058_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21736_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01059_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21737_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01060_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21738_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01061_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21739_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01062_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21740_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01063_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21741_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01064_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21742_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01065_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21743_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01066_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21744_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01067_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21745_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01068_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21746_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01069_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21747_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01070_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21748_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01071_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21749_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01072_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21750_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01073_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21751_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01074_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21752_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01075_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21753_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01076_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21754_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01077_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21755_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01078_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21756_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01079_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21757_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01080_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21758_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01081_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21759_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01082_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01083_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01084_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21762_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01085_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21763_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01086_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21764_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01087_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21765_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01088_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21766_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01089_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21767_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01090_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21768_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01091_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21769_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01092_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21770_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01093_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21771_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01094_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21772_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01095_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21773_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01096_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01097_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21775_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01098_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21776_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01099_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21777_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01100_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21778_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01101_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21779_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01102_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01103_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21781_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01104_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21782_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01105_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21783_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01106_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21784_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01107_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01108_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21786_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01109_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21787_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01110_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21788_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01111_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21789_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01112_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21790_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01113_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21791_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01114_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21792_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01115_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21793_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01116_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21794_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01117_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21795_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01118_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21796_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01119_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01120_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21798_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01121_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21799_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01122_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21800_ (.CLK(net153),
    .D(_01123_),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(net154),
    .D(_01124_),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21802_ (.CLK(net155),
    .D(_01125_),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21803_ (.CLK(net156),
    .D(_01126_),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21804_ (.CLK(net157),
    .D(_01127_),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(net158),
    .D(_01128_),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(net159),
    .D(_01129_),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21807_ (.CLK(net160),
    .D(_01130_),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(net161),
    .D(_01131_),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(net162),
    .D(_01132_),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(net163),
    .D(_01133_),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(net164),
    .D(_01134_),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(net165),
    .D(_01135_),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(net166),
    .D(_01136_),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(net167),
    .D(_01137_),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21815_ (.CLK(net168),
    .D(_01138_),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21816_ (.CLK(net169),
    .D(_01139_),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21817_ (.CLK(net170),
    .D(_01140_),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(net171),
    .D(_01141_),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21819_ (.CLK(net172),
    .D(_01142_),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21820_ (.CLK(net173),
    .D(_01143_),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(net174),
    .D(_01144_),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21822_ (.CLK(net175),
    .D(_01145_),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21823_ (.CLK(net176),
    .D(_01146_),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21824_ (.CLK(net177),
    .D(_01147_),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21825_ (.CLK(net178),
    .D(_01148_),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21826_ (.CLK(net179),
    .D(_01149_),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21827_ (.CLK(net180),
    .D(_01150_),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21828_ (.CLK(net181),
    .D(_01151_),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21829_ (.CLK(net182),
    .D(_01152_),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21830_ (.CLK(net183),
    .D(_01153_),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21831_ (.CLK(net184),
    .D(_01154_),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21832_ (.CLK(net185),
    .D(_01155_),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21833_ (.CLK(net186),
    .D(_01156_),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(net187),
    .D(_01157_),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(net188),
    .D(_01158_),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(net189),
    .D(_01159_),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(net190),
    .D(_01160_),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(net191),
    .D(_01161_),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21839_ (.CLK(net192),
    .D(_01162_),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(net193),
    .D(_01163_),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21841_ (.CLK(net194),
    .D(_01164_),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21842_ (.CLK(net195),
    .D(_01165_),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21843_ (.CLK(net196),
    .D(_01166_),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21844_ (.CLK(net197),
    .D(_01167_),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(net198),
    .D(_01168_),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21846_ (.CLK(net199),
    .D(_01169_),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21847_ (.CLK(net200),
    .D(_01170_),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21848_ (.CLK(net201),
    .D(_01171_),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(net202),
    .D(_01172_),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(net203),
    .D(_01173_),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(net204),
    .D(_01174_),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(net205),
    .D(_01175_),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21853_ (.CLK(net206),
    .D(_01176_),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(net207),
    .D(_01177_),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(net208),
    .D(_01178_),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(net209),
    .D(_01179_),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(net210),
    .D(_01180_),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(net211),
    .D(_01181_),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(net212),
    .D(_01182_),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(net213),
    .D(_01183_),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(net214),
    .D(_01184_),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(net215),
    .D(_01185_),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21863_ (.CLK(net216),
    .D(_01186_),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01187_),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01188_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01189_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01190_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01191_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01192_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01193_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01194_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01195_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21873_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01196_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21874_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01197_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01198_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01199_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01200_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21878_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01201_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21879_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01202_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21880_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01203_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01204_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21882_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01205_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01206_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01207_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01208_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01209_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01210_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01211_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01212_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01213_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01214_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01215_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01216_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01217_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21895_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01218_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01219_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01220_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21898_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01221_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01222_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01223_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01224_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01225_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01226_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01227_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01228_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01229_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01230_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01231_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21909_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01232_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01233_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21911_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01234_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01235_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01236_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(clknet_leaf_86_i_clk),
    .D(_01237_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21915_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01238_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01239_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01240_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01241_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01242_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01243_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01244_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01245_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01246_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01247_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01248_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21926_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01249_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01250_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01251_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01252_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21930_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01253_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21931_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01254_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01255_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01256_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01257_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01258_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01259_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01260_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(clknet_leaf_12_i_clk),
    .D(_01261_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01262_),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01263_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01264_),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01265_),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(clknet_leaf_17_i_clk),
    .D(_01266_),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_2 _21944_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01267_),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01268_),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21946_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01269_),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21947_ (.CLK(clknet_leaf_14_i_clk),
    .D(_01270_),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21948_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01271_),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21949_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01272_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21950_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01273_),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(clknet_leaf_16_i_clk),
    .D(_01274_),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(clknet_leaf_17_i_clk),
    .D(_01275_),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(clknet_leaf_17_i_clk),
    .D(_01276_),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(clknet_leaf_20_i_clk),
    .D(_01277_),
    .Q(\rbzero.spi_registers.got_new_texadd3 ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(net217),
    .D(_01278_),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(net218),
    .D(_01279_),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(net219),
    .D(_01280_),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21958_ (.CLK(net220),
    .D(_01281_),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(net221),
    .D(_01282_),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21960_ (.CLK(net222),
    .D(_01283_),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(net223),
    .D(_01284_),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(net224),
    .D(_01285_),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21963_ (.CLK(net225),
    .D(_01286_),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(net226),
    .D(_01287_),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(net227),
    .D(_01288_),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(net228),
    .D(_01289_),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21967_ (.CLK(net229),
    .D(_01290_),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(net230),
    .D(_01291_),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(net231),
    .D(_01292_),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(net232),
    .D(_01293_),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21971_ (.CLK(net233),
    .D(_01294_),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(net234),
    .D(_01295_),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(net235),
    .D(_01296_),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(net236),
    .D(_01297_),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(net237),
    .D(_01298_),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(net238),
    .D(_01299_),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(net239),
    .D(_01300_),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(net240),
    .D(_01301_),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(net241),
    .D(_01302_),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(net242),
    .D(_01303_),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(net243),
    .D(_01304_),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(net244),
    .D(_01305_),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(net245),
    .D(_01306_),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(net246),
    .D(_01307_),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(net247),
    .D(_01308_),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(net248),
    .D(_01309_),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(net249),
    .D(_01310_),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(net250),
    .D(_01311_),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(net251),
    .D(_01312_),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(net252),
    .D(_01313_),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21991_ (.CLK(net253),
    .D(_01314_),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21992_ (.CLK(net254),
    .D(_01315_),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(net255),
    .D(_01316_),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(net256),
    .D(_01317_),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(net257),
    .D(_01318_),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(net258),
    .D(_01319_),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(net259),
    .D(_01320_),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21998_ (.CLK(net260),
    .D(_01321_),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(net261),
    .D(_01322_),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(net262),
    .D(_01323_),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(net263),
    .D(_01324_),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(net264),
    .D(_01325_),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(net265),
    .D(_01326_),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(net266),
    .D(_01327_),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(net267),
    .D(_01328_),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(net268),
    .D(_01329_),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(net269),
    .D(_01330_),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(net270),
    .D(_01331_),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(net271),
    .D(_01332_),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(net272),
    .D(_01333_),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(net273),
    .D(_01334_),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22012_ (.CLK(net274),
    .D(_01335_),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22013_ (.CLK(net275),
    .D(_01336_),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(net276),
    .D(_01337_),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(net277),
    .D(_01338_),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(net278),
    .D(_01339_),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(net279),
    .D(_01340_),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(net280),
    .D(_01341_),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(net281),
    .D(_01342_),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(net282),
    .D(_01343_),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(net283),
    .D(_01344_),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22022_ (.CLK(net284),
    .D(_01345_),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(net285),
    .D(_01346_),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(net286),
    .D(_01347_),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(net287),
    .D(_01348_),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(net288),
    .D(_01349_),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(net289),
    .D(_01350_),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(net290),
    .D(_01351_),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(net291),
    .D(_01352_),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(net292),
    .D(_01353_),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(net293),
    .D(_01354_),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(net294),
    .D(_01355_),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22033_ (.CLK(net295),
    .D(_01356_),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(net296),
    .D(_01357_),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(net297),
    .D(_01358_),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22036_ (.CLK(net298),
    .D(_01359_),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(net299),
    .D(_01360_),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(net300),
    .D(_01361_),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(net301),
    .D(_01362_),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(net302),
    .D(_01363_),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(net303),
    .D(_01364_),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(net304),
    .D(_01365_),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(net305),
    .D(_01366_),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(net306),
    .D(_01367_),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(net307),
    .D(_01368_),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22046_ (.CLK(net308),
    .D(_01369_),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22047_ (.CLK(net309),
    .D(_01370_),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22048_ (.CLK(net310),
    .D(_01371_),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22049_ (.CLK(net311),
    .D(_01372_),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22050_ (.CLK(net312),
    .D(_01373_),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22051_ (.CLK(net313),
    .D(_01374_),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22052_ (.CLK(net314),
    .D(_01375_),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22053_ (.CLK(net315),
    .D(_01376_),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22054_ (.CLK(net316),
    .D(_01377_),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22055_ (.CLK(net317),
    .D(_01378_),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22056_ (.CLK(net318),
    .D(_01379_),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22057_ (.CLK(net319),
    .D(_01380_),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22058_ (.CLK(net320),
    .D(_01381_),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22059_ (.CLK(net321),
    .D(_01382_),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22060_ (.CLK(net322),
    .D(_01383_),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22061_ (.CLK(net323),
    .D(_01384_),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22062_ (.CLK(net324),
    .D(_01385_),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22063_ (.CLK(net325),
    .D(_01386_),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22064_ (.CLK(net326),
    .D(_01387_),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22065_ (.CLK(net327),
    .D(_01388_),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22066_ (.CLK(net328),
    .D(_01389_),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22067_ (.CLK(net329),
    .D(_01390_),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22068_ (.CLK(net330),
    .D(_01391_),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22069_ (.CLK(net331),
    .D(_01392_),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22070_ (.CLK(net332),
    .D(_01393_),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22071_ (.CLK(net333),
    .D(_01394_),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22072_ (.CLK(net334),
    .D(_01395_),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22073_ (.CLK(net335),
    .D(_01396_),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22074_ (.CLK(net336),
    .D(_01397_),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22075_ (.CLK(net337),
    .D(_01398_),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22076_ (.CLK(net338),
    .D(_01399_),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22077_ (.CLK(net339),
    .D(_01400_),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22078_ (.CLK(net340),
    .D(_01401_),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22079_ (.CLK(net341),
    .D(_01402_),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22080_ (.CLK(net342),
    .D(_01403_),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22081_ (.CLK(net343),
    .D(_01404_),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22082_ (.CLK(net344),
    .D(_01405_),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22083_ (.CLK(net345),
    .D(_01406_),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22084_ (.CLK(net346),
    .D(_01407_),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22085_ (.CLK(net347),
    .D(_01408_),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22086_ (.CLK(net348),
    .D(_01409_),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22087_ (.CLK(net349),
    .D(_01410_),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22088_ (.CLK(net350),
    .D(_01411_),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22089_ (.CLK(net351),
    .D(_01412_),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22090_ (.CLK(net352),
    .D(_01413_),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22091_ (.CLK(net353),
    .D(_01414_),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22092_ (.CLK(net354),
    .D(_01415_),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22093_ (.CLK(net355),
    .D(_01416_),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22094_ (.CLK(net356),
    .D(_01417_),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22095_ (.CLK(net357),
    .D(_01418_),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22096_ (.CLK(net358),
    .D(_01419_),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22097_ (.CLK(net359),
    .D(_01420_),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22098_ (.CLK(net360),
    .D(_01421_),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22099_ (.CLK(net361),
    .D(_01422_),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22100_ (.CLK(net362),
    .D(_01423_),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22101_ (.CLK(net363),
    .D(_01424_),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22102_ (.CLK(net364),
    .D(_01425_),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22103_ (.CLK(net365),
    .D(_01426_),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22104_ (.CLK(net366),
    .D(_01427_),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22105_ (.CLK(net367),
    .D(_01428_),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22106_ (.CLK(net368),
    .D(_01429_),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22107_ (.CLK(net369),
    .D(_01430_),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22108_ (.CLK(net370),
    .D(_01431_),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22109_ (.CLK(net371),
    .D(_01432_),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22110_ (.CLK(net372),
    .D(_01433_),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22111_ (.CLK(net373),
    .D(_01434_),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22112_ (.CLK(net374),
    .D(_01435_),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22113_ (.CLK(net375),
    .D(_01436_),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22114_ (.CLK(net376),
    .D(_01437_),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22115_ (.CLK(net377),
    .D(_01438_),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22116_ (.CLK(net378),
    .D(_01439_),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22117_ (.CLK(net379),
    .D(_01440_),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22118_ (.CLK(net380),
    .D(_01441_),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22119_ (.CLK(net381),
    .D(_01442_),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22120_ (.CLK(net382),
    .D(_01443_),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22121_ (.CLK(net383),
    .D(_01444_),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22122_ (.CLK(net384),
    .D(_01445_),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22123_ (.CLK(net385),
    .D(_01446_),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22124_ (.CLK(net386),
    .D(_01447_),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22125_ (.CLK(net387),
    .D(_01448_),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22126_ (.CLK(net388),
    .D(_01449_),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22127_ (.CLK(net389),
    .D(_01450_),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22128_ (.CLK(net390),
    .D(_01451_),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22129_ (.CLK(net391),
    .D(_01452_),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22130_ (.CLK(net392),
    .D(_01453_),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22131_ (.CLK(net393),
    .D(_01454_),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22132_ (.CLK(net394),
    .D(_01455_),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22133_ (.CLK(net395),
    .D(_01456_),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22134_ (.CLK(net396),
    .D(_01457_),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22135_ (.CLK(net397),
    .D(_01458_),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22136_ (.CLK(net398),
    .D(_01459_),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22137_ (.CLK(net399),
    .D(_01460_),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22138_ (.CLK(net400),
    .D(_01461_),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22139_ (.CLK(net401),
    .D(_01462_),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22140_ (.CLK(net402),
    .D(_01463_),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22141_ (.CLK(net403),
    .D(_01464_),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22142_ (.CLK(net404),
    .D(_01465_),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22143_ (.CLK(net405),
    .D(_01466_),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22144_ (.CLK(net406),
    .D(_01467_),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22145_ (.CLK(net407),
    .D(_01468_),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22146_ (.CLK(net408),
    .D(_01469_),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22147_ (.CLK(net409),
    .D(_01470_),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22148_ (.CLK(net410),
    .D(_01471_),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22149_ (.CLK(net411),
    .D(_01472_),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22150_ (.CLK(net412),
    .D(_01473_),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22151_ (.CLK(net413),
    .D(_01474_),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22152_ (.CLK(net414),
    .D(_01475_),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22153_ (.CLK(net415),
    .D(_01476_),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22154_ (.CLK(net416),
    .D(_01477_),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22155_ (.CLK(net417),
    .D(_01478_),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22156_ (.CLK(net418),
    .D(_01479_),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22157_ (.CLK(net419),
    .D(_01480_),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22158_ (.CLK(net420),
    .D(_01481_),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22159_ (.CLK(net421),
    .D(_01482_),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22160_ (.CLK(net422),
    .D(_01483_),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22161_ (.CLK(net423),
    .D(_01484_),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22162_ (.CLK(net424),
    .D(_01485_),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22163_ (.CLK(net425),
    .D(_01486_),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22164_ (.CLK(net426),
    .D(_01487_),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22165_ (.CLK(net427),
    .D(_01488_),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22166_ (.CLK(net428),
    .D(_01489_),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22167_ (.CLK(net429),
    .D(_01490_),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22168_ (.CLK(net430),
    .D(_01491_),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22169_ (.CLK(net431),
    .D(_01492_),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22170_ (.CLK(net432),
    .D(_01493_),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22171_ (.CLK(net433),
    .D(_01494_),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22172_ (.CLK(net434),
    .D(_01495_),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22173_ (.CLK(net435),
    .D(_01496_),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22174_ (.CLK(net436),
    .D(_01497_),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22175_ (.CLK(net437),
    .D(_01498_),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22176_ (.CLK(net438),
    .D(_01499_),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22177_ (.CLK(net439),
    .D(_01500_),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22178_ (.CLK(net440),
    .D(_01501_),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22179_ (.CLK(net441),
    .D(_01502_),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22180_ (.CLK(net442),
    .D(_01503_),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22181_ (.CLK(net443),
    .D(_01504_),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22182_ (.CLK(net444),
    .D(_01505_),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22183_ (.CLK(net445),
    .D(_01506_),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22184_ (.CLK(net446),
    .D(_01507_),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22185_ (.CLK(net447),
    .D(_01508_),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22186_ (.CLK(net448),
    .D(_01509_),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22187_ (.CLK(net449),
    .D(_01510_),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22188_ (.CLK(net450),
    .D(_01511_),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22189_ (.CLK(net451),
    .D(_01512_),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22190_ (.CLK(net452),
    .D(_01513_),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22191_ (.CLK(net453),
    .D(_01514_),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22192_ (.CLK(net454),
    .D(_01515_),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22193_ (.CLK(net455),
    .D(_01516_),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22194_ (.CLK(net456),
    .D(_01517_),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22195_ (.CLK(net457),
    .D(_01518_),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22196_ (.CLK(net458),
    .D(_01519_),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22197_ (.CLK(net459),
    .D(_01520_),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22198_ (.CLK(net460),
    .D(_01521_),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22199_ (.CLK(net461),
    .D(_01522_),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22200_ (.CLK(net462),
    .D(_01523_),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22201_ (.CLK(net463),
    .D(_01524_),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22202_ (.CLK(net464),
    .D(_01525_),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22203_ (.CLK(net465),
    .D(_01526_),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22204_ (.CLK(net466),
    .D(_01527_),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22205_ (.CLK(net467),
    .D(_01528_),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22206_ (.CLK(net468),
    .D(_01529_),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22207_ (.CLK(net469),
    .D(_01530_),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22208_ (.CLK(net470),
    .D(_01531_),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22209_ (.CLK(net471),
    .D(_01532_),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22210_ (.CLK(net472),
    .D(_01533_),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22211_ (.CLK(net473),
    .D(_01534_),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22212_ (.CLK(net474),
    .D(_01535_),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22213_ (.CLK(net475),
    .D(_01536_),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22214_ (.CLK(net476),
    .D(_01537_),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22215_ (.CLK(net477),
    .D(_01538_),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22216_ (.CLK(net478),
    .D(_01539_),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22217_ (.CLK(net479),
    .D(_01540_),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22218_ (.CLK(net480),
    .D(_01541_),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22219_ (.CLK(net481),
    .D(_01542_),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22220_ (.CLK(net482),
    .D(_01543_),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22221_ (.CLK(net483),
    .D(_01544_),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22222_ (.CLK(net484),
    .D(_01545_),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22223_ (.CLK(net485),
    .D(_01546_),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22224_ (.CLK(net486),
    .D(_01547_),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22225_ (.CLK(net487),
    .D(_01548_),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22226_ (.CLK(net488),
    .D(_01549_),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22227_ (.CLK(net489),
    .D(_01550_),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22228_ (.CLK(net490),
    .D(_01551_),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22229_ (.CLK(net491),
    .D(_01552_),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22230_ (.CLK(net492),
    .D(_01553_),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22231_ (.CLK(net493),
    .D(_01554_),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22232_ (.CLK(net494),
    .D(_01555_),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22233_ (.CLK(net495),
    .D(_01556_),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22234_ (.CLK(net496),
    .D(_01557_),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22235_ (.CLK(net497),
    .D(_01558_),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22236_ (.CLK(net498),
    .D(_01559_),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22237_ (.CLK(net499),
    .D(_01560_),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22238_ (.CLK(net500),
    .D(_01561_),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22239_ (.CLK(net501),
    .D(_01562_),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22240_ (.CLK(net502),
    .D(_01563_),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22241_ (.CLK(net503),
    .D(_01564_),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22242_ (.CLK(net504),
    .D(_01565_),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22243_ (.CLK(net505),
    .D(_01566_),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22244_ (.CLK(net506),
    .D(_01567_),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22245_ (.CLK(net507),
    .D(_01568_),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22246_ (.CLK(net508),
    .D(_01569_),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22247_ (.CLK(net509),
    .D(_01570_),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22248_ (.CLK(net510),
    .D(_01571_),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22249_ (.CLK(net511),
    .D(_01572_),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22250_ (.CLK(net512),
    .D(_01573_),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22251_ (.CLK(net133),
    .D(_01574_),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22252_ (.CLK(net134),
    .D(_01575_),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22253_ (.CLK(net135),
    .D(_01576_),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22254_ (.CLK(net136),
    .D(_01577_),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22255_ (.CLK(net137),
    .D(_01578_),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22256_ (.CLK(net138),
    .D(_01579_),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22257_ (.CLK(net139),
    .D(_01580_),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22258_ (.CLK(net140),
    .D(_01581_),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22259_ (.CLK(net141),
    .D(_01582_),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22260_ (.CLK(net142),
    .D(_01583_),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22261_ (.CLK(net143),
    .D(_01584_),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22262_ (.CLK(net144),
    .D(_01585_),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22263_ (.CLK(net145),
    .D(_01586_),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22264_ (.CLK(net146),
    .D(_01587_),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22265_ (.CLK(net147),
    .D(_01588_),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22266_ (.CLK(net148),
    .D(_01589_),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22267_ (.CLK(net149),
    .D(_01590_),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22268_ (.CLK(net150),
    .D(_01591_),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22269_ (.CLK(net151),
    .D(_01592_),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22270_ (.CLK(net152),
    .D(_01593_),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22271_ (.CLK(net129),
    .D(_01594_),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22272_ (.CLK(net130),
    .D(_01595_),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22273_ (.CLK(net131),
    .D(_01596_),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22274_ (.CLK(net132),
    .D(_01597_),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22275_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01598_),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22276_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01599_),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22277_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01600_),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _22278_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01601_),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _22279_ (.CLK(clknet_leaf_65_i_clk),
    .D(_01602_),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22280_ (.CLK(clknet_leaf_65_i_clk),
    .D(_01603_),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22281_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01604_),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22282_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01605_),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22283_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01606_),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _22284_ (.CLK(clknet_leaf_66_i_clk),
    .D(_01607_),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _22285_ (.CLK(clknet_leaf_65_i_clk),
    .D(_01608_),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _22286_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01609_),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _22287_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01610_),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _22288_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01611_),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22289_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01612_),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22290_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01613_),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_2 _22291_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01614_),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22292_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01615_),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22293_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01616_),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22294_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01617_),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22295_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01618_),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22296_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01619_),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22297_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01620_),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22298_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01621_),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_4 _22299_ (.CLK(clknet_leaf_64_i_clk),
    .D(_01622_),
    .Q(\rbzero.trace_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22300_ (.CLK(clknet_leaf_64_i_clk),
    .D(_01623_),
    .Q(\rbzero.trace_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22301_ (.CLK(clknet_leaf_64_i_clk),
    .D(_01624_),
    .Q(\rbzero.trace_state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _22302_ (.CLK(clknet_leaf_48_i_clk),
    .D(_01625_),
    .Q(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22303_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01626_),
    .Q(\reg_gpout[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22304_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01627_),
    .Q(\reg_gpout[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22305_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01628_),
    .Q(\reg_gpout[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22306_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01629_),
    .Q(\reg_gpout[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22307_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01630_),
    .Q(\reg_gpout[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22308_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01631_),
    .Q(\reg_gpout[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22309_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01632_),
    .Q(reg_hsync));
 sky130_fd_sc_hd__dfxtp_1 _22310_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01633_),
    .Q(reg_vsync));
 sky130_fd_sc_hd__dfxtp_1 _22311_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01634_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22312_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01635_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22313_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01636_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22314_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01637_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22315_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01638_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22316_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01639_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22317_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01640_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22318_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01641_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22319_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01642_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22320_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01643_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22321_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01644_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22322_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01645_),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22323_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01646_),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22324_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01647_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22325_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01648_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22326_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01649_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22327_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01650_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22328_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01651_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22329_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01652_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22330_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01653_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22331_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01654_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22332_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01655_),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22333_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01656_),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22334_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01657_),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22335_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01658_),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22336_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01659_),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22337_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01660_),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22338_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01661_),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22339_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01662_),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.HI(net111));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_122 (.HI(net122));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_124 (.HI(net124));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_125 (.HI(net125));
 sky130_fd_sc_hd__inv_2 _11576__1 (.A(clknet_1_1__leaf__04767_),
    .Y(net126));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.HI(net110));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(i_debug_map_overlay),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(i_debug_trace_overlay),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(i_debug_vec_overlay),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(i_gpout0_sel[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(i_gpout0_sel[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(i_gpout0_sel[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(i_gpout0_sel[3]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(i_gpout0_sel[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(i_gpout0_sel[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(i_gpout1_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(i_gpout1_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(i_gpout1_sel[2]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(i_gpout1_sel[3]),
    .X(net13));
 sky130_fd_sc_hd__buf_6 input14 (.A(i_gpout1_sel[4]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(i_gpout1_sel[5]),
    .X(net15));
 sky130_fd_sc_hd__buf_6 input16 (.A(i_gpout2_sel[0]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(i_gpout2_sel[1]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(i_gpout2_sel[2]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(i_gpout2_sel[3]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(i_gpout2_sel[4]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(i_gpout2_sel[5]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(i_gpout3_sel[0]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(i_gpout3_sel[1]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(i_gpout3_sel[2]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(i_gpout3_sel[3]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(i_gpout3_sel[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(i_gpout3_sel[5]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(i_gpout4_sel[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(i_gpout4_sel[1]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(i_gpout4_sel[2]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(i_gpout4_sel[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(i_gpout4_sel[4]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(i_gpout4_sel[5]),
    .X(net33));
 sky130_fd_sc_hd__buf_6 input34 (.A(i_gpout5_sel[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_8 input35 (.A(i_gpout5_sel[1]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(i_gpout5_sel[2]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(i_gpout5_sel[3]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(i_gpout5_sel[4]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(i_gpout5_sel[5]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_16 input40 (.A(i_mode[0]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_16 input41 (.A(i_mode[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_8 input42 (.A(i_mode[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(i_reg_csb),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(i_reg_mosi),
    .X(net44));
 sky130_fd_sc_hd__buf_6 input45 (.A(i_reg_outs_enb),
    .X(net45));
 sky130_fd_sc_hd__buf_8 input46 (.A(i_reg_sclk),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(i_reset_lock_a),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_reset_lock_b),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(i_test_wb_clk_i),
    .X(net49));
 sky130_fd_sc_hd__buf_6 input50 (.A(i_tex_in[0]),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input51 (.A(i_tex_in[1]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(i_tex_in[2]),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input53 (.A(i_tex_in[3]),
    .X(net53));
 sky130_fd_sc_hd__buf_8 input54 (.A(i_vec_csb),
    .X(net54));
 sky130_fd_sc_hd__buf_4 input55 (.A(i_vec_mosi),
    .X(net55));
 sky130_fd_sc_hd__buf_8 input56 (.A(i_vec_sclk),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(o_hsync));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(o_reset));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(o_tex_csb));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(o_tex_out0));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net126),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(o_vsync));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_76 (.LO(net76));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_1_0__leaf__04767_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 net99_3 (.A(clknet_1_0__leaf__04767_),
    .Y(net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_opt_2_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_opt_3_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_opt_4_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_opt_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_opt_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05795_ (.A(_05795_),
    .X(clknet_0__05795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05795_ (.A(clknet_0__05795_),
    .X(clknet_1_0__leaf__05795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05795_ (.A(clknet_0__05795_),
    .X(clknet_1_1__leaf__05795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04767_ (.A(_04767_),
    .X(clknet_0__04767_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04767_ (.A(clknet_0__04767_),
    .X(clknet_1_0__leaf__04767_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04767_ (.A(clknet_0__04767_),
    .X(clknet_1_1__leaf__04767_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05854_ (.A(_05854_),
    .X(clknet_0__05854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05854_ (.A(clknet_0__05854_),
    .X(clknet_1_0__leaf__05854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05854_ (.A(clknet_0__05854_),
    .X(clknet_1_1__leaf__05854_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__06092_ (.A(_06092_),
    .X(clknet_0__06092_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__06092_ (.A(clknet_0__06092_),
    .X(clknet_1_0__leaf__06092_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__06092_ (.A(clknet_0__06092_),
    .X(clknet_1_1__leaf__06092_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03944_ (.A(_03944_),
    .X(clknet_0__03944_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03944_ (.A(clknet_0__03944_),
    .X(clknet_1_0__leaf__03944_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03944_ (.A(clknet_0__03944_),
    .X(clknet_1_1__leaf__03944_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03943_ (.A(_03943_),
    .X(clknet_0__03943_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03943_ (.A(clknet_0__03943_),
    .X(clknet_1_0__leaf__03943_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03943_ (.A(clknet_0__03943_),
    .X(clknet_1_1__leaf__03943_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03932_ (.A(_03932_),
    .X(clknet_0__03932_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03932_ (.A(clknet_0__03932_),
    .X(clknet_1_0__leaf__03932_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03932_ (.A(clknet_0__03932_),
    .X(clknet_1_1__leaf__03932_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03942_ (.A(_03942_),
    .X(clknet_0__03942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03942_ (.A(clknet_0__03942_),
    .X(clknet_1_0__leaf__03942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03942_ (.A(clknet_0__03942_),
    .X(clknet_1_1__leaf__03942_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03941_ (.A(_03941_),
    .X(clknet_0__03941_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03941_ (.A(clknet_0__03941_),
    .X(clknet_1_0__leaf__03941_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03941_ (.A(clknet_0__03941_),
    .X(clknet_1_1__leaf__03941_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03940_ (.A(_03940_),
    .X(clknet_0__03940_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03940_ (.A(clknet_0__03940_),
    .X(clknet_1_0__leaf__03940_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03940_ (.A(clknet_0__03940_),
    .X(clknet_1_1__leaf__03940_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03939_ (.A(_03939_),
    .X(clknet_0__03939_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03939_ (.A(clknet_0__03939_),
    .X(clknet_1_0__leaf__03939_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03939_ (.A(clknet_0__03939_),
    .X(clknet_1_1__leaf__03939_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03938_ (.A(_03938_),
    .X(clknet_0__03938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03938_ (.A(clknet_0__03938_),
    .X(clknet_1_0__leaf__03938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03938_ (.A(clknet_0__03938_),
    .X(clknet_1_1__leaf__03938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03937_ (.A(_03937_),
    .X(clknet_0__03937_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03937_ (.A(clknet_0__03937_),
    .X(clknet_1_0__leaf__03937_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03937_ (.A(clknet_0__03937_),
    .X(clknet_1_1__leaf__03937_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03936_ (.A(_03936_),
    .X(clknet_0__03936_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03936_ (.A(clknet_0__03936_),
    .X(clknet_1_0__leaf__03936_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03936_ (.A(clknet_0__03936_),
    .X(clknet_1_1__leaf__03936_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03935_ (.A(_03935_),
    .X(clknet_0__03935_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03935_ (.A(clknet_0__03935_),
    .X(clknet_1_0__leaf__03935_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03935_ (.A(clknet_0__03935_),
    .X(clknet_1_1__leaf__03935_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03934_ (.A(_03934_),
    .X(clknet_0__03934_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03934_ (.A(clknet_0__03934_),
    .X(clknet_1_0__leaf__03934_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03934_ (.A(clknet_0__03934_),
    .X(clknet_1_1__leaf__03934_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03933_ (.A(_03933_),
    .X(clknet_0__03933_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03933_ (.A(clknet_0__03933_),
    .X(clknet_1_0__leaf__03933_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03933_ (.A(clknet_0__03933_),
    .X(clknet_1_1__leaf__03933_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03921_ (.A(_03921_),
    .X(clknet_0__03921_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03921_ (.A(clknet_0__03921_),
    .X(clknet_1_0__leaf__03921_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03921_ (.A(clknet_0__03921_),
    .X(clknet_1_1__leaf__03921_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03931_ (.A(_03931_),
    .X(clknet_0__03931_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03931_ (.A(clknet_0__03931_),
    .X(clknet_1_0__leaf__03931_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03931_ (.A(clknet_0__03931_),
    .X(clknet_1_1__leaf__03931_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03930_ (.A(_03930_),
    .X(clknet_0__03930_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03930_ (.A(clknet_0__03930_),
    .X(clknet_1_0__leaf__03930_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03930_ (.A(clknet_0__03930_),
    .X(clknet_1_1__leaf__03930_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03929_ (.A(_03929_),
    .X(clknet_0__03929_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03929_ (.A(clknet_0__03929_),
    .X(clknet_1_0__leaf__03929_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03929_ (.A(clknet_0__03929_),
    .X(clknet_1_1__leaf__03929_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03928_ (.A(_03928_),
    .X(clknet_0__03928_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03928_ (.A(clknet_0__03928_),
    .X(clknet_1_0__leaf__03928_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03928_ (.A(clknet_0__03928_),
    .X(clknet_1_1__leaf__03928_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03927_ (.A(_03927_),
    .X(clknet_0__03927_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03927_ (.A(clknet_0__03927_),
    .X(clknet_1_0__leaf__03927_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03927_ (.A(clknet_0__03927_),
    .X(clknet_1_1__leaf__03927_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03926_ (.A(_03926_),
    .X(clknet_0__03926_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03926_ (.A(clknet_0__03926_),
    .X(clknet_1_0__leaf__03926_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03926_ (.A(clknet_0__03926_),
    .X(clknet_1_1__leaf__03926_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03925_ (.A(_03925_),
    .X(clknet_0__03925_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03925_ (.A(clknet_0__03925_),
    .X(clknet_1_0__leaf__03925_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03925_ (.A(clknet_0__03925_),
    .X(clknet_1_1__leaf__03925_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03924_ (.A(_03924_),
    .X(clknet_0__03924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03924_ (.A(clknet_0__03924_),
    .X(clknet_1_0__leaf__03924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03924_ (.A(clknet_0__03924_),
    .X(clknet_1_1__leaf__03924_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03923_ (.A(_03923_),
    .X(clknet_0__03923_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03923_ (.A(clknet_0__03923_),
    .X(clknet_1_0__leaf__03923_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03923_ (.A(clknet_0__03923_),
    .X(clknet_1_1__leaf__03923_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03922_ (.A(_03922_),
    .X(clknet_0__03922_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03922_ (.A(clknet_0__03922_),
    .X(clknet_1_0__leaf__03922_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03922_ (.A(clknet_0__03922_),
    .X(clknet_1_1__leaf__03922_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03711_ (.A(_03711_),
    .X(clknet_0__03711_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03711_ (.A(clknet_0__03711_),
    .X(clknet_1_0__leaf__03711_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03711_ (.A(clknet_0__03711_),
    .X(clknet_1_1__leaf__03711_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03920_ (.A(_03920_),
    .X(clknet_0__03920_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03920_ (.A(clknet_0__03920_),
    .X(clknet_1_0__leaf__03920_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03920_ (.A(clknet_0__03920_),
    .X(clknet_1_1__leaf__03920_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03919_ (.A(_03919_),
    .X(clknet_0__03919_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03919_ (.A(clknet_0__03919_),
    .X(clknet_1_0__leaf__03919_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03919_ (.A(clknet_0__03919_),
    .X(clknet_1_1__leaf__03919_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03918_ (.A(_03918_),
    .X(clknet_0__03918_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03918_ (.A(clknet_0__03918_),
    .X(clknet_1_0__leaf__03918_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03918_ (.A(clknet_0__03918_),
    .X(clknet_1_1__leaf__03918_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03917_ (.A(_03917_),
    .X(clknet_0__03917_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03917_ (.A(clknet_0__03917_),
    .X(clknet_1_0__leaf__03917_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03917_ (.A(clknet_0__03917_),
    .X(clknet_1_1__leaf__03917_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03916_ (.A(_03916_),
    .X(clknet_0__03916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03916_ (.A(clknet_0__03916_),
    .X(clknet_1_0__leaf__03916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03916_ (.A(clknet_0__03916_),
    .X(clknet_1_1__leaf__03916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03915_ (.A(_03915_),
    .X(clknet_0__03915_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03915_ (.A(clknet_0__03915_),
    .X(clknet_1_0__leaf__03915_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03915_ (.A(clknet_0__03915_),
    .X(clknet_1_1__leaf__03915_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03914_ (.A(_03914_),
    .X(clknet_0__03914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03914_ (.A(clknet_0__03914_),
    .X(clknet_1_0__leaf__03914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03914_ (.A(clknet_0__03914_),
    .X(clknet_1_1__leaf__03914_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03913_ (.A(_03913_),
    .X(clknet_0__03913_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03913_ (.A(clknet_0__03913_),
    .X(clknet_1_0__leaf__03913_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03913_ (.A(clknet_0__03913_),
    .X(clknet_1_1__leaf__03913_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03912_ (.A(_03912_),
    .X(clknet_0__03912_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03912_ (.A(clknet_0__03912_),
    .X(clknet_1_0__leaf__03912_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03912_ (.A(clknet_0__03912_),
    .X(clknet_1_1__leaf__03912_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03712_ (.A(_03712_),
    .X(clknet_0__03712_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03712_ (.A(clknet_0__03712_),
    .X(clknet_1_0__leaf__03712_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03712_ (.A(clknet_0__03712_),
    .X(clknet_1_1__leaf__03712_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03704_ (.A(_03704_),
    .X(clknet_0__03704_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03704_ (.A(clknet_0__03704_),
    .X(clknet_1_0__leaf__03704_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03704_ (.A(clknet_0__03704_),
    .X(clknet_1_1__leaf__03704_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03710_ (.A(_03710_),
    .X(clknet_0__03710_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03710_ (.A(clknet_0__03710_),
    .X(clknet_1_0__leaf__03710_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03710_ (.A(clknet_0__03710_),
    .X(clknet_1_1__leaf__03710_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03709_ (.A(_03709_),
    .X(clknet_0__03709_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03709_ (.A(clknet_0__03709_),
    .X(clknet_1_0__leaf__03709_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03709_ (.A(clknet_0__03709_),
    .X(clknet_1_1__leaf__03709_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03708_ (.A(_03708_),
    .X(clknet_0__03708_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03708_ (.A(clknet_0__03708_),
    .X(clknet_1_0__leaf__03708_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03708_ (.A(clknet_0__03708_),
    .X(clknet_1_1__leaf__03708_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03707_ (.A(_03707_),
    .X(clknet_0__03707_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03707_ (.A(clknet_0__03707_),
    .X(clknet_1_0__leaf__03707_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03707_ (.A(clknet_0__03707_),
    .X(clknet_1_1__leaf__03707_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03706_ (.A(_03706_),
    .X(clknet_0__03706_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03706_ (.A(clknet_0__03706_),
    .X(clknet_1_0__leaf__03706_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03706_ (.A(clknet_0__03706_),
    .X(clknet_1_1__leaf__03706_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03705_ (.A(_03705_),
    .X(clknet_0__03705_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03705_ (.A(clknet_0__03705_),
    .X(clknet_1_0__leaf__03705_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03705_ (.A(clknet_0__03705_),
    .X(clknet_1_1__leaf__03705_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__06036_ (.A(_06036_),
    .X(clknet_0__06036_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__06036_ (.A(clknet_0__06036_),
    .X(clknet_1_0__leaf__06036_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__06036_ (.A(clknet_0__06036_),
    .X(clknet_1_1__leaf__06036_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05977_ (.A(_05977_),
    .X(clknet_0__05977_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05977_ (.A(clknet_0__05977_),
    .X(clknet_1_0__leaf__05977_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05977_ (.A(clknet_0__05977_),
    .X(clknet_1_1__leaf__05977_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05916_ (.A(_05916_),
    .X(clknet_0__05916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05916_ (.A(clknet_0__05916_),
    .X(clknet_1_0__leaf__05916_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05916_ (.A(clknet_0__05916_),
    .X(clknet_1_1__leaf__05916_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rbzero.tex_r1[40] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\rbzero.spi_registers.new_other[10] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\rbzero.spi_registers.new_vinf ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\rbzero.spi_registers.new_other[7] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\rbzero.spi_registers.new_other[8] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\rbzero.spi_registers.new_other[1] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\rbzero.spi_registers.new_other[2] ),
    .X(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_04955_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_05053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_05351_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_08207_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_08249_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_08355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_08355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_08355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_08556_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_09883_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_09887_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_09889_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_09946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_09946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\rbzero.texV[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\rbzero.texu_hot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_04563_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_04970_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_05053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_05727_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_08481_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_09938_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_10030_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net53));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1226 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1226 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_982 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1252 ();
 assign o_rgb[0] = net76;
 assign o_rgb[10] = net84;
 assign o_rgb[11] = net85;
 assign o_rgb[12] = net86;
 assign o_rgb[13] = net87;
 assign o_rgb[16] = net88;
 assign o_rgb[17] = net89;
 assign o_rgb[18] = net90;
 assign o_rgb[19] = net91;
 assign o_rgb[1] = net77;
 assign o_rgb[20] = net92;
 assign o_rgb[21] = net93;
 assign o_rgb[2] = net78;
 assign o_rgb[3] = net79;
 assign o_rgb[4] = net80;
 assign o_rgb[5] = net81;
 assign o_rgb[8] = net82;
 assign o_rgb[9] = net83;
 assign ones[0] = net110;
 assign ones[10] = net120;
 assign ones[11] = net121;
 assign ones[12] = net122;
 assign ones[13] = net123;
 assign ones[14] = net124;
 assign ones[15] = net125;
 assign ones[1] = net111;
 assign ones[2] = net112;
 assign ones[3] = net113;
 assign ones[4] = net114;
 assign ones[5] = net115;
 assign ones[6] = net116;
 assign ones[7] = net117;
 assign ones[8] = net118;
 assign ones[9] = net119;
 assign zeros[0] = net94;
 assign zeros[10] = net104;
 assign zeros[11] = net105;
 assign zeros[12] = net106;
 assign zeros[13] = net107;
 assign zeros[14] = net108;
 assign zeros[15] = net109;
 assign zeros[1] = net95;
 assign zeros[2] = net96;
 assign zeros[3] = net97;
 assign zeros[4] = net98;
 assign zeros[5] = net99;
 assign zeros[6] = net100;
 assign zeros[7] = net101;
 assign zeros[8] = net102;
 assign zeros[9] = net103;
endmodule

