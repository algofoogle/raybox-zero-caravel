magic
tech sky130A
magscale 1 2
timestamp 1699236789
<< nwell >>
rect 1066 117765 116970 118086
rect 1066 116677 116970 117243
rect 1066 115589 116970 116155
rect 1066 114501 116970 115067
rect 1066 113413 116970 113979
rect 1066 112325 116970 112891
rect 1066 111237 116970 111803
rect 1066 110149 116970 110715
rect 1066 109061 116970 109627
rect 1066 107973 116970 108539
rect 1066 106885 116970 107451
rect 1066 105797 116970 106363
rect 1066 104709 116970 105275
rect 1066 103621 116970 104187
rect 1066 102533 116970 103099
rect 1066 101445 116970 102011
rect 1066 100357 116970 100923
rect 1066 99269 116970 99835
rect 1066 98181 116970 98747
rect 1066 97093 116970 97659
rect 1066 96005 116970 96571
rect 1066 94917 116970 95483
rect 1066 93829 116970 94395
rect 1066 92741 116970 93307
rect 1066 91653 116970 92219
rect 1066 90565 116970 91131
rect 1066 89477 116970 90043
rect 1066 88389 116970 88955
rect 1066 87301 116970 87867
rect 1066 86213 116970 86779
rect 1066 85125 116970 85691
rect 1066 84037 116970 84603
rect 1066 82949 116970 83515
rect 1066 81861 116970 82427
rect 1066 80773 116970 81339
rect 1066 79685 116970 80251
rect 1066 78597 116970 79163
rect 1066 77509 116970 78075
rect 1066 76421 116970 76987
rect 1066 75333 116970 75899
rect 1066 74245 116970 74811
rect 1066 73157 116970 73723
rect 1066 72069 116970 72635
rect 1066 70981 116970 71547
rect 1066 69893 116970 70459
rect 1066 68805 116970 69371
rect 1066 67717 116970 68283
rect 1066 66629 116970 67195
rect 1066 65541 116970 66107
rect 1066 64453 116970 65019
rect 1066 63365 116970 63931
rect 1066 62277 116970 62843
rect 1066 61189 116970 61755
rect 1066 60101 116970 60667
rect 1066 59013 116970 59579
rect 1066 57925 116970 58491
rect 1066 56837 116970 57403
rect 1066 55749 116970 56315
rect 1066 54661 116970 55227
rect 1066 53573 116970 54139
rect 1066 52485 116970 53051
rect 1066 51397 116970 51963
rect 1066 50309 116970 50875
rect 1066 49221 116970 49787
rect 1066 48133 116970 48699
rect 1066 47045 116970 47611
rect 1066 45957 116970 46523
rect 1066 44869 116970 45435
rect 1066 43781 116970 44347
rect 1066 42693 116970 43259
rect 1066 41605 116970 42171
rect 1066 40517 116970 41083
rect 1066 39429 116970 39995
rect 1066 38341 116970 38907
rect 1066 37253 116970 37819
rect 1066 36165 116970 36731
rect 1066 35077 116970 35643
rect 1066 33989 116970 34555
rect 1066 32901 116970 33467
rect 1066 31813 116970 32379
rect 1066 30725 116970 31291
rect 1066 29637 116970 30203
rect 1066 28549 116970 29115
rect 1066 27461 116970 28027
rect 1066 26373 116970 26939
rect 1066 25285 116970 25851
rect 1066 24197 116970 24763
rect 1066 23109 116970 23675
rect 1066 22021 116970 22587
rect 1066 20933 116970 21499
rect 1066 19845 116970 20411
rect 1066 18757 116970 19323
rect 1066 17669 116970 18235
rect 1066 16581 116970 17147
rect 1066 15493 116970 16059
rect 1066 14405 116970 14971
rect 1066 13317 116970 13883
rect 1066 12229 116970 12795
rect 1066 11141 116970 11707
rect 1066 10053 116970 10619
rect 1066 8965 116970 9531
rect 1066 7877 116970 8443
rect 1066 6789 116970 7355
rect 1066 5701 116970 6267
rect 1066 4613 116970 5179
rect 1066 3525 116970 4091
rect 1066 2437 116970 3003
<< obsli1 >>
rect 1104 2159 116932 118065
<< obsm1 >>
rect 1104 2128 117194 119400
<< metal2 >>
rect 2686 119451 2742 120251
rect 4986 119451 5042 120251
rect 7286 119451 7342 120251
rect 9586 119451 9642 120251
rect 11886 119451 11942 120251
rect 14186 119451 14242 120251
rect 16486 119451 16542 120251
rect 18786 119451 18842 120251
rect 21086 119451 21142 120251
rect 23386 119451 23442 120251
rect 25686 119451 25742 120251
rect 27986 119451 28042 120251
rect 30286 119451 30342 120251
rect 32586 119451 32642 120251
rect 34886 119451 34942 120251
rect 37186 119451 37242 120251
rect 39486 119451 39542 120251
rect 41786 119451 41842 120251
rect 44086 119451 44142 120251
rect 46386 119451 46442 120251
rect 48686 119451 48742 120251
rect 50986 119451 51042 120251
rect 53286 119451 53342 120251
rect 55586 119451 55642 120251
rect 57886 119451 57942 120251
rect 60186 119451 60242 120251
rect 62486 119451 62542 120251
rect 64786 119451 64842 120251
rect 67086 119451 67142 120251
rect 69386 119451 69442 120251
rect 71686 119451 71742 120251
rect 73986 119451 74042 120251
rect 76286 119451 76342 120251
rect 78586 119451 78642 120251
rect 80886 119451 80942 120251
rect 83186 119451 83242 120251
rect 85486 119451 85542 120251
rect 87786 119451 87842 120251
rect 90086 119451 90142 120251
rect 92386 119451 92442 120251
rect 94686 119451 94742 120251
rect 96986 119451 97042 120251
rect 99286 119451 99342 120251
rect 101586 119451 101642 120251
rect 103886 119451 103942 120251
rect 106186 119451 106242 120251
rect 108486 119451 108542 120251
rect 110786 119451 110842 120251
rect 113086 119451 113142 120251
rect 115386 119451 115442 120251
rect 3054 0 3110 800
rect 5998 0 6054 800
rect 8942 0 8998 800
rect 11886 0 11942 800
rect 14830 0 14886 800
rect 17774 0 17830 800
rect 20718 0 20774 800
rect 23662 0 23718 800
rect 26606 0 26662 800
rect 29550 0 29606 800
rect 32494 0 32550 800
rect 35438 0 35494 800
rect 38382 0 38438 800
rect 41326 0 41382 800
rect 44270 0 44326 800
rect 47214 0 47270 800
rect 50158 0 50214 800
rect 53102 0 53158 800
rect 56046 0 56102 800
rect 58990 0 59046 800
rect 61934 0 61990 800
rect 64878 0 64934 800
rect 67822 0 67878 800
rect 70766 0 70822 800
rect 73710 0 73766 800
rect 76654 0 76710 800
rect 79598 0 79654 800
rect 82542 0 82598 800
rect 85486 0 85542 800
rect 88430 0 88486 800
rect 91374 0 91430 800
rect 94318 0 94374 800
rect 97262 0 97318 800
rect 100206 0 100262 800
rect 103150 0 103206 800
rect 106094 0 106150 800
rect 109038 0 109094 800
rect 111982 0 112038 800
rect 114926 0 114982 800
<< obsm2 >>
rect 3056 119395 4930 119490
rect 5098 119395 7230 119490
rect 7398 119395 9530 119490
rect 9698 119395 11830 119490
rect 11998 119395 14130 119490
rect 14298 119395 16430 119490
rect 16598 119395 18730 119490
rect 18898 119395 21030 119490
rect 21198 119395 23330 119490
rect 23498 119395 25630 119490
rect 25798 119395 27930 119490
rect 28098 119395 30230 119490
rect 30398 119395 32530 119490
rect 32698 119395 34830 119490
rect 34998 119395 37130 119490
rect 37298 119395 39430 119490
rect 39598 119395 41730 119490
rect 41898 119395 44030 119490
rect 44198 119395 46330 119490
rect 46498 119395 48630 119490
rect 48798 119395 50930 119490
rect 51098 119395 53230 119490
rect 53398 119395 55530 119490
rect 55698 119395 57830 119490
rect 57998 119395 60130 119490
rect 60298 119395 62430 119490
rect 62598 119395 64730 119490
rect 64898 119395 67030 119490
rect 67198 119395 69330 119490
rect 69498 119395 71630 119490
rect 71798 119395 73930 119490
rect 74098 119395 76230 119490
rect 76398 119395 78530 119490
rect 78698 119395 80830 119490
rect 80998 119395 83130 119490
rect 83298 119395 85430 119490
rect 85598 119395 87730 119490
rect 87898 119395 90030 119490
rect 90198 119395 92330 119490
rect 92498 119395 94630 119490
rect 94798 119395 96930 119490
rect 97098 119395 99230 119490
rect 99398 119395 101530 119490
rect 101698 119395 103830 119490
rect 103998 119395 106130 119490
rect 106298 119395 108430 119490
rect 108598 119395 110730 119490
rect 110898 119395 113030 119490
rect 113198 119395 115330 119490
rect 115498 119395 117188 119490
rect 3056 856 117188 119395
rect 3166 734 5942 856
rect 6110 734 8886 856
rect 9054 734 11830 856
rect 11998 734 14774 856
rect 14942 734 17718 856
rect 17886 734 20662 856
rect 20830 734 23606 856
rect 23774 734 26550 856
rect 26718 734 29494 856
rect 29662 734 32438 856
rect 32606 734 35382 856
rect 35550 734 38326 856
rect 38494 734 41270 856
rect 41438 734 44214 856
rect 44382 734 47158 856
rect 47326 734 50102 856
rect 50270 734 53046 856
rect 53214 734 55990 856
rect 56158 734 58934 856
rect 59102 734 61878 856
rect 62046 734 64822 856
rect 64990 734 67766 856
rect 67934 734 70710 856
rect 70878 734 73654 856
rect 73822 734 76598 856
rect 76766 734 79542 856
rect 79710 734 82486 856
rect 82654 734 85430 856
rect 85598 734 88374 856
rect 88542 734 91318 856
rect 91486 734 94262 856
rect 94430 734 97206 856
rect 97374 734 100150 856
rect 100318 734 103094 856
rect 103262 734 106038 856
rect 106206 734 108982 856
rect 109150 734 111926 856
rect 112094 734 114870 856
rect 115038 734 117188 856
<< metal3 >>
rect 117307 114248 118107 114368
rect 117307 111528 118107 111648
rect 117307 108808 118107 108928
rect 117307 106088 118107 106208
rect 117307 103368 118107 103488
rect 117307 100648 118107 100768
rect 117307 97928 118107 98048
rect 117307 95208 118107 95328
rect 117307 92488 118107 92608
rect 117307 89768 118107 89888
rect 117307 87048 118107 87168
rect 117307 84328 118107 84448
rect 117307 81608 118107 81728
rect 117307 78888 118107 79008
rect 117307 76168 118107 76288
rect 117307 73448 118107 73568
rect 117307 70728 118107 70848
rect 117307 68008 118107 68128
rect 117307 65288 118107 65408
rect 117307 62568 118107 62688
rect 117307 59848 118107 59968
rect 117307 57128 118107 57248
rect 117307 54408 118107 54528
rect 117307 51688 118107 51808
rect 117307 48968 118107 49088
rect 117307 46248 118107 46368
rect 117307 43528 118107 43648
rect 117307 40808 118107 40928
rect 117307 38088 118107 38208
rect 117307 35368 118107 35488
rect 117307 32648 118107 32768
rect 117307 29928 118107 30048
rect 117307 27208 118107 27328
rect 117307 24488 118107 24608
rect 117307 21768 118107 21888
rect 117307 19048 118107 19168
rect 117307 16328 118107 16448
rect 117307 13608 118107 13728
rect 117307 10888 118107 11008
rect 117307 8168 118107 8288
rect 117307 5448 118107 5568
<< obsm3 >>
rect 4210 114448 117307 118285
rect 4210 114168 117227 114448
rect 4210 111728 117307 114168
rect 4210 111448 117227 111728
rect 4210 109008 117307 111448
rect 4210 108728 117227 109008
rect 4210 106288 117307 108728
rect 4210 106008 117227 106288
rect 4210 103568 117307 106008
rect 4210 103288 117227 103568
rect 4210 100848 117307 103288
rect 4210 100568 117227 100848
rect 4210 98128 117307 100568
rect 4210 97848 117227 98128
rect 4210 95408 117307 97848
rect 4210 95128 117227 95408
rect 4210 92688 117307 95128
rect 4210 92408 117227 92688
rect 4210 89968 117307 92408
rect 4210 89688 117227 89968
rect 4210 87248 117307 89688
rect 4210 86968 117227 87248
rect 4210 84528 117307 86968
rect 4210 84248 117227 84528
rect 4210 81808 117307 84248
rect 4210 81528 117227 81808
rect 4210 79088 117307 81528
rect 4210 78808 117227 79088
rect 4210 76368 117307 78808
rect 4210 76088 117227 76368
rect 4210 73648 117307 76088
rect 4210 73368 117227 73648
rect 4210 70928 117307 73368
rect 4210 70648 117227 70928
rect 4210 68208 117307 70648
rect 4210 67928 117227 68208
rect 4210 65488 117307 67928
rect 4210 65208 117227 65488
rect 4210 62768 117307 65208
rect 4210 62488 117227 62768
rect 4210 60048 117307 62488
rect 4210 59768 117227 60048
rect 4210 57328 117307 59768
rect 4210 57048 117227 57328
rect 4210 54608 117307 57048
rect 4210 54328 117227 54608
rect 4210 51888 117307 54328
rect 4210 51608 117227 51888
rect 4210 49168 117307 51608
rect 4210 48888 117227 49168
rect 4210 46448 117307 48888
rect 4210 46168 117227 46448
rect 4210 43728 117307 46168
rect 4210 43448 117227 43728
rect 4210 41008 117307 43448
rect 4210 40728 117227 41008
rect 4210 38288 117307 40728
rect 4210 38008 117227 38288
rect 4210 35568 117307 38008
rect 4210 35288 117227 35568
rect 4210 32848 117307 35288
rect 4210 32568 117227 32848
rect 4210 30128 117307 32568
rect 4210 29848 117227 30128
rect 4210 27408 117307 29848
rect 4210 27128 117227 27408
rect 4210 24688 117307 27128
rect 4210 24408 117227 24688
rect 4210 21968 117307 24408
rect 4210 21688 117227 21968
rect 4210 19248 117307 21688
rect 4210 18968 117227 19248
rect 4210 16528 117307 18968
rect 4210 16248 117227 16528
rect 4210 13808 117307 16248
rect 4210 13528 117227 13808
rect 4210 11088 117307 13528
rect 4210 10808 117227 11088
rect 4210 8368 117307 10808
rect 4210 8088 117227 8368
rect 4210 5648 117307 8088
rect 4210 5368 117227 5648
rect 4210 2143 117307 5368
<< metal4 >>
rect 4208 2128 4528 118096
rect 19568 2128 19888 118096
rect 34928 2128 35248 118096
rect 50288 2128 50608 118096
rect 65648 2128 65968 118096
rect 81008 2128 81328 118096
rect 96368 2128 96688 118096
rect 111728 2128 112048 118096
<< obsm4 >>
rect 8523 2619 19488 117469
rect 19968 2619 34848 117469
rect 35328 2619 50208 117469
rect 50688 2619 65568 117469
rect 66048 2619 80928 117469
rect 81408 2619 96288 117469
rect 96768 2619 111648 117469
rect 112128 2619 115309 117469
<< labels >>
rlabel metal2 s 115386 119451 115442 120251 6 i_clk
port 1 nsew signal input
rlabel metal3 s 117307 70728 118107 70848 6 i_debug_map_overlay
port 2 nsew signal input
rlabel metal3 s 117307 51688 118107 51808 6 i_debug_trace_overlay
port 3 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 i_debug_vec_overlay
port 4 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 i_gpout0_sel[0]
port 5 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 i_gpout0_sel[1]
port 6 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 i_gpout0_sel[2]
port 7 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 i_gpout0_sel[3]
port 8 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 i_gpout0_sel[4]
port 9 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 i_gpout0_sel[5]
port 10 nsew signal input
rlabel metal3 s 117307 19048 118107 19168 6 i_gpout1_sel[0]
port 11 nsew signal input
rlabel metal3 s 117307 21768 118107 21888 6 i_gpout1_sel[1]
port 12 nsew signal input
rlabel metal3 s 117307 24488 118107 24608 6 i_gpout1_sel[2]
port 13 nsew signal input
rlabel metal3 s 117307 27208 118107 27328 6 i_gpout1_sel[3]
port 14 nsew signal input
rlabel metal3 s 117307 29928 118107 30048 6 i_gpout1_sel[4]
port 15 nsew signal input
rlabel metal3 s 117307 32648 118107 32768 6 i_gpout1_sel[5]
port 16 nsew signal input
rlabel metal3 s 117307 35368 118107 35488 6 i_gpout2_sel[0]
port 17 nsew signal input
rlabel metal3 s 117307 38088 118107 38208 6 i_gpout2_sel[1]
port 18 nsew signal input
rlabel metal3 s 117307 40808 118107 40928 6 i_gpout2_sel[2]
port 19 nsew signal input
rlabel metal3 s 117307 43528 118107 43648 6 i_gpout2_sel[3]
port 20 nsew signal input
rlabel metal3 s 117307 46248 118107 46368 6 i_gpout2_sel[4]
port 21 nsew signal input
rlabel metal3 s 117307 48968 118107 49088 6 i_gpout2_sel[5]
port 22 nsew signal input
rlabel metal3 s 117307 54408 118107 54528 6 i_gpout3_sel[0]
port 23 nsew signal input
rlabel metal3 s 117307 57128 118107 57248 6 i_gpout3_sel[1]
port 24 nsew signal input
rlabel metal3 s 117307 59848 118107 59968 6 i_gpout3_sel[2]
port 25 nsew signal input
rlabel metal3 s 117307 62568 118107 62688 6 i_gpout3_sel[3]
port 26 nsew signal input
rlabel metal3 s 117307 65288 118107 65408 6 i_gpout3_sel[4]
port 27 nsew signal input
rlabel metal3 s 117307 68008 118107 68128 6 i_gpout3_sel[5]
port 28 nsew signal input
rlabel metal3 s 117307 73448 118107 73568 6 i_gpout4_sel[0]
port 29 nsew signal input
rlabel metal3 s 117307 76168 118107 76288 6 i_gpout4_sel[1]
port 30 nsew signal input
rlabel metal3 s 117307 78888 118107 79008 6 i_gpout4_sel[2]
port 31 nsew signal input
rlabel metal3 s 117307 81608 118107 81728 6 i_gpout4_sel[3]
port 32 nsew signal input
rlabel metal3 s 117307 84328 118107 84448 6 i_gpout4_sel[4]
port 33 nsew signal input
rlabel metal3 s 117307 87048 118107 87168 6 i_gpout4_sel[5]
port 34 nsew signal input
rlabel metal3 s 117307 89768 118107 89888 6 i_gpout5_sel[0]
port 35 nsew signal input
rlabel metal3 s 117307 92488 118107 92608 6 i_gpout5_sel[1]
port 36 nsew signal input
rlabel metal3 s 117307 95208 118107 95328 6 i_gpout5_sel[2]
port 37 nsew signal input
rlabel metal3 s 117307 97928 118107 98048 6 i_gpout5_sel[3]
port 38 nsew signal input
rlabel metal3 s 117307 100648 118107 100768 6 i_gpout5_sel[4]
port 39 nsew signal input
rlabel metal3 s 117307 103368 118107 103488 6 i_gpout5_sel[5]
port 40 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 i_la_invalid
port 41 nsew signal input
rlabel metal3 s 117307 106088 118107 106208 6 i_mode[0]
port 42 nsew signal input
rlabel metal3 s 117307 108808 118107 108928 6 i_mode[1]
port 43 nsew signal input
rlabel metal3 s 117307 111528 118107 111648 6 i_mode[2]
port 44 nsew signal input
rlabel metal3 s 117307 8168 118107 8288 6 i_reg_csb
port 45 nsew signal input
rlabel metal3 s 117307 10888 118107 11008 6 i_reg_mosi
port 46 nsew signal input
rlabel metal3 s 117307 13608 118107 13728 6 i_reg_outs_enb
port 47 nsew signal input
rlabel metal3 s 117307 16328 118107 16448 6 i_reg_sclk
port 48 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 i_reset_lock_a
port 49 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 i_reset_lock_b
port 50 nsew signal input
rlabel metal3 s 117307 114248 118107 114368 6 i_spare_0
port 51 nsew signal input
rlabel metal2 s 2686 119451 2742 120251 6 i_spare_1
port 52 nsew signal input
rlabel metal3 s 117307 5448 118107 5568 6 i_test_uc2
port 53 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 i_test_wci
port 54 nsew signal input
rlabel metal2 s 11886 119451 11942 120251 6 i_tex_in[0]
port 55 nsew signal input
rlabel metal2 s 9586 119451 9642 120251 6 i_tex_in[1]
port 56 nsew signal input
rlabel metal2 s 7286 119451 7342 120251 6 i_tex_in[2]
port 57 nsew signal input
rlabel metal2 s 4986 119451 5042 120251 6 i_tex_in[3]
port 58 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 i_vec_csb
port 59 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 i_vec_mosi
port 60 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 i_vec_sclk
port 61 nsew signal input
rlabel metal2 s 25686 119451 25742 120251 6 o_gpout[0]
port 62 nsew signal output
rlabel metal2 s 23386 119451 23442 120251 6 o_gpout[1]
port 63 nsew signal output
rlabel metal2 s 21086 119451 21142 120251 6 o_gpout[2]
port 64 nsew signal output
rlabel metal2 s 18786 119451 18842 120251 6 o_gpout[3]
port 65 nsew signal output
rlabel metal2 s 16486 119451 16542 120251 6 o_gpout[4]
port 66 nsew signal output
rlabel metal2 s 14186 119451 14242 120251 6 o_gpout[5]
port 67 nsew signal output
rlabel metal2 s 39486 119451 39542 120251 6 o_hsync
port 68 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 o_reset
port 69 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 o_rgb[0]
port 70 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 o_rgb[10]
port 71 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 o_rgb[11]
port 72 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 o_rgb[12]
port 73 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 o_rgb[13]
port 74 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 o_rgb[14]
port 75 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 o_rgb[15]
port 76 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 o_rgb[16]
port 77 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 o_rgb[17]
port 78 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 o_rgb[18]
port 79 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 o_rgb[19]
port 80 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 o_rgb[1]
port 81 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 o_rgb[20]
port 82 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 o_rgb[21]
port 83 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 o_rgb[22]
port 84 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 o_rgb[23]
port 85 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 o_rgb[2]
port 86 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 o_rgb[3]
port 87 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 o_rgb[4]
port 88 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 o_rgb[5]
port 89 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 o_rgb[6]
port 90 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 o_rgb[7]
port 91 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 o_rgb[8]
port 92 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 o_rgb[9]
port 93 nsew signal output
rlabel metal2 s 34886 119451 34942 120251 6 o_tex_csb
port 94 nsew signal output
rlabel metal2 s 32586 119451 32642 120251 6 o_tex_oeb0
port 95 nsew signal output
rlabel metal2 s 30286 119451 30342 120251 6 o_tex_out0
port 96 nsew signal output
rlabel metal2 s 27986 119451 28042 120251 6 o_tex_sclk
port 97 nsew signal output
rlabel metal2 s 37186 119451 37242 120251 6 o_vsync
port 98 nsew signal output
rlabel metal2 s 113086 119451 113142 120251 6 ones[0]
port 99 nsew signal output
rlabel metal2 s 90086 119451 90142 120251 6 ones[10]
port 100 nsew signal output
rlabel metal2 s 87786 119451 87842 120251 6 ones[11]
port 101 nsew signal output
rlabel metal2 s 85486 119451 85542 120251 6 ones[12]
port 102 nsew signal output
rlabel metal2 s 83186 119451 83242 120251 6 ones[13]
port 103 nsew signal output
rlabel metal2 s 80886 119451 80942 120251 6 ones[14]
port 104 nsew signal output
rlabel metal2 s 78586 119451 78642 120251 6 ones[15]
port 105 nsew signal output
rlabel metal2 s 110786 119451 110842 120251 6 ones[1]
port 106 nsew signal output
rlabel metal2 s 108486 119451 108542 120251 6 ones[2]
port 107 nsew signal output
rlabel metal2 s 106186 119451 106242 120251 6 ones[3]
port 108 nsew signal output
rlabel metal2 s 103886 119451 103942 120251 6 ones[4]
port 109 nsew signal output
rlabel metal2 s 101586 119451 101642 120251 6 ones[5]
port 110 nsew signal output
rlabel metal2 s 99286 119451 99342 120251 6 ones[6]
port 111 nsew signal output
rlabel metal2 s 96986 119451 97042 120251 6 ones[7]
port 112 nsew signal output
rlabel metal2 s 94686 119451 94742 120251 6 ones[8]
port 113 nsew signal output
rlabel metal2 s 92386 119451 92442 120251 6 ones[9]
port 114 nsew signal output
rlabel metal4 s 4208 2128 4528 118096 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 118096 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 118096 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 118096 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 118096 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 118096 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 118096 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 118096 6 vssd1
port 116 nsew ground bidirectional
rlabel metal2 s 76286 119451 76342 120251 6 zeros[0]
port 117 nsew signal output
rlabel metal2 s 53286 119451 53342 120251 6 zeros[10]
port 118 nsew signal output
rlabel metal2 s 50986 119451 51042 120251 6 zeros[11]
port 119 nsew signal output
rlabel metal2 s 48686 119451 48742 120251 6 zeros[12]
port 120 nsew signal output
rlabel metal2 s 46386 119451 46442 120251 6 zeros[13]
port 121 nsew signal output
rlabel metal2 s 44086 119451 44142 120251 6 zeros[14]
port 122 nsew signal output
rlabel metal2 s 41786 119451 41842 120251 6 zeros[15]
port 123 nsew signal output
rlabel metal2 s 73986 119451 74042 120251 6 zeros[1]
port 124 nsew signal output
rlabel metal2 s 71686 119451 71742 120251 6 zeros[2]
port 125 nsew signal output
rlabel metal2 s 69386 119451 69442 120251 6 zeros[3]
port 126 nsew signal output
rlabel metal2 s 67086 119451 67142 120251 6 zeros[4]
port 127 nsew signal output
rlabel metal2 s 64786 119451 64842 120251 6 zeros[5]
port 128 nsew signal output
rlabel metal2 s 62486 119451 62542 120251 6 zeros[6]
port 129 nsew signal output
rlabel metal2 s 60186 119451 60242 120251 6 zeros[7]
port 130 nsew signal output
rlabel metal2 s 57886 119451 57942 120251 6 zeros[8]
port 131 nsew signal output
rlabel metal2 s 55586 119451 55642 120251 6 zeros[9]
port 132 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 118107 120251
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 41325106
string GDS_FILE /home/zerotoasic/asic_tools/raybox-zero-caravel/openlane/top_ew_algofoogle/runs/23_11_06_12_28/results/signoff/top_ew_algofoogle.magic.gds
string GDS_START 1496174
<< end >>

