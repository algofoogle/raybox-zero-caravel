VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_ew_algofoogle
  CLASS BLOCK ;
  FOREIGN top_ew_algofoogle ;
  ORIGIN 0.000 0.000 ;
  SIZE 561.710 BY 572.430 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 14.320 561.710 14.920 ;
    END
  END i_clk
  PIN i_debug_map_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 342.760 561.710 343.360 ;
    END
  END i_debug_map_overlay
  PIN i_debug_trace_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 242.800 561.710 243.400 ;
    END
  END i_debug_trace_overlay
  PIN i_debug_vec_overlay
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END i_debug_vec_overlay
  PIN i_gpout0_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END i_gpout0_sel[0]
  PIN i_gpout0_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END i_gpout0_sel[1]
  PIN i_gpout0_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END i_gpout0_sel[2]
  PIN i_gpout0_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END i_gpout0_sel[3]
  PIN i_gpout0_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END i_gpout0_sel[4]
  PIN i_gpout0_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END i_gpout0_sel[5]
  PIN i_gpout1_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 71.440 561.710 72.040 ;
    END
  END i_gpout1_sel[0]
  PIN i_gpout1_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 85.720 561.710 86.320 ;
    END
  END i_gpout1_sel[1]
  PIN i_gpout1_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 100.000 561.710 100.600 ;
    END
  END i_gpout1_sel[2]
  PIN i_gpout1_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 114.280 561.710 114.880 ;
    END
  END i_gpout1_sel[3]
  PIN i_gpout1_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 128.560 561.710 129.160 ;
    END
  END i_gpout1_sel[4]
  PIN i_gpout1_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 142.840 561.710 143.440 ;
    END
  END i_gpout1_sel[5]
  PIN i_gpout2_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 157.120 561.710 157.720 ;
    END
  END i_gpout2_sel[0]
  PIN i_gpout2_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 171.400 561.710 172.000 ;
    END
  END i_gpout2_sel[1]
  PIN i_gpout2_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 185.680 561.710 186.280 ;
    END
  END i_gpout2_sel[2]
  PIN i_gpout2_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 199.960 561.710 200.560 ;
    END
  END i_gpout2_sel[3]
  PIN i_gpout2_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 214.240 561.710 214.840 ;
    END
  END i_gpout2_sel[4]
  PIN i_gpout2_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 228.520 561.710 229.120 ;
    END
  END i_gpout2_sel[5]
  PIN i_gpout3_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 257.080 561.710 257.680 ;
    END
  END i_gpout3_sel[0]
  PIN i_gpout3_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 271.360 561.710 271.960 ;
    END
  END i_gpout3_sel[1]
  PIN i_gpout3_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 285.640 561.710 286.240 ;
    END
  END i_gpout3_sel[2]
  PIN i_gpout3_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 299.920 561.710 300.520 ;
    END
  END i_gpout3_sel[3]
  PIN i_gpout3_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 314.200 561.710 314.800 ;
    END
  END i_gpout3_sel[4]
  PIN i_gpout3_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 328.480 561.710 329.080 ;
    END
  END i_gpout3_sel[5]
  PIN i_gpout4_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 357.040 561.710 357.640 ;
    END
  END i_gpout4_sel[0]
  PIN i_gpout4_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 371.320 561.710 371.920 ;
    END
  END i_gpout4_sel[1]
  PIN i_gpout4_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 385.600 561.710 386.200 ;
    END
  END i_gpout4_sel[2]
  PIN i_gpout4_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 399.880 561.710 400.480 ;
    END
  END i_gpout4_sel[3]
  PIN i_gpout4_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 414.160 561.710 414.760 ;
    END
  END i_gpout4_sel[4]
  PIN i_gpout4_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 428.440 561.710 429.040 ;
    END
  END i_gpout4_sel[5]
  PIN i_gpout5_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 442.720 561.710 443.320 ;
    END
  END i_gpout5_sel[0]
  PIN i_gpout5_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 457.000 561.710 457.600 ;
    END
  END i_gpout5_sel[1]
  PIN i_gpout5_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 471.280 561.710 471.880 ;
    END
  END i_gpout5_sel[2]
  PIN i_gpout5_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 485.560 561.710 486.160 ;
    END
  END i_gpout5_sel[3]
  PIN i_gpout5_sel[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 499.840 561.710 500.440 ;
    END
  END i_gpout5_sel[4]
  PIN i_gpout5_sel[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 514.120 561.710 514.720 ;
    END
  END i_gpout5_sel[5]
  PIN i_la_invalid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END i_la_invalid
  PIN i_mode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 528.400 561.710 529.000 ;
    END
  END i_mode[0]
  PIN i_mode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 542.680 561.710 543.280 ;
    END
  END i_mode[1]
  PIN i_mode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 556.960 561.710 557.560 ;
    END
  END i_mode[2]
  PIN i_reg_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 28.600 561.710 29.200 ;
    END
  END i_reg_csb
  PIN i_reg_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 42.880 561.710 43.480 ;
    END
  END i_reg_mosi
  PIN i_reg_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 557.710 57.160 561.710 57.760 ;
    END
  END i_reg_sclk
  PIN i_reset_lock_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END i_reset_lock_a
  PIN i_reset_lock_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END i_reset_lock_b
  PIN i_tex_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 568.430 44.990 572.430 ;
    END
  END i_tex_in[0]
  PIN i_tex_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 568.430 33.490 572.430 ;
    END
  END i_tex_in[1]
  PIN i_tex_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 568.430 21.990 572.430 ;
    END
  END i_tex_in[2]
  PIN i_tex_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 568.430 10.490 572.430 ;
    END
  END i_tex_in[3]
  PIN i_vec_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END i_vec_csb
  PIN i_vec_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END i_vec_mosi
  PIN i_vec_sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END i_vec_sclk
  PIN o_gpout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 568.430 113.990 572.430 ;
    END
  END o_gpout[0]
  PIN o_gpout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 568.430 102.490 572.430 ;
    END
  END o_gpout[1]
  PIN o_gpout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 568.430 90.990 572.430 ;
    END
  END o_gpout[2]
  PIN o_gpout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 568.430 79.490 572.430 ;
    END
  END o_gpout[3]
  PIN o_gpout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 568.430 67.990 572.430 ;
    END
  END o_gpout[4]
  PIN o_gpout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 568.430 56.490 572.430 ;
    END
  END o_gpout[5]
  PIN o_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 568.430 182.990 572.430 ;
    END
  END o_hsync
  PIN o_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END o_reset
  PIN o_rgb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END o_rgb[0]
  PIN o_rgb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END o_rgb[10]
  PIN o_rgb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END o_rgb[11]
  PIN o_rgb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END o_rgb[12]
  PIN o_rgb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END o_rgb[13]
  PIN o_rgb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END o_rgb[14]
  PIN o_rgb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END o_rgb[15]
  PIN o_rgb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END o_rgb[16]
  PIN o_rgb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END o_rgb[17]
  PIN o_rgb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END o_rgb[18]
  PIN o_rgb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END o_rgb[19]
  PIN o_rgb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END o_rgb[1]
  PIN o_rgb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END o_rgb[20]
  PIN o_rgb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END o_rgb[21]
  PIN o_rgb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END o_rgb[22]
  PIN o_rgb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END o_rgb[23]
  PIN o_rgb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END o_rgb[2]
  PIN o_rgb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END o_rgb[3]
  PIN o_rgb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END o_rgb[4]
  PIN o_rgb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END o_rgb[5]
  PIN o_rgb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END o_rgb[6]
  PIN o_rgb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END o_rgb[7]
  PIN o_rgb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END o_rgb[8]
  PIN o_rgb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END o_rgb[9]
  PIN o_tex_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 568.430 159.990 572.430 ;
    END
  END o_tex_csb
  PIN o_tex_oeb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 568.430 148.490 572.430 ;
    END
  END o_tex_oeb0
  PIN o_tex_out0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 568.430 136.990 572.430 ;
    END
  END o_tex_out0
  PIN o_tex_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 568.430 125.490 572.430 ;
    END
  END o_tex_sclk
  PIN o_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 568.430 171.490 572.430 ;
    END
  END o_vsync
  PIN ones[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 568.430 550.990 572.430 ;
    END
  END ones[0]
  PIN ones[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 568.430 435.990 572.430 ;
    END
  END ones[10]
  PIN ones[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 568.430 424.490 572.430 ;
    END
  END ones[11]
  PIN ones[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 568.430 412.990 572.430 ;
    END
  END ones[12]
  PIN ones[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 568.430 401.490 572.430 ;
    END
  END ones[13]
  PIN ones[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 568.430 389.990 572.430 ;
    END
  END ones[14]
  PIN ones[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 568.430 378.490 572.430 ;
    END
  END ones[15]
  PIN ones[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 568.430 539.490 572.430 ;
    END
  END ones[1]
  PIN ones[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 568.430 527.990 572.430 ;
    END
  END ones[2]
  PIN ones[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 568.430 516.490 572.430 ;
    END
  END ones[3]
  PIN ones[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 568.430 504.990 572.430 ;
    END
  END ones[4]
  PIN ones[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 568.430 493.490 572.430 ;
    END
  END ones[5]
  PIN ones[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 568.430 481.990 572.430 ;
    END
  END ones[6]
  PIN ones[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 568.430 470.490 572.430 ;
    END
  END ones[7]
  PIN ones[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 568.430 458.990 572.430 ;
    END
  END ones[8]
  PIN ones[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 568.430 447.490 572.430 ;
    END
  END ones[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 560.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 560.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 560.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 560.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 560.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 560.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 560.560 ;
    END
  END vssd1
  PIN zeros[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 568.430 366.990 572.430 ;
    END
  END zeros[0]
  PIN zeros[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 568.430 251.990 572.430 ;
    END
  END zeros[10]
  PIN zeros[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 568.430 240.490 572.430 ;
    END
  END zeros[11]
  PIN zeros[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 568.430 228.990 572.430 ;
    END
  END zeros[12]
  PIN zeros[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 568.430 217.490 572.430 ;
    END
  END zeros[13]
  PIN zeros[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 568.430 205.990 572.430 ;
    END
  END zeros[14]
  PIN zeros[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 568.430 194.490 572.430 ;
    END
  END zeros[15]
  PIN zeros[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 568.430 355.490 572.430 ;
    END
  END zeros[1]
  PIN zeros[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 568.430 343.990 572.430 ;
    END
  END zeros[2]
  PIN zeros[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 568.430 332.490 572.430 ;
    END
  END zeros[3]
  PIN zeros[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 568.430 320.990 572.430 ;
    END
  END zeros[4]
  PIN zeros[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 568.430 309.490 572.430 ;
    END
  END zeros[5]
  PIN zeros[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 568.430 297.990 572.430 ;
    END
  END zeros[6]
  PIN zeros[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 568.430 286.490 572.430 ;
    END
  END zeros[7]
  PIN zeros[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 568.430 274.990 572.430 ;
    END
  END zeros[8]
  PIN zeros[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 568.430 263.490 572.430 ;
    END
  END zeros[9]
  OBS
      LAYER nwell ;
        RECT 5.330 556.185 556.330 559.015 ;
        RECT 5.330 550.745 556.330 553.575 ;
        RECT 5.330 545.305 556.330 548.135 ;
        RECT 5.330 539.865 556.330 542.695 ;
        RECT 5.330 534.425 556.330 537.255 ;
        RECT 5.330 528.985 556.330 531.815 ;
        RECT 5.330 523.545 556.330 526.375 ;
        RECT 5.330 518.105 556.330 520.935 ;
        RECT 5.330 512.665 556.330 515.495 ;
        RECT 5.330 507.225 556.330 510.055 ;
        RECT 5.330 501.785 556.330 504.615 ;
        RECT 5.330 496.345 556.330 499.175 ;
        RECT 5.330 490.905 556.330 493.735 ;
        RECT 5.330 485.465 556.330 488.295 ;
        RECT 5.330 480.025 556.330 482.855 ;
        RECT 5.330 474.585 556.330 477.415 ;
        RECT 5.330 469.145 556.330 471.975 ;
        RECT 5.330 463.705 556.330 466.535 ;
        RECT 5.330 458.265 556.330 461.095 ;
        RECT 5.330 452.825 556.330 455.655 ;
        RECT 5.330 447.385 556.330 450.215 ;
        RECT 5.330 441.945 556.330 444.775 ;
        RECT 5.330 436.505 556.330 439.335 ;
        RECT 5.330 431.065 556.330 433.895 ;
        RECT 5.330 425.625 556.330 428.455 ;
        RECT 5.330 420.185 556.330 423.015 ;
        RECT 5.330 414.745 556.330 417.575 ;
        RECT 5.330 409.305 556.330 412.135 ;
        RECT 5.330 403.865 556.330 406.695 ;
        RECT 5.330 398.425 556.330 401.255 ;
        RECT 5.330 392.985 556.330 395.815 ;
        RECT 5.330 387.545 556.330 390.375 ;
        RECT 5.330 382.105 556.330 384.935 ;
        RECT 5.330 376.665 556.330 379.495 ;
        RECT 5.330 371.225 556.330 374.055 ;
        RECT 5.330 365.785 556.330 368.615 ;
        RECT 5.330 360.345 556.330 363.175 ;
        RECT 5.330 354.905 556.330 357.735 ;
        RECT 5.330 349.465 556.330 352.295 ;
        RECT 5.330 344.025 556.330 346.855 ;
        RECT 5.330 338.585 556.330 341.415 ;
        RECT 5.330 333.145 556.330 335.975 ;
        RECT 5.330 327.705 556.330 330.535 ;
        RECT 5.330 322.265 556.330 325.095 ;
        RECT 5.330 316.825 556.330 319.655 ;
        RECT 5.330 311.385 556.330 314.215 ;
        RECT 5.330 305.945 556.330 308.775 ;
        RECT 5.330 300.505 556.330 303.335 ;
        RECT 5.330 295.065 556.330 297.895 ;
        RECT 5.330 289.625 556.330 292.455 ;
        RECT 5.330 284.185 556.330 287.015 ;
        RECT 5.330 278.745 556.330 281.575 ;
        RECT 5.330 273.305 556.330 276.135 ;
        RECT 5.330 267.865 556.330 270.695 ;
        RECT 5.330 262.425 556.330 265.255 ;
        RECT 5.330 256.985 556.330 259.815 ;
        RECT 5.330 251.545 556.330 254.375 ;
        RECT 5.330 246.105 556.330 248.935 ;
        RECT 5.330 240.665 556.330 243.495 ;
        RECT 5.330 235.225 556.330 238.055 ;
        RECT 5.330 229.785 556.330 232.615 ;
        RECT 5.330 224.345 556.330 227.175 ;
        RECT 5.330 218.905 556.330 221.735 ;
        RECT 5.330 213.465 556.330 216.295 ;
        RECT 5.330 208.025 556.330 210.855 ;
        RECT 5.330 202.585 556.330 205.415 ;
        RECT 5.330 197.145 556.330 199.975 ;
        RECT 5.330 191.705 556.330 194.535 ;
        RECT 5.330 186.265 556.330 189.095 ;
        RECT 5.330 180.825 556.330 183.655 ;
        RECT 5.330 175.385 556.330 178.215 ;
        RECT 5.330 169.945 556.330 172.775 ;
        RECT 5.330 164.505 556.330 167.335 ;
        RECT 5.330 159.065 556.330 161.895 ;
        RECT 5.330 153.625 556.330 156.455 ;
        RECT 5.330 148.185 556.330 151.015 ;
        RECT 5.330 142.745 556.330 145.575 ;
        RECT 5.330 137.305 556.330 140.135 ;
        RECT 5.330 131.865 556.330 134.695 ;
        RECT 5.330 126.425 556.330 129.255 ;
        RECT 5.330 120.985 556.330 123.815 ;
        RECT 5.330 115.545 556.330 118.375 ;
        RECT 5.330 110.105 556.330 112.935 ;
        RECT 5.330 104.665 556.330 107.495 ;
        RECT 5.330 99.225 556.330 102.055 ;
        RECT 5.330 93.785 556.330 96.615 ;
        RECT 5.330 88.345 556.330 91.175 ;
        RECT 5.330 82.905 556.330 85.735 ;
        RECT 5.330 77.465 556.330 80.295 ;
        RECT 5.330 72.025 556.330 74.855 ;
        RECT 5.330 66.585 556.330 69.415 ;
        RECT 5.330 61.145 556.330 63.975 ;
        RECT 5.330 55.705 556.330 58.535 ;
        RECT 5.330 50.265 556.330 53.095 ;
        RECT 5.330 44.825 556.330 47.655 ;
        RECT 5.330 39.385 556.330 42.215 ;
        RECT 5.330 33.945 556.330 36.775 ;
        RECT 5.330 28.505 556.330 31.335 ;
        RECT 5.330 23.065 556.330 25.895 ;
        RECT 5.330 17.625 556.330 20.455 ;
        RECT 5.330 12.185 556.330 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 556.140 560.405 ;
      LAYER met1 ;
        RECT 5.520 9.560 556.140 560.560 ;
      LAYER met2 ;
        RECT 8.380 568.150 9.930 568.890 ;
        RECT 10.770 568.150 21.430 568.890 ;
        RECT 22.270 568.150 32.930 568.890 ;
        RECT 33.770 568.150 44.430 568.890 ;
        RECT 45.270 568.150 55.930 568.890 ;
        RECT 56.770 568.150 67.430 568.890 ;
        RECT 68.270 568.150 78.930 568.890 ;
        RECT 79.770 568.150 90.430 568.890 ;
        RECT 91.270 568.150 101.930 568.890 ;
        RECT 102.770 568.150 113.430 568.890 ;
        RECT 114.270 568.150 124.930 568.890 ;
        RECT 125.770 568.150 136.430 568.890 ;
        RECT 137.270 568.150 147.930 568.890 ;
        RECT 148.770 568.150 159.430 568.890 ;
        RECT 160.270 568.150 170.930 568.890 ;
        RECT 171.770 568.150 182.430 568.890 ;
        RECT 183.270 568.150 193.930 568.890 ;
        RECT 194.770 568.150 205.430 568.890 ;
        RECT 206.270 568.150 216.930 568.890 ;
        RECT 217.770 568.150 228.430 568.890 ;
        RECT 229.270 568.150 239.930 568.890 ;
        RECT 240.770 568.150 251.430 568.890 ;
        RECT 252.270 568.150 262.930 568.890 ;
        RECT 263.770 568.150 274.430 568.890 ;
        RECT 275.270 568.150 285.930 568.890 ;
        RECT 286.770 568.150 297.430 568.890 ;
        RECT 298.270 568.150 308.930 568.890 ;
        RECT 309.770 568.150 320.430 568.890 ;
        RECT 321.270 568.150 331.930 568.890 ;
        RECT 332.770 568.150 343.430 568.890 ;
        RECT 344.270 568.150 354.930 568.890 ;
        RECT 355.770 568.150 366.430 568.890 ;
        RECT 367.270 568.150 377.930 568.890 ;
        RECT 378.770 568.150 389.430 568.890 ;
        RECT 390.270 568.150 400.930 568.890 ;
        RECT 401.770 568.150 412.430 568.890 ;
        RECT 413.270 568.150 423.930 568.890 ;
        RECT 424.770 568.150 435.430 568.890 ;
        RECT 436.270 568.150 446.930 568.890 ;
        RECT 447.770 568.150 458.430 568.890 ;
        RECT 459.270 568.150 469.930 568.890 ;
        RECT 470.770 568.150 481.430 568.890 ;
        RECT 482.270 568.150 492.930 568.890 ;
        RECT 493.770 568.150 504.430 568.890 ;
        RECT 505.270 568.150 515.930 568.890 ;
        RECT 516.770 568.150 527.430 568.890 ;
        RECT 528.270 568.150 538.930 568.890 ;
        RECT 539.770 568.150 550.430 568.890 ;
        RECT 551.270 568.150 554.660 568.890 ;
        RECT 8.380 4.280 554.660 568.150 ;
        RECT 8.930 3.670 22.810 4.280 ;
        RECT 23.650 3.670 37.530 4.280 ;
        RECT 38.370 3.670 52.250 4.280 ;
        RECT 53.090 3.670 66.970 4.280 ;
        RECT 67.810 3.670 81.690 4.280 ;
        RECT 82.530 3.670 96.410 4.280 ;
        RECT 97.250 3.670 111.130 4.280 ;
        RECT 111.970 3.670 125.850 4.280 ;
        RECT 126.690 3.670 140.570 4.280 ;
        RECT 141.410 3.670 155.290 4.280 ;
        RECT 156.130 3.670 170.010 4.280 ;
        RECT 170.850 3.670 184.730 4.280 ;
        RECT 185.570 3.670 199.450 4.280 ;
        RECT 200.290 3.670 214.170 4.280 ;
        RECT 215.010 3.670 228.890 4.280 ;
        RECT 229.730 3.670 243.610 4.280 ;
        RECT 244.450 3.670 258.330 4.280 ;
        RECT 259.170 3.670 273.050 4.280 ;
        RECT 273.890 3.670 287.770 4.280 ;
        RECT 288.610 3.670 302.490 4.280 ;
        RECT 303.330 3.670 317.210 4.280 ;
        RECT 318.050 3.670 331.930 4.280 ;
        RECT 332.770 3.670 346.650 4.280 ;
        RECT 347.490 3.670 361.370 4.280 ;
        RECT 362.210 3.670 376.090 4.280 ;
        RECT 376.930 3.670 390.810 4.280 ;
        RECT 391.650 3.670 405.530 4.280 ;
        RECT 406.370 3.670 420.250 4.280 ;
        RECT 421.090 3.670 434.970 4.280 ;
        RECT 435.810 3.670 449.690 4.280 ;
        RECT 450.530 3.670 464.410 4.280 ;
        RECT 465.250 3.670 479.130 4.280 ;
        RECT 479.970 3.670 493.850 4.280 ;
        RECT 494.690 3.670 508.570 4.280 ;
        RECT 509.410 3.670 523.290 4.280 ;
        RECT 524.130 3.670 538.010 4.280 ;
        RECT 538.850 3.670 552.730 4.280 ;
        RECT 553.570 3.670 554.660 4.280 ;
      LAYER met3 ;
        RECT 21.050 557.960 557.710 560.485 ;
        RECT 21.050 556.560 557.310 557.960 ;
        RECT 21.050 543.680 557.710 556.560 ;
        RECT 21.050 542.280 557.310 543.680 ;
        RECT 21.050 529.400 557.710 542.280 ;
        RECT 21.050 528.000 557.310 529.400 ;
        RECT 21.050 515.120 557.710 528.000 ;
        RECT 21.050 513.720 557.310 515.120 ;
        RECT 21.050 500.840 557.710 513.720 ;
        RECT 21.050 499.440 557.310 500.840 ;
        RECT 21.050 486.560 557.710 499.440 ;
        RECT 21.050 485.160 557.310 486.560 ;
        RECT 21.050 472.280 557.710 485.160 ;
        RECT 21.050 470.880 557.310 472.280 ;
        RECT 21.050 458.000 557.710 470.880 ;
        RECT 21.050 456.600 557.310 458.000 ;
        RECT 21.050 443.720 557.710 456.600 ;
        RECT 21.050 442.320 557.310 443.720 ;
        RECT 21.050 429.440 557.710 442.320 ;
        RECT 21.050 428.040 557.310 429.440 ;
        RECT 21.050 415.160 557.710 428.040 ;
        RECT 21.050 413.760 557.310 415.160 ;
        RECT 21.050 400.880 557.710 413.760 ;
        RECT 21.050 399.480 557.310 400.880 ;
        RECT 21.050 386.600 557.710 399.480 ;
        RECT 21.050 385.200 557.310 386.600 ;
        RECT 21.050 372.320 557.710 385.200 ;
        RECT 21.050 370.920 557.310 372.320 ;
        RECT 21.050 358.040 557.710 370.920 ;
        RECT 21.050 356.640 557.310 358.040 ;
        RECT 21.050 343.760 557.710 356.640 ;
        RECT 21.050 342.360 557.310 343.760 ;
        RECT 21.050 329.480 557.710 342.360 ;
        RECT 21.050 328.080 557.310 329.480 ;
        RECT 21.050 315.200 557.710 328.080 ;
        RECT 21.050 313.800 557.310 315.200 ;
        RECT 21.050 300.920 557.710 313.800 ;
        RECT 21.050 299.520 557.310 300.920 ;
        RECT 21.050 286.640 557.710 299.520 ;
        RECT 21.050 285.240 557.310 286.640 ;
        RECT 21.050 272.360 557.710 285.240 ;
        RECT 21.050 270.960 557.310 272.360 ;
        RECT 21.050 258.080 557.710 270.960 ;
        RECT 21.050 256.680 557.310 258.080 ;
        RECT 21.050 243.800 557.710 256.680 ;
        RECT 21.050 242.400 557.310 243.800 ;
        RECT 21.050 229.520 557.710 242.400 ;
        RECT 21.050 228.120 557.310 229.520 ;
        RECT 21.050 215.240 557.710 228.120 ;
        RECT 21.050 213.840 557.310 215.240 ;
        RECT 21.050 200.960 557.710 213.840 ;
        RECT 21.050 199.560 557.310 200.960 ;
        RECT 21.050 186.680 557.710 199.560 ;
        RECT 21.050 185.280 557.310 186.680 ;
        RECT 21.050 172.400 557.710 185.280 ;
        RECT 21.050 171.000 557.310 172.400 ;
        RECT 21.050 158.120 557.710 171.000 ;
        RECT 21.050 156.720 557.310 158.120 ;
        RECT 21.050 143.840 557.710 156.720 ;
        RECT 21.050 142.440 557.310 143.840 ;
        RECT 21.050 129.560 557.710 142.440 ;
        RECT 21.050 128.160 557.310 129.560 ;
        RECT 21.050 115.280 557.710 128.160 ;
        RECT 21.050 113.880 557.310 115.280 ;
        RECT 21.050 101.000 557.710 113.880 ;
        RECT 21.050 99.600 557.310 101.000 ;
        RECT 21.050 86.720 557.710 99.600 ;
        RECT 21.050 85.320 557.310 86.720 ;
        RECT 21.050 72.440 557.710 85.320 ;
        RECT 21.050 71.040 557.310 72.440 ;
        RECT 21.050 58.160 557.710 71.040 ;
        RECT 21.050 56.760 557.310 58.160 ;
        RECT 21.050 43.880 557.710 56.760 ;
        RECT 21.050 42.480 557.310 43.880 ;
        RECT 21.050 29.600 557.710 42.480 ;
        RECT 21.050 28.200 557.310 29.600 ;
        RECT 21.050 15.320 557.710 28.200 ;
        RECT 21.050 13.920 557.310 15.320 ;
        RECT 21.050 10.715 557.710 13.920 ;
      LAYER met4 ;
        RECT 115.295 12.415 174.240 559.465 ;
        RECT 176.640 12.415 251.040 559.465 ;
        RECT 253.440 12.415 327.840 559.465 ;
        RECT 330.240 12.415 404.640 559.465 ;
        RECT 407.040 12.415 481.440 559.465 ;
        RECT 483.840 12.415 489.145 559.465 ;
  END
END top_ew_algofoogle
END LIBRARY

