// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_outs_enb,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_spare_0,
    i_spare_1,
    i_test_uc2,
    i_test_wci,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_outs_enb;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_spare_0;
 input i_spare_1;
 input i_test_uc2;
 input i_test_wci;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire _00000_;
 wire _00001_;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire clknet_leaf_0_i_clk;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net78;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net79;
 wire net94;
 wire net95;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net112;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdx[5] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_mapdy[5] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.side_hot ;
 wire \rbzero.spi_registers.buf_floor[0] ;
 wire \rbzero.spi_registers.buf_floor[1] ;
 wire \rbzero.spi_registers.buf_floor[2] ;
 wire \rbzero.spi_registers.buf_floor[3] ;
 wire \rbzero.spi_registers.buf_floor[4] ;
 wire \rbzero.spi_registers.buf_floor[5] ;
 wire \rbzero.spi_registers.buf_leak[0] ;
 wire \rbzero.spi_registers.buf_leak[1] ;
 wire \rbzero.spi_registers.buf_leak[2] ;
 wire \rbzero.spi_registers.buf_leak[3] ;
 wire \rbzero.spi_registers.buf_leak[4] ;
 wire \rbzero.spi_registers.buf_leak[5] ;
 wire \rbzero.spi_registers.buf_mapdx[0] ;
 wire \rbzero.spi_registers.buf_mapdx[1] ;
 wire \rbzero.spi_registers.buf_mapdx[2] ;
 wire \rbzero.spi_registers.buf_mapdx[3] ;
 wire \rbzero.spi_registers.buf_mapdx[4] ;
 wire \rbzero.spi_registers.buf_mapdx[5] ;
 wire \rbzero.spi_registers.buf_mapdxw[0] ;
 wire \rbzero.spi_registers.buf_mapdxw[1] ;
 wire \rbzero.spi_registers.buf_mapdy[0] ;
 wire \rbzero.spi_registers.buf_mapdy[1] ;
 wire \rbzero.spi_registers.buf_mapdy[2] ;
 wire \rbzero.spi_registers.buf_mapdy[3] ;
 wire \rbzero.spi_registers.buf_mapdy[4] ;
 wire \rbzero.spi_registers.buf_mapdy[5] ;
 wire \rbzero.spi_registers.buf_mapdyw[0] ;
 wire \rbzero.spi_registers.buf_mapdyw[1] ;
 wire \rbzero.spi_registers.buf_otherx[0] ;
 wire \rbzero.spi_registers.buf_otherx[1] ;
 wire \rbzero.spi_registers.buf_otherx[2] ;
 wire \rbzero.spi_registers.buf_otherx[3] ;
 wire \rbzero.spi_registers.buf_otherx[4] ;
 wire \rbzero.spi_registers.buf_othery[0] ;
 wire \rbzero.spi_registers.buf_othery[1] ;
 wire \rbzero.spi_registers.buf_othery[2] ;
 wire \rbzero.spi_registers.buf_othery[3] ;
 wire \rbzero.spi_registers.buf_othery[4] ;
 wire \rbzero.spi_registers.buf_sky[0] ;
 wire \rbzero.spi_registers.buf_sky[1] ;
 wire \rbzero.spi_registers.buf_sky[2] ;
 wire \rbzero.spi_registers.buf_sky[3] ;
 wire \rbzero.spi_registers.buf_sky[4] ;
 wire \rbzero.spi_registers.buf_sky[5] ;
 wire \rbzero.spi_registers.buf_texadd0[0] ;
 wire \rbzero.spi_registers.buf_texadd0[10] ;
 wire \rbzero.spi_registers.buf_texadd0[11] ;
 wire \rbzero.spi_registers.buf_texadd0[12] ;
 wire \rbzero.spi_registers.buf_texadd0[13] ;
 wire \rbzero.spi_registers.buf_texadd0[14] ;
 wire \rbzero.spi_registers.buf_texadd0[15] ;
 wire \rbzero.spi_registers.buf_texadd0[16] ;
 wire \rbzero.spi_registers.buf_texadd0[17] ;
 wire \rbzero.spi_registers.buf_texadd0[18] ;
 wire \rbzero.spi_registers.buf_texadd0[19] ;
 wire \rbzero.spi_registers.buf_texadd0[1] ;
 wire \rbzero.spi_registers.buf_texadd0[20] ;
 wire \rbzero.spi_registers.buf_texadd0[21] ;
 wire \rbzero.spi_registers.buf_texadd0[22] ;
 wire \rbzero.spi_registers.buf_texadd0[23] ;
 wire \rbzero.spi_registers.buf_texadd0[2] ;
 wire \rbzero.spi_registers.buf_texadd0[3] ;
 wire \rbzero.spi_registers.buf_texadd0[4] ;
 wire \rbzero.spi_registers.buf_texadd0[5] ;
 wire \rbzero.spi_registers.buf_texadd0[6] ;
 wire \rbzero.spi_registers.buf_texadd0[7] ;
 wire \rbzero.spi_registers.buf_texadd0[8] ;
 wire \rbzero.spi_registers.buf_texadd0[9] ;
 wire \rbzero.spi_registers.buf_texadd1[0] ;
 wire \rbzero.spi_registers.buf_texadd1[10] ;
 wire \rbzero.spi_registers.buf_texadd1[11] ;
 wire \rbzero.spi_registers.buf_texadd1[12] ;
 wire \rbzero.spi_registers.buf_texadd1[13] ;
 wire \rbzero.spi_registers.buf_texadd1[14] ;
 wire \rbzero.spi_registers.buf_texadd1[15] ;
 wire \rbzero.spi_registers.buf_texadd1[16] ;
 wire \rbzero.spi_registers.buf_texadd1[17] ;
 wire \rbzero.spi_registers.buf_texadd1[18] ;
 wire \rbzero.spi_registers.buf_texadd1[19] ;
 wire \rbzero.spi_registers.buf_texadd1[1] ;
 wire \rbzero.spi_registers.buf_texadd1[20] ;
 wire \rbzero.spi_registers.buf_texadd1[21] ;
 wire \rbzero.spi_registers.buf_texadd1[22] ;
 wire \rbzero.spi_registers.buf_texadd1[23] ;
 wire \rbzero.spi_registers.buf_texadd1[2] ;
 wire \rbzero.spi_registers.buf_texadd1[3] ;
 wire \rbzero.spi_registers.buf_texadd1[4] ;
 wire \rbzero.spi_registers.buf_texadd1[5] ;
 wire \rbzero.spi_registers.buf_texadd1[6] ;
 wire \rbzero.spi_registers.buf_texadd1[7] ;
 wire \rbzero.spi_registers.buf_texadd1[8] ;
 wire \rbzero.spi_registers.buf_texadd1[9] ;
 wire \rbzero.spi_registers.buf_texadd2[0] ;
 wire \rbzero.spi_registers.buf_texadd2[10] ;
 wire \rbzero.spi_registers.buf_texadd2[11] ;
 wire \rbzero.spi_registers.buf_texadd2[12] ;
 wire \rbzero.spi_registers.buf_texadd2[13] ;
 wire \rbzero.spi_registers.buf_texadd2[14] ;
 wire \rbzero.spi_registers.buf_texadd2[15] ;
 wire \rbzero.spi_registers.buf_texadd2[16] ;
 wire \rbzero.spi_registers.buf_texadd2[17] ;
 wire \rbzero.spi_registers.buf_texadd2[18] ;
 wire \rbzero.spi_registers.buf_texadd2[19] ;
 wire \rbzero.spi_registers.buf_texadd2[1] ;
 wire \rbzero.spi_registers.buf_texadd2[20] ;
 wire \rbzero.spi_registers.buf_texadd2[21] ;
 wire \rbzero.spi_registers.buf_texadd2[22] ;
 wire \rbzero.spi_registers.buf_texadd2[23] ;
 wire \rbzero.spi_registers.buf_texadd2[2] ;
 wire \rbzero.spi_registers.buf_texadd2[3] ;
 wire \rbzero.spi_registers.buf_texadd2[4] ;
 wire \rbzero.spi_registers.buf_texadd2[5] ;
 wire \rbzero.spi_registers.buf_texadd2[6] ;
 wire \rbzero.spi_registers.buf_texadd2[7] ;
 wire \rbzero.spi_registers.buf_texadd2[8] ;
 wire \rbzero.spi_registers.buf_texadd2[9] ;
 wire \rbzero.spi_registers.buf_texadd3[0] ;
 wire \rbzero.spi_registers.buf_texadd3[10] ;
 wire \rbzero.spi_registers.buf_texadd3[11] ;
 wire \rbzero.spi_registers.buf_texadd3[12] ;
 wire \rbzero.spi_registers.buf_texadd3[13] ;
 wire \rbzero.spi_registers.buf_texadd3[14] ;
 wire \rbzero.spi_registers.buf_texadd3[15] ;
 wire \rbzero.spi_registers.buf_texadd3[16] ;
 wire \rbzero.spi_registers.buf_texadd3[17] ;
 wire \rbzero.spi_registers.buf_texadd3[18] ;
 wire \rbzero.spi_registers.buf_texadd3[19] ;
 wire \rbzero.spi_registers.buf_texadd3[1] ;
 wire \rbzero.spi_registers.buf_texadd3[20] ;
 wire \rbzero.spi_registers.buf_texadd3[21] ;
 wire \rbzero.spi_registers.buf_texadd3[22] ;
 wire \rbzero.spi_registers.buf_texadd3[23] ;
 wire \rbzero.spi_registers.buf_texadd3[2] ;
 wire \rbzero.spi_registers.buf_texadd3[3] ;
 wire \rbzero.spi_registers.buf_texadd3[4] ;
 wire \rbzero.spi_registers.buf_texadd3[5] ;
 wire \rbzero.spi_registers.buf_texadd3[6] ;
 wire \rbzero.spi_registers.buf_texadd3[7] ;
 wire \rbzero.spi_registers.buf_texadd3[8] ;
 wire \rbzero.spi_registers.buf_texadd3[9] ;
 wire \rbzero.spi_registers.buf_vinf ;
 wire \rbzero.spi_registers.buf_vshift[0] ;
 wire \rbzero.spi_registers.buf_vshift[1] ;
 wire \rbzero.spi_registers.buf_vshift[2] ;
 wire \rbzero.spi_registers.buf_vshift[3] ;
 wire \rbzero.spi_registers.buf_vshift[4] ;
 wire \rbzero.spi_registers.buf_vshift[5] ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[16] ;
 wire \rbzero.spi_registers.spi_buffer[17] ;
 wire \rbzero.spi_registers.spi_buffer[18] ;
 wire \rbzero.spi_registers.spi_buffer[19] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[20] ;
 wire \rbzero.spi_registers.spi_buffer[21] ;
 wire \rbzero.spi_registers.spi_buffer[22] ;
 wire \rbzero.spi_registers.spi_buffer[23] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.texadd0[0] ;
 wire \rbzero.spi_registers.texadd0[10] ;
 wire \rbzero.spi_registers.texadd0[11] ;
 wire \rbzero.spi_registers.texadd0[12] ;
 wire \rbzero.spi_registers.texadd0[13] ;
 wire \rbzero.spi_registers.texadd0[14] ;
 wire \rbzero.spi_registers.texadd0[15] ;
 wire \rbzero.spi_registers.texadd0[16] ;
 wire \rbzero.spi_registers.texadd0[17] ;
 wire \rbzero.spi_registers.texadd0[18] ;
 wire \rbzero.spi_registers.texadd0[19] ;
 wire \rbzero.spi_registers.texadd0[1] ;
 wire \rbzero.spi_registers.texadd0[20] ;
 wire \rbzero.spi_registers.texadd0[21] ;
 wire \rbzero.spi_registers.texadd0[22] ;
 wire \rbzero.spi_registers.texadd0[23] ;
 wire \rbzero.spi_registers.texadd0[2] ;
 wire \rbzero.spi_registers.texadd0[3] ;
 wire \rbzero.spi_registers.texadd0[4] ;
 wire \rbzero.spi_registers.texadd0[5] ;
 wire \rbzero.spi_registers.texadd0[6] ;
 wire \rbzero.spi_registers.texadd0[7] ;
 wire \rbzero.spi_registers.texadd0[8] ;
 wire \rbzero.spi_registers.texadd0[9] ;
 wire \rbzero.spi_registers.texadd1[0] ;
 wire \rbzero.spi_registers.texadd1[10] ;
 wire \rbzero.spi_registers.texadd1[11] ;
 wire \rbzero.spi_registers.texadd1[12] ;
 wire \rbzero.spi_registers.texadd1[13] ;
 wire \rbzero.spi_registers.texadd1[14] ;
 wire \rbzero.spi_registers.texadd1[15] ;
 wire \rbzero.spi_registers.texadd1[16] ;
 wire \rbzero.spi_registers.texadd1[17] ;
 wire \rbzero.spi_registers.texadd1[18] ;
 wire \rbzero.spi_registers.texadd1[19] ;
 wire \rbzero.spi_registers.texadd1[1] ;
 wire \rbzero.spi_registers.texadd1[20] ;
 wire \rbzero.spi_registers.texadd1[21] ;
 wire \rbzero.spi_registers.texadd1[22] ;
 wire \rbzero.spi_registers.texadd1[23] ;
 wire \rbzero.spi_registers.texadd1[2] ;
 wire \rbzero.spi_registers.texadd1[3] ;
 wire \rbzero.spi_registers.texadd1[4] ;
 wire \rbzero.spi_registers.texadd1[5] ;
 wire \rbzero.spi_registers.texadd1[6] ;
 wire \rbzero.spi_registers.texadd1[7] ;
 wire \rbzero.spi_registers.texadd1[8] ;
 wire \rbzero.spi_registers.texadd1[9] ;
 wire \rbzero.spi_registers.texadd2[0] ;
 wire \rbzero.spi_registers.texadd2[10] ;
 wire \rbzero.spi_registers.texadd2[11] ;
 wire \rbzero.spi_registers.texadd2[12] ;
 wire \rbzero.spi_registers.texadd2[13] ;
 wire \rbzero.spi_registers.texadd2[14] ;
 wire \rbzero.spi_registers.texadd2[15] ;
 wire \rbzero.spi_registers.texadd2[16] ;
 wire \rbzero.spi_registers.texadd2[17] ;
 wire \rbzero.spi_registers.texadd2[18] ;
 wire \rbzero.spi_registers.texadd2[19] ;
 wire \rbzero.spi_registers.texadd2[1] ;
 wire \rbzero.spi_registers.texadd2[20] ;
 wire \rbzero.spi_registers.texadd2[21] ;
 wire \rbzero.spi_registers.texadd2[22] ;
 wire \rbzero.spi_registers.texadd2[23] ;
 wire \rbzero.spi_registers.texadd2[2] ;
 wire \rbzero.spi_registers.texadd2[3] ;
 wire \rbzero.spi_registers.texadd2[4] ;
 wire \rbzero.spi_registers.texadd2[5] ;
 wire \rbzero.spi_registers.texadd2[6] ;
 wire \rbzero.spi_registers.texadd2[7] ;
 wire \rbzero.spi_registers.texadd2[8] ;
 wire \rbzero.spi_registers.texadd2[9] ;
 wire \rbzero.spi_registers.texadd3[0] ;
 wire \rbzero.spi_registers.texadd3[10] ;
 wire \rbzero.spi_registers.texadd3[11] ;
 wire \rbzero.spi_registers.texadd3[12] ;
 wire \rbzero.spi_registers.texadd3[13] ;
 wire \rbzero.spi_registers.texadd3[14] ;
 wire \rbzero.spi_registers.texadd3[15] ;
 wire \rbzero.spi_registers.texadd3[16] ;
 wire \rbzero.spi_registers.texadd3[17] ;
 wire \rbzero.spi_registers.texadd3[18] ;
 wire \rbzero.spi_registers.texadd3[19] ;
 wire \rbzero.spi_registers.texadd3[1] ;
 wire \rbzero.spi_registers.texadd3[20] ;
 wire \rbzero.spi_registers.texadd3[21] ;
 wire \rbzero.spi_registers.texadd3[22] ;
 wire \rbzero.spi_registers.texadd3[23] ;
 wire \rbzero.spi_registers.texadd3[2] ;
 wire \rbzero.spi_registers.texadd3[3] ;
 wire \rbzero.spi_registers.texadd3[4] ;
 wire \rbzero.spi_registers.texadd3[5] ;
 wire \rbzero.spi_registers.texadd3[6] ;
 wire \rbzero.spi_registers.texadd3[7] ;
 wire \rbzero.spi_registers.texadd3[8] ;
 wire \rbzero.spi_registers.texadd3[9] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.texu_hot[0] ;
 wire \rbzero.texu_hot[1] ;
 wire \rbzero.texu_hot[2] ;
 wire \rbzero.texu_hot[3] ;
 wire \rbzero.texu_hot[4] ;
 wire \rbzero.texu_hot[5] ;
 wire \rbzero.trace_state[0] ;
 wire \rbzero.trace_state[1] ;
 wire \rbzero.trace_state[2] ;
 wire \rbzero.trace_state[3] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_hot[0] ;
 wire \rbzero.wall_hot[1] ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \reg_gpout[0] ;
 wire \reg_gpout[1] ;
 wire \reg_gpout[2] ;
 wire \reg_gpout[3] ;
 wire \reg_gpout[4] ;
 wire \reg_gpout[5] ;
 wire reg_hsync;
 wire \reg_rgb[14] ;
 wire \reg_rgb[15] ;
 wire \reg_rgb[22] ;
 wire \reg_rgb[23] ;
 wire \reg_rgb[6] ;
 wire \reg_rgb[7] ;
 wire reg_vsync;
 wire net96;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net130;
 wire net76;
 wire net77;
 wire net128;
 wire net129;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_100_i_clk;
 wire clknet_leaf_101_i_clk;
 wire clknet_leaf_102_i_clk;
 wire clknet_leaf_104_i_clk;
 wire clknet_leaf_105_i_clk;
 wire clknet_leaf_106_i_clk;
 wire clknet_leaf_107_i_clk;
 wire clknet_leaf_108_i_clk;
 wire clknet_leaf_109_i_clk;
 wire clknet_leaf_111_i_clk;
 wire clknet_leaf_112_i_clk;
 wire clknet_leaf_113_i_clk;
 wire clknet_leaf_114_i_clk;
 wire clknet_leaf_116_i_clk;
 wire clknet_leaf_117_i_clk;
 wire clknet_leaf_118_i_clk;
 wire clknet_leaf_119_i_clk;
 wire clknet_leaf_120_i_clk;
 wire clknet_leaf_121_i_clk;
 wire clknet_leaf_122_i_clk;
 wire clknet_leaf_123_i_clk;
 wire clknet_leaf_124_i_clk;
 wire clknet_leaf_125_i_clk;
 wire clknet_leaf_126_i_clk;
 wire clknet_leaf_127_i_clk;
 wire clknet_leaf_128_i_clk;
 wire clknet_leaf_129_i_clk;
 wire clknet_leaf_130_i_clk;
 wire clknet_leaf_131_i_clk;
 wire clknet_leaf_132_i_clk;
 wire clknet_leaf_133_i_clk;
 wire clknet_leaf_134_i_clk;
 wire clknet_leaf_135_i_clk;
 wire clknet_leaf_136_i_clk;
 wire clknet_leaf_137_i_clk;
 wire clknet_leaf_138_i_clk;
 wire clknet_leaf_139_i_clk;
 wire clknet_leaf_140_i_clk;
 wire clknet_leaf_141_i_clk;
 wire clknet_leaf_142_i_clk;
 wire clknet_leaf_143_i_clk;
 wire clknet_leaf_144_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_0_1_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_1_1_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_2_1_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_2_3_1_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_4_0_0_i_clk;
 wire clknet_4_1_0_i_clk;
 wire clknet_4_2_0_i_clk;
 wire clknet_4_3_0_i_clk;
 wire clknet_4_4_0_i_clk;
 wire clknet_4_5_0_i_clk;
 wire clknet_4_6_0_i_clk;
 wire clknet_4_7_0_i_clk;
 wire clknet_4_8_0_i_clk;
 wire clknet_4_9_0_i_clk;
 wire clknet_4_10_0_i_clk;
 wire clknet_4_11_0_i_clk;
 wire clknet_4_12_0_i_clk;
 wire clknet_4_13_0_i_clk;
 wire clknet_4_14_0_i_clk;
 wire clknet_4_15_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_opt_2_0_i_clk;
 wire clknet_opt_3_0_i_clk;
 wire clknet_opt_4_0_i_clk;
 wire clknet_opt_5_0_i_clk;
 wire clknet_opt_6_0_i_clk;
 wire clknet_opt_7_0_i_clk;
 wire clknet_opt_8_0_i_clk;
 wire clknet_0__05731_;
 wire clknet_1_0__leaf__05731_;
 wire clknet_1_1__leaf__05731_;
 wire clknet_0__05991_;
 wire clknet_1_0__leaf__05991_;
 wire clknet_1_1__leaf__05991_;
 wire clknet_0__05762_;
 wire clknet_1_0__leaf__05762_;
 wire clknet_1_1__leaf__05762_;
 wire clknet_0__03849_;
 wire clknet_1_0__leaf__03849_;
 wire clknet_1_1__leaf__03849_;
 wire clknet_0__03848_;
 wire clknet_1_0__leaf__03848_;
 wire clknet_1_1__leaf__03848_;
 wire clknet_0__03837_;
 wire clknet_1_0__leaf__03837_;
 wire clknet_1_1__leaf__03837_;
 wire clknet_0__03847_;
 wire clknet_1_0__leaf__03847_;
 wire clknet_1_1__leaf__03847_;
 wire clknet_0__03846_;
 wire clknet_1_0__leaf__03846_;
 wire clknet_1_1__leaf__03846_;
 wire clknet_0__03845_;
 wire clknet_1_0__leaf__03845_;
 wire clknet_1_1__leaf__03845_;
 wire clknet_0__03844_;
 wire clknet_1_0__leaf__03844_;
 wire clknet_1_1__leaf__03844_;
 wire clknet_0__03843_;
 wire clknet_1_0__leaf__03843_;
 wire clknet_1_1__leaf__03843_;
 wire clknet_0__03842_;
 wire clknet_1_0__leaf__03842_;
 wire clknet_1_1__leaf__03842_;
 wire clknet_0__03841_;
 wire clknet_1_0__leaf__03841_;
 wire clknet_1_1__leaf__03841_;
 wire clknet_0__03840_;
 wire clknet_1_0__leaf__03840_;
 wire clknet_1_1__leaf__03840_;
 wire clknet_0__03839_;
 wire clknet_1_0__leaf__03839_;
 wire clknet_1_1__leaf__03839_;
 wire clknet_0__03838_;
 wire clknet_1_0__leaf__03838_;
 wire clknet_1_1__leaf__03838_;
 wire clknet_0__03826_;
 wire clknet_1_0__leaf__03826_;
 wire clknet_1_1__leaf__03826_;
 wire clknet_0__03836_;
 wire clknet_1_0__leaf__03836_;
 wire clknet_1_1__leaf__03836_;
 wire clknet_0__03835_;
 wire clknet_1_0__leaf__03835_;
 wire clknet_1_1__leaf__03835_;
 wire clknet_0__03834_;
 wire clknet_1_0__leaf__03834_;
 wire clknet_1_1__leaf__03834_;
 wire clknet_0__03833_;
 wire clknet_1_0__leaf__03833_;
 wire clknet_1_1__leaf__03833_;
 wire clknet_0__03832_;
 wire clknet_1_0__leaf__03832_;
 wire clknet_1_1__leaf__03832_;
 wire clknet_0__03831_;
 wire clknet_1_0__leaf__03831_;
 wire clknet_1_1__leaf__03831_;
 wire clknet_0__03830_;
 wire clknet_1_0__leaf__03830_;
 wire clknet_1_1__leaf__03830_;
 wire clknet_0__03829_;
 wire clknet_1_0__leaf__03829_;
 wire clknet_1_1__leaf__03829_;
 wire clknet_0__03828_;
 wire clknet_1_0__leaf__03828_;
 wire clknet_1_1__leaf__03828_;
 wire clknet_0__03827_;
 wire clknet_1_0__leaf__03827_;
 wire clknet_1_1__leaf__03827_;
 wire clknet_0__03616_;
 wire clknet_1_0__leaf__03616_;
 wire clknet_1_1__leaf__03616_;
 wire clknet_0__03825_;
 wire clknet_1_0__leaf__03825_;
 wire clknet_1_1__leaf__03825_;
 wire clknet_0__03824_;
 wire clknet_1_0__leaf__03824_;
 wire clknet_1_1__leaf__03824_;
 wire clknet_0__03823_;
 wire clknet_1_0__leaf__03823_;
 wire clknet_1_1__leaf__03823_;
 wire clknet_0__03822_;
 wire clknet_1_0__leaf__03822_;
 wire clknet_1_1__leaf__03822_;
 wire clknet_0__03821_;
 wire clknet_1_0__leaf__03821_;
 wire clknet_1_1__leaf__03821_;
 wire clknet_0__03820_;
 wire clknet_1_0__leaf__03820_;
 wire clknet_1_1__leaf__03820_;
 wire clknet_0__03819_;
 wire clknet_1_0__leaf__03819_;
 wire clknet_1_1__leaf__03819_;
 wire clknet_0__03818_;
 wire clknet_1_0__leaf__03818_;
 wire clknet_1_1__leaf__03818_;
 wire clknet_0__03817_;
 wire clknet_1_0__leaf__03817_;
 wire clknet_1_1__leaf__03817_;
 wire clknet_0__03617_;
 wire clknet_1_0__leaf__03617_;
 wire clknet_1_1__leaf__03617_;
 wire clknet_0__03609_;
 wire clknet_1_0__leaf__03609_;
 wire clknet_1_1__leaf__03609_;
 wire clknet_0__03615_;
 wire clknet_1_0__leaf__03615_;
 wire clknet_1_1__leaf__03615_;
 wire clknet_0__03614_;
 wire clknet_1_0__leaf__03614_;
 wire clknet_1_1__leaf__03614_;
 wire clknet_0__03613_;
 wire clknet_1_0__leaf__03613_;
 wire clknet_1_1__leaf__03613_;
 wire clknet_0__03612_;
 wire clknet_1_0__leaf__03612_;
 wire clknet_1_1__leaf__03612_;
 wire clknet_0__03611_;
 wire clknet_1_0__leaf__03611_;
 wire clknet_1_1__leaf__03611_;
 wire clknet_0__03610_;
 wire clknet_1_0__leaf__03610_;
 wire clknet_1_1__leaf__03610_;
 wire clknet_0__05944_;
 wire clknet_1_0__leaf__05944_;
 wire clknet_1_1__leaf__05944_;
 wire clknet_0__05893_;
 wire clknet_1_0__leaf__05893_;
 wire clknet_1_1__leaf__05893_;
 wire clknet_0__05839_;
 wire clknet_1_0__leaf__05839_;
 wire clknet_1_1__leaf__05839_;
 wire clknet_0__05786_;
 wire clknet_1_0__leaf__05786_;
 wire clknet_1_1__leaf__05786_;
 wire net75;
 wire net514;
 wire net515;
 wire net516;

 sky130_fd_sc_hd__buf_4 _10449_ (.A(\gpout0.hpos[0] ),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_4 _10450_ (.A(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__buf_4 _10451_ (.A(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__buf_4 _10452_ (.A(\gpout0.hpos[7] ),
    .X(_04013_));
 sky130_fd_sc_hd__clkbuf_4 _10453_ (.A(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__xor2_4 _10454_ (.A(net47),
    .B(net48),
    .X(_04015_));
 sky130_fd_sc_hd__buf_4 _10455_ (.A(\gpout0.hpos[8] ),
    .X(_04016_));
 sky130_fd_sc_hd__clkbuf_4 _10456_ (.A(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__clkbuf_4 _10457_ (.A(\gpout0.hpos[9] ),
    .X(_04018_));
 sky130_fd_sc_hd__and2b_1 _10458_ (.A_N(_04017_),
    .B(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__and4_4 _10459_ (.A(_04012_),
    .B(_04014_),
    .C(_04015_),
    .D(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__buf_4 _10460_ (.A(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_4 _10461_ (.A(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(\rbzero.tex_r1[63] ),
    .A1(net51),
    .S(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__clkbuf_1 _10463_ (.A(_04023_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[63] ),
    .S(_04022_),
    .X(_04024_));
 sky130_fd_sc_hd__clkbuf_1 _10465_ (.A(_04024_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _10466_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_04022_),
    .X(_04025_));
 sky130_fd_sc_hd__clkbuf_1 _10467_ (.A(_04025_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(_04022_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_1 _10469_ (.A(_04026_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_04022_),
    .X(_04027_));
 sky130_fd_sc_hd__clkbuf_1 _10471_ (.A(_04027_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_04022_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_1 _10473_ (.A(_04028_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _10474_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_04022_),
    .X(_04029_));
 sky130_fd_sc_hd__clkbuf_1 _10475_ (.A(_04029_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(_04022_),
    .X(_04030_));
 sky130_fd_sc_hd__clkbuf_1 _10477_ (.A(_04030_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _10478_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_04022_),
    .X(_04031_));
 sky130_fd_sc_hd__clkbuf_1 _10479_ (.A(_04031_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(_04022_),
    .X(_04032_));
 sky130_fd_sc_hd__clkbuf_1 _10481_ (.A(_04032_),
    .X(_01577_));
 sky130_fd_sc_hd__clkbuf_4 _10482_ (.A(_04021_),
    .X(_04033_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__clkbuf_1 _10484_ (.A(_04034_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(_04033_),
    .X(_04035_));
 sky130_fd_sc_hd__clkbuf_1 _10486_ (.A(_04035_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_04033_),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_1 _10488_ (.A(_04036_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_04033_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _10490_ (.A(_04037_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_04033_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _10492_ (.A(_04038_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(_04033_),
    .X(_04039_));
 sky130_fd_sc_hd__clkbuf_1 _10494_ (.A(_04039_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_04033_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_1 _10496_ (.A(_04040_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(_04033_),
    .X(_04041_));
 sky130_fd_sc_hd__clkbuf_1 _10498_ (.A(_04041_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _10499_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_04033_),
    .X(_04042_));
 sky130_fd_sc_hd__clkbuf_1 _10500_ (.A(_04042_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(_04033_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(_04043_),
    .X(_01567_));
 sky130_fd_sc_hd__clkbuf_4 _10503_ (.A(_04021_),
    .X(_04044_));
 sky130_fd_sc_hd__mux2_1 _10504_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _10505_ (.A(_04045_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(_04044_),
    .X(_04046_));
 sky130_fd_sc_hd__clkbuf_1 _10507_ (.A(_04046_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_04044_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_1 _10509_ (.A(_04047_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(_04044_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_1 _10511_ (.A(_04048_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _10512_ (.A0(\rbzero.tex_r1[39] ),
    .A1(net75),
    .S(_04044_),
    .X(_04049_));
 sky130_fd_sc_hd__clkbuf_1 _10513_ (.A(_04049_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(_04044_),
    .X(_04050_));
 sky130_fd_sc_hd__clkbuf_1 _10515_ (.A(_04050_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04044_),
    .X(_04051_));
 sky130_fd_sc_hd__clkbuf_1 _10517_ (.A(_04051_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_04044_),
    .X(_04052_));
 sky130_fd_sc_hd__clkbuf_1 _10519_ (.A(_04052_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _10520_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_04044_),
    .X(_04053_));
 sky130_fd_sc_hd__clkbuf_1 _10521_ (.A(_04053_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(_04044_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_1 _10523_ (.A(_04054_),
    .X(_01557_));
 sky130_fd_sc_hd__clkbuf_4 _10524_ (.A(_04021_),
    .X(_04055_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_1 _10526_ (.A(_04056_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _10527_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(_04055_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_1 _10528_ (.A(_04057_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_04055_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _10530_ (.A(_04058_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(_04055_),
    .X(_04059_));
 sky130_fd_sc_hd__clkbuf_1 _10532_ (.A(_04059_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _10533_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_04055_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _10534_ (.A(_04060_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(_04055_),
    .X(_04061_));
 sky130_fd_sc_hd__clkbuf_1 _10536_ (.A(_04061_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_04055_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_1 _10538_ (.A(_04062_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(_04055_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _10540_ (.A(_04063_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_04055_),
    .X(_04064_));
 sky130_fd_sc_hd__clkbuf_1 _10542_ (.A(_04064_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(_04055_),
    .X(_04065_));
 sky130_fd_sc_hd__clkbuf_1 _10544_ (.A(_04065_),
    .X(_01547_));
 sky130_fd_sc_hd__clkbuf_4 _10545_ (.A(_04021_),
    .X(_04066_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_04067_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(_04066_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_1 _10549_ (.A(_04068_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_04066_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _10551_ (.A(_04069_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(_04066_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_1 _10553_ (.A(_04070_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _10554_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_04066_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _10555_ (.A(_04071_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10556_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(_04066_),
    .X(_04072_));
 sky130_fd_sc_hd__clkbuf_1 _10557_ (.A(_04072_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_04066_),
    .X(_04073_));
 sky130_fd_sc_hd__clkbuf_1 _10559_ (.A(_04073_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(_04066_),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _10561_ (.A(_04074_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_04066_),
    .X(_04075_));
 sky130_fd_sc_hd__clkbuf_1 _10563_ (.A(_04075_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(_04066_),
    .X(_04076_));
 sky130_fd_sc_hd__clkbuf_1 _10565_ (.A(_04076_),
    .X(_01537_));
 sky130_fd_sc_hd__clkbuf_4 _10566_ (.A(_04021_),
    .X(_04077_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__clkbuf_1 _10568_ (.A(_04078_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_04077_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _10570_ (.A(_04079_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10571_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_04077_),
    .X(_04080_));
 sky130_fd_sc_hd__clkbuf_1 _10572_ (.A(_04080_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(_04077_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_1 _10574_ (.A(_04081_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_04077_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _10576_ (.A(_04082_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10577_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_04077_),
    .X(_04083_));
 sky130_fd_sc_hd__clkbuf_1 _10578_ (.A(_04083_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04077_),
    .X(_04084_));
 sky130_fd_sc_hd__clkbuf_1 _10580_ (.A(_04084_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(_04077_),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _10582_ (.A(_04085_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04077_),
    .X(_04086_));
 sky130_fd_sc_hd__clkbuf_1 _10584_ (.A(_04086_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(_04077_),
    .X(_04087_));
 sky130_fd_sc_hd__clkbuf_1 _10586_ (.A(_04087_),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_4 _10587_ (.A(_04021_),
    .X(_04088_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_1 _10589_ (.A(_04089_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_04088_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_1 _10591_ (.A(_04090_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10592_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_04088_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _10593_ (.A(_04091_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\rbzero.tex_r1[0] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(_04088_),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _10595_ (.A(_04092_),
    .X(_01523_));
 sky130_fd_sc_hd__inv_2 _10596_ (.A(_04013_),
    .Y(_04093_));
 sky130_fd_sc_hd__inv_6 _10597_ (.A(_04015_),
    .Y(_04094_));
 sky130_fd_sc_hd__or4b_4 _10598_ (.A(_04011_),
    .B(_04093_),
    .C(_04094_),
    .D_N(_04019_),
    .X(_04095_));
 sky130_fd_sc_hd__buf_4 _10599_ (.A(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_4 _10600_ (.A(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(net51),
    .A1(\rbzero.tex_r0[63] ),
    .S(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_04098_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04097_),
    .X(_04099_));
 sky130_fd_sc_hd__clkbuf_1 _10604_ (.A(_04099_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_04097_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_04100_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04097_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(_04101_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(_04097_),
    .X(_04102_));
 sky130_fd_sc_hd__clkbuf_1 _10610_ (.A(_04102_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04097_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _10612_ (.A(_04103_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(_04097_),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_04104_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04097_),
    .X(_04105_));
 sky130_fd_sc_hd__clkbuf_1 _10616_ (.A(_04105_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10617_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(_04097_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _10618_ (.A(_04106_),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _10619_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04097_),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _10620_ (.A(_04107_),
    .X(_01513_));
 sky130_fd_sc_hd__clkbuf_4 _10621_ (.A(_04096_),
    .X(_04108_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_04109_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04108_),
    .X(_04110_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_04110_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_04108_),
    .X(_04111_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(_04111_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_04108_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_04112_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(_04108_),
    .X(_04113_));
 sky130_fd_sc_hd__clkbuf_1 _10631_ (.A(_04113_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04108_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_04114_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(_04108_),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _10635_ (.A(_04115_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04108_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _10637_ (.A(_04116_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_04108_),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_04117_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04108_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _10641_ (.A(_04118_),
    .X(_01503_));
 sky130_fd_sc_hd__clkbuf_4 _10642_ (.A(_04096_),
    .X(_04119_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(_04120_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04119_),
    .X(_04121_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(_04121_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(_04119_),
    .X(_04122_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(_04122_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04119_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(_04123_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(_04119_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _10652_ (.A(_04124_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04119_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _10654_ (.A(_04125_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(_04119_),
    .X(_04126_));
 sky130_fd_sc_hd__clkbuf_1 _10656_ (.A(_04126_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04119_),
    .X(_04127_));
 sky130_fd_sc_hd__clkbuf_1 _10658_ (.A(_04127_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(_04119_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _10660_ (.A(_04128_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04119_),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_1 _10662_ (.A(_04129_),
    .X(_01493_));
 sky130_fd_sc_hd__clkbuf_4 _10663_ (.A(_04096_),
    .X(_04130_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(_04131_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04130_),
    .X(_04132_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(_04132_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(_04130_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(_04133_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04130_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(_04134_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(_04130_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_1 _10673_ (.A(_04135_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04130_),
    .X(_04136_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_04136_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_04130_),
    .X(_04137_));
 sky130_fd_sc_hd__clkbuf_1 _10677_ (.A(_04137_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04130_),
    .X(_04138_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_04138_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(_04130_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_04139_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04130_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_1 _10683_ (.A(_04140_),
    .X(_01483_));
 sky130_fd_sc_hd__clkbuf_4 _10684_ (.A(_04096_),
    .X(_04141_));
 sky130_fd_sc_hd__mux2_1 _10685_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(_04141_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _10686_ (.A(_04142_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04141_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _10688_ (.A(_04143_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(_04141_),
    .X(_04144_));
 sky130_fd_sc_hd__clkbuf_1 _10690_ (.A(_04144_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04141_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _10692_ (.A(_04145_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _10693_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(_04141_),
    .X(_04146_));
 sky130_fd_sc_hd__clkbuf_1 _10694_ (.A(_04146_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04141_),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _10696_ (.A(_04147_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(_04141_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_1 _10698_ (.A(_04148_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04141_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_1 _10700_ (.A(_04149_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(_04141_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _10702_ (.A(_04150_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04141_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _10704_ (.A(_04151_),
    .X(_01473_));
 sky130_fd_sc_hd__clkbuf_4 _10705_ (.A(_04096_),
    .X(_04152_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(_04153_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04152_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(_04154_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(_04152_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(_04155_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04152_),
    .X(_04156_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(_04156_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_04152_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _10715_ (.A(_04157_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04152_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _10717_ (.A(_04158_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(_04152_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _10719_ (.A(_04159_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04152_),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_04160_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(_04152_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _10723_ (.A(_04161_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04152_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10725_ (.A(_04162_),
    .X(_01463_));
 sky130_fd_sc_hd__buf_4 _10726_ (.A(_04096_),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(_04164_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _10729_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_04163_),
    .X(_04165_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(_04165_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10731_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_04163_),
    .X(_04166_));
 sky130_fd_sc_hd__clkbuf_1 _10732_ (.A(_04166_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04163_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _10734_ (.A(_04167_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10735_ (.A0(\rbzero.tex_g1[63] ),
    .A1(net52),
    .S(_04088_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _10736_ (.A(_04168_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[63] ),
    .S(_04088_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _10738_ (.A(_04169_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10739_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_04088_),
    .X(_04170_));
 sky130_fd_sc_hd__clkbuf_1 _10740_ (.A(_04170_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(_04088_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _10742_ (.A(_04171_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04088_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _10744_ (.A(_04172_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_04088_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _10746_ (.A(_04173_),
    .X(_01453_));
 sky130_fd_sc_hd__clkbuf_4 _10747_ (.A(_04021_),
    .X(_04174_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _10749_ (.A(_04175_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(_04174_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _10751_ (.A(_04176_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_04174_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(_04177_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(_04174_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _10755_ (.A(_04178_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_04174_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _10757_ (.A(_04179_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(_04174_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_04180_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04174_),
    .X(_04181_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_04181_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(_04174_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_04182_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04174_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_04183_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_04174_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(_04184_),
    .X(_01443_));
 sky130_fd_sc_hd__buf_4 _10768_ (.A(_04020_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_4 _10769_ (.A(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _10771_ (.A(_04187_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(_04186_),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _10773_ (.A(_04188_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_04186_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _10775_ (.A(_04189_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(_04186_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _10777_ (.A(_04190_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10778_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_04186_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _10779_ (.A(_04191_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10780_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(_04186_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _10781_ (.A(_04192_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10782_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_04186_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _10783_ (.A(_04193_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10784_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_04186_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _10785_ (.A(_04194_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10786_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_04186_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _10787_ (.A(_04195_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _10788_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(_04186_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _10789_ (.A(_04196_),
    .X(_01433_));
 sky130_fd_sc_hd__clkbuf_4 _10790_ (.A(_04185_),
    .X(_04197_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_04198_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(_04197_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _10794_ (.A(_04199_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_04197_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_04200_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(_04197_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _10798_ (.A(_04201_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_04197_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _10800_ (.A(_04202_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10801_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(_04197_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _10802_ (.A(_04203_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_04197_),
    .X(_04204_));
 sky130_fd_sc_hd__clkbuf_1 _10804_ (.A(_04204_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10805_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(_04197_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _10806_ (.A(_04205_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_04197_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _10808_ (.A(_04206_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _10809_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(_04197_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _10810_ (.A(_04207_),
    .X(_01423_));
 sky130_fd_sc_hd__clkbuf_4 _10811_ (.A(_04185_),
    .X(_04208_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(_04209_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(_04208_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _10815_ (.A(_04210_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_04208_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_04211_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(_04208_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _10819_ (.A(_04212_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _10820_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04208_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _10821_ (.A(_04213_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10822_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(_04208_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _10823_ (.A(_04214_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_04208_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _10825_ (.A(_04215_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10826_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(_04208_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _10827_ (.A(_04216_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04208_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _10829_ (.A(_04217_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _10830_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(_04208_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _10831_ (.A(_04218_),
    .X(_01413_));
 sky130_fd_sc_hd__clkbuf_4 _10832_ (.A(_04185_),
    .X(_04219_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_04220_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(_04219_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(_04221_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_04219_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(_04222_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(_04219_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(_04223_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10841_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_04219_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _10842_ (.A(_04224_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(_04219_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _10844_ (.A(_04225_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_04219_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _10846_ (.A(_04226_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(_04219_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _10848_ (.A(_04227_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_04219_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_04228_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(_04219_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _10852_ (.A(_04229_),
    .X(_01403_));
 sky130_fd_sc_hd__buf_4 _10853_ (.A(_04185_),
    .X(_04230_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _10855_ (.A(_04231_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _10856_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(_04230_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _10857_ (.A(_04232_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _10858_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_04230_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _10859_ (.A(_04233_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _10860_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(_04230_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _10861_ (.A(_04234_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_04230_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _10863_ (.A(_04235_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(_04230_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _10865_ (.A(_04236_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_04230_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(_04237_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(\rbzero.tex_g1[0] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_04230_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(_04238_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(net52),
    .A1(\rbzero.tex_g0[63] ),
    .S(_04163_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _10871_ (.A(_04239_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_04163_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_04240_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(_04163_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(_04241_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04163_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(_04242_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_04163_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_04243_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04163_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(_04244_),
    .X(_01389_));
 sky130_fd_sc_hd__clkbuf_4 _10882_ (.A(_04096_),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _10884_ (.A(_04246_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_04245_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(_04247_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(_04245_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_04248_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04245_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_04249_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(_04245_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_04250_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_04245_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_04251_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(_04245_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(_04252_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_04245_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_04253_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(_04245_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_04254_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04245_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_04255_),
    .X(_01379_));
 sky130_fd_sc_hd__buf_4 _10903_ (.A(_04095_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_4 _10904_ (.A(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(_04258_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04257_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_04259_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(_04257_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_04260_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_04257_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_04261_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(_04257_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(_04262_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _10915_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04257_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _10916_ (.A(_04263_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _10917_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_04257_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _10918_ (.A(_04264_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _10919_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04257_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _10920_ (.A(_04265_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(_04257_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _10922_ (.A(_04266_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _10923_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04257_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _10924_ (.A(_04267_),
    .X(_01369_));
 sky130_fd_sc_hd__clkbuf_4 _10925_ (.A(_04256_),
    .X(_04268_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(_04269_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04268_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_04270_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(_04268_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _10931_ (.A(_04271_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04268_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _10933_ (.A(_04272_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _10934_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(_04268_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _10935_ (.A(_04273_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04268_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_1 _10937_ (.A(_04274_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(_04268_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _10939_ (.A(_04275_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _10940_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_04268_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _10941_ (.A(_04276_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _10942_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(_04268_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _10943_ (.A(_04277_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _10944_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04268_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _10945_ (.A(_04278_),
    .X(_01359_));
 sky130_fd_sc_hd__clkbuf_4 _10946_ (.A(_04256_),
    .X(_04279_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_04280_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_04279_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_04281_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(_04279_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _10952_ (.A(_04282_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _10953_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_04279_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _10954_ (.A(_04283_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(_04279_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _10956_ (.A(_04284_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04279_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _10958_ (.A(_04285_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _10959_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(_04279_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _10960_ (.A(_04286_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04279_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _10962_ (.A(_04287_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10963_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(_04279_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _10964_ (.A(_04288_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_04279_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _10966_ (.A(_04289_),
    .X(_01349_));
 sky130_fd_sc_hd__clkbuf_4 _10967_ (.A(_04256_),
    .X(_04290_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_04291_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04290_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(_04292_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(_04290_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(_04293_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_04290_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _10975_ (.A(_04294_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10976_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(_04290_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _10977_ (.A(_04295_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _10978_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04290_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _10979_ (.A(_04296_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _10980_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_04290_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _10981_ (.A(_04297_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_04290_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _10983_ (.A(_04298_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(_04290_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(_04299_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04290_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _10987_ (.A(_04300_),
    .X(_01339_));
 sky130_fd_sc_hd__buf_4 _10988_ (.A(_04256_),
    .X(_04301_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _10990_ (.A(_04302_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04301_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _10992_ (.A(_04303_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(_04301_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _10994_ (.A(_04304_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04301_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _10996_ (.A(_04305_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(_04301_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _10998_ (.A(_04306_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_04301_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _11000_ (.A(_04307_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_04301_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _11002_ (.A(_04308_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_04301_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(_04309_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\rbzero.tex_b1[63] ),
    .A1(net53),
    .S(_04230_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_04310_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[63] ),
    .S(_04230_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _11008_ (.A(_04311_),
    .X(_01329_));
 sky130_fd_sc_hd__clkbuf_4 _11009_ (.A(_04185_),
    .X(_04312_));
 sky130_fd_sc_hd__mux2_1 _11010_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _11011_ (.A(_04313_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(_04312_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _11013_ (.A(_04314_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04312_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _11015_ (.A(_04315_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(_04312_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _11017_ (.A(_04316_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_04312_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _11019_ (.A(_04317_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(_04312_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _11021_ (.A(_04318_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_04312_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _11023_ (.A(_04319_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(_04312_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _11025_ (.A(_04320_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04312_),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_1 _11027_ (.A(_04321_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(_04312_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _11029_ (.A(_04322_),
    .X(_01319_));
 sky130_fd_sc_hd__clkbuf_4 _11030_ (.A(_04185_),
    .X(_04323_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _11032_ (.A(_04324_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(_04323_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _11034_ (.A(_04325_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04323_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _11036_ (.A(_04326_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(_04323_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _11038_ (.A(_04327_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04323_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _11040_ (.A(_04328_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(_04323_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _11042_ (.A(_04329_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04323_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _11044_ (.A(_04330_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(_04323_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _11046_ (.A(_04331_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_04323_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_04332_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(_04323_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _11050_ (.A(_04333_),
    .X(_01309_));
 sky130_fd_sc_hd__clkbuf_4 _11051_ (.A(_04185_),
    .X(_04334_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _11053_ (.A(_04335_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(_04334_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(_04336_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_04334_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _11057_ (.A(_04337_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(_04334_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _11059_ (.A(_04338_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04334_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(_04339_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(_04334_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(_04340_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_04334_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(_04341_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(_04334_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(_04342_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_04334_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(_04343_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(_04334_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _11071_ (.A(_04344_),
    .X(_01299_));
 sky130_fd_sc_hd__clkbuf_4 _11072_ (.A(_04185_),
    .X(_04345_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _11074_ (.A(_04346_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(_04345_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _11076_ (.A(_04347_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_04345_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _11078_ (.A(_04348_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_04345_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _11080_ (.A(_04349_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_04345_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _11082_ (.A(_04350_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(_04345_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _11084_ (.A(_04351_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_04345_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _11086_ (.A(_04352_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(_04345_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _11088_ (.A(_04353_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_04345_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _11090_ (.A(_04354_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _11091_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_04345_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _11092_ (.A(_04355_),
    .X(_01289_));
 sky130_fd_sc_hd__clkbuf_4 _11093_ (.A(_04185_),
    .X(_04356_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(_04357_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(_04356_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(_04358_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04356_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(_04359_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(_04356_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(_04360_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_04356_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _11103_ (.A(_04361_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(_04356_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _11105_ (.A(_04362_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04356_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _11107_ (.A(_04363_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_04356_),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _11109_ (.A(_04364_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04356_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _11111_ (.A(_04365_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(_04356_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _11113_ (.A(_04366_),
    .X(_01279_));
 sky130_fd_sc_hd__clkbuf_4 _11114_ (.A(_04020_),
    .X(_04367_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(_04368_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(_04367_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(_04369_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04367_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_1 _11120_ (.A(_04370_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_04367_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _11122_ (.A(_04371_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _11123_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04367_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _11124_ (.A(_04372_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(_04367_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _11126_ (.A(_04373_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04367_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _11128_ (.A(_04374_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_04367_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(_04375_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _11131_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04367_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _11132_ (.A(_04376_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _11133_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_04367_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _11134_ (.A(_04377_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _11135_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_04021_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _11136_ (.A(_04378_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _11137_ (.A0(\rbzero.tex_b1[0] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_04021_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _11138_ (.A(_04379_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _11139_ (.A0(net53),
    .A1(\rbzero.tex_b0[63] ),
    .S(_04301_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _11140_ (.A(_04380_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _11141_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_04301_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _11142_ (.A(_04381_),
    .X(_01172_));
 sky130_fd_sc_hd__clkbuf_4 _11143_ (.A(_04256_),
    .X(_04382_));
 sky130_fd_sc_hd__mux2_1 _11144_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_04382_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _11145_ (.A(_04383_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_04382_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _11147_ (.A(_04384_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(_04382_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _11149_ (.A(_04385_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_04382_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _11151_ (.A(_04386_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(_04382_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _11153_ (.A(_04387_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_04382_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(_04388_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(_04382_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _11157_ (.A(_04389_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _11158_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_04382_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _11159_ (.A(_04390_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(_04382_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _11161_ (.A(_04391_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_04382_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _11163_ (.A(_04392_),
    .X(_01162_));
 sky130_fd_sc_hd__clkbuf_4 _11164_ (.A(_04256_),
    .X(_04393_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _11166_ (.A(_04394_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04393_),
    .X(_04395_));
 sky130_fd_sc_hd__clkbuf_1 _11168_ (.A(_04395_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(_04393_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(_04396_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_04393_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(_04397_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(_04393_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _11174_ (.A(_04398_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_04393_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _11176_ (.A(_04399_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _11177_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_04393_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _11178_ (.A(_04400_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _11179_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_04393_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _11180_ (.A(_04401_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _11181_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_04393_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _11182_ (.A(_04402_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_04393_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _11184_ (.A(_04403_),
    .X(_01152_));
 sky130_fd_sc_hd__clkbuf_4 _11185_ (.A(_04256_),
    .X(_04404_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _11187_ (.A(_04405_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_04404_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(_04406_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(_04404_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _11191_ (.A(_04407_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_04404_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_1 _11193_ (.A(_04408_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(_04404_),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_1 _11195_ (.A(_04409_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _11196_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04404_),
    .X(_04410_));
 sky130_fd_sc_hd__clkbuf_1 _11197_ (.A(_04410_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_04404_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _11199_ (.A(_04411_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_04404_),
    .X(_04412_));
 sky130_fd_sc_hd__clkbuf_1 _11201_ (.A(_04412_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _11202_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(_04404_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _11203_ (.A(_04413_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _11204_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_04404_),
    .X(_04414_));
 sky130_fd_sc_hd__clkbuf_1 _11205_ (.A(_04414_),
    .X(_01142_));
 sky130_fd_sc_hd__clkbuf_4 _11206_ (.A(_04256_),
    .X(_04415_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(_04416_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_04415_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(_04417_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(_04415_),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_1 _11212_ (.A(_04418_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_04415_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _11214_ (.A(_04419_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _11215_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(_04415_),
    .X(_04420_));
 sky130_fd_sc_hd__clkbuf_1 _11216_ (.A(_04420_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_04415_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_1 _11218_ (.A(_04421_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(_04415_),
    .X(_04422_));
 sky130_fd_sc_hd__clkbuf_1 _11220_ (.A(_04422_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _11221_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04415_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _11222_ (.A(_04423_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _11223_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(_04415_),
    .X(_04424_));
 sky130_fd_sc_hd__clkbuf_1 _11224_ (.A(_04424_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _11225_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_04415_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _11226_ (.A(_04425_),
    .X(_01132_));
 sky130_fd_sc_hd__clkbuf_4 _11227_ (.A(_04256_),
    .X(_04426_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _11229_ (.A(_04427_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _11230_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04426_),
    .X(_04428_));
 sky130_fd_sc_hd__clkbuf_1 _11231_ (.A(_04428_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(_04426_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _11233_ (.A(_04429_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_04426_),
    .X(_04430_));
 sky130_fd_sc_hd__clkbuf_1 _11235_ (.A(_04430_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(_04426_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _11237_ (.A(_04431_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04426_),
    .X(_04432_));
 sky130_fd_sc_hd__clkbuf_1 _11239_ (.A(_04432_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(_04426_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _11241_ (.A(_04433_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _11242_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_04426_),
    .X(_04434_));
 sky130_fd_sc_hd__clkbuf_1 _11243_ (.A(_04434_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_04426_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _11245_ (.A(_04435_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _11246_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_04426_),
    .X(_04436_));
 sky130_fd_sc_hd__clkbuf_1 _11247_ (.A(_04436_),
    .X(_01122_));
 sky130_fd_sc_hd__clkbuf_4 _11248_ (.A(_04095_),
    .X(_04437_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__clkbuf_1 _11250_ (.A(_04438_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_04437_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _11252_ (.A(_04439_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _11253_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(_04437_),
    .X(_04440_));
 sky130_fd_sc_hd__clkbuf_1 _11254_ (.A(_04440_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_04437_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _11256_ (.A(_04441_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _11257_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(_04437_),
    .X(_04442_));
 sky130_fd_sc_hd__clkbuf_1 _11258_ (.A(_04442_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_04437_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _11260_ (.A(_04443_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _11261_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(_04437_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_1 _11262_ (.A(_04444_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _11263_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04437_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _11264_ (.A(_04445_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _11265_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(_04437_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _11266_ (.A(_04446_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _11267_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_04437_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _11268_ (.A(_04447_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _11269_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_04096_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _11270_ (.A(_04448_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _11271_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04096_),
    .X(_04449_));
 sky130_fd_sc_hd__clkbuf_1 _11272_ (.A(_04449_),
    .X(_01110_));
 sky130_fd_sc_hd__buf_6 _11273_ (.A(_04094_),
    .X(_04450_));
 sky130_fd_sc_hd__buf_8 _11274_ (.A(_04450_),
    .X(net65));
 sky130_fd_sc_hd__buf_4 _11275_ (.A(\gpout0.hpos[5] ),
    .X(_04451_));
 sky130_fd_sc_hd__buf_4 _11276_ (.A(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__buf_4 _11277_ (.A(\gpout0.hpos[3] ),
    .X(_04453_));
 sky130_fd_sc_hd__inv_2 _11278_ (.A(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__clkinv_4 _11279_ (.A(\gpout0.hpos[4] ),
    .Y(_04455_));
 sky130_fd_sc_hd__nor2_2 _11280_ (.A(_04454_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__buf_4 _11281_ (.A(\gpout0.hpos[6] ),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_4 _11282_ (.A(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__o21ai_1 _11283_ (.A1(_04452_),
    .A2(_04456_),
    .B1(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__and3_1 _11284_ (.A(\gpout0.hpos[3] ),
    .B(\gpout0.hpos[5] ),
    .C(\gpout0.hpos[4] ),
    .X(_04460_));
 sky130_fd_sc_hd__or3b_1 _11285_ (.A(_04014_),
    .B(_04017_),
    .C_N(_04018_),
    .X(_04461_));
 sky130_fd_sc_hd__or3_1 _11286_ (.A(_04459_),
    .B(_04460_),
    .C(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__buf_4 _11287_ (.A(_04462_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 _11288_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_04463_));
 sky130_fd_sc_hd__buf_2 _11289_ (.A(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__or2_2 _11290_ (.A(\rbzero.trace_state[1] ),
    .B(\rbzero.trace_state[0] ),
    .X(_04465_));
 sky130_fd_sc_hd__clkinv_2 _11291_ (.A(\rbzero.vga_sync.vsync ),
    .Y(_04466_));
 sky130_fd_sc_hd__nand2_1 _11292_ (.A(_04466_),
    .B(_04015_),
    .Y(_04467_));
 sky130_fd_sc_hd__inv_2 _11293_ (.A(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__buf_4 _11294_ (.A(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__o31a_1 _11295_ (.A1(\rbzero.trace_state[3] ),
    .A2(\rbzero.trace_state[2] ),
    .A3(_04465_),
    .B1(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__buf_2 _11296_ (.A(\rbzero.trace_state[0] ),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_4 _11297_ (.A(\rbzero.trace_state[1] ),
    .X(_04472_));
 sky130_fd_sc_hd__nand2b_2 _11298_ (.A_N(\rbzero.trace_state[2] ),
    .B(\rbzero.trace_state[3] ),
    .Y(_04473_));
 sky130_fd_sc_hd__nor2_1 _11299_ (.A(_04472_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__nor2_1 _11300_ (.A(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .Y(_04475_));
 sky130_fd_sc_hd__and3_1 _11301_ (.A(_04472_),
    .B(_04471_),
    .C(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__a21oi_1 _11302_ (.A1(_04471_),
    .A2(_04474_),
    .B1(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__buf_4 _11303_ (.A(_04469_),
    .X(_04478_));
 sky130_fd_sc_hd__a32o_1 _11304_ (.A1(_04464_),
    .A2(_04470_),
    .A3(_04477_),
    .B1(_04476_),
    .B2(_04478_),
    .X(_00001_));
 sky130_fd_sc_hd__a21bo_2 _11305_ (.A1(_04093_),
    .A2(_04459_),
    .B1_N(_04019_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 _11306_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_4 _11307_ (.A(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__a21bo_1 _11308_ (.A1(_04480_),
    .A2(_04477_),
    .B1_N(_04470_),
    .X(_00000_));
 sky130_fd_sc_hd__inv_4 _11309_ (.A(\gpout0.hpos[6] ),
    .Y(_04481_));
 sky130_fd_sc_hd__buf_4 _11310_ (.A(_04453_),
    .X(_04482_));
 sky130_fd_sc_hd__buf_4 _11311_ (.A(\gpout0.hpos[4] ),
    .X(_04483_));
 sky130_fd_sc_hd__buf_4 _11312_ (.A(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__or2_1 _11313_ (.A(_04482_),
    .B(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__inv_2 _11314_ (.A(\rbzero.wall_hot[1] ),
    .Y(_04486_));
 sky130_fd_sc_hd__clkbuf_4 _11315_ (.A(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__nand2_1 _11316_ (.A(_04487_),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04488_));
 sky130_fd_sc_hd__buf_2 _11317_ (.A(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_4 _11318_ (.A(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__nor2_2 _11319_ (.A(_04487_),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04491_));
 sky130_fd_sc_hd__buf_2 _11320_ (.A(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__and2_1 _11321_ (.A(\rbzero.spi_registers.texadd1[19] ),
    .B(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__buf_4 _11322_ (.A(_04487_),
    .X(_04494_));
 sky130_fd_sc_hd__and2_2 _11323_ (.A(\rbzero.wall_hot[1] ),
    .B(\rbzero.wall_hot[0] ),
    .X(_04495_));
 sky130_fd_sc_hd__buf_2 _11324_ (.A(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__clkbuf_4 _11325_ (.A(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__and2_1 _11326_ (.A(_04486_),
    .B(\rbzero.wall_hot[0] ),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_4 _11327_ (.A(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__clkbuf_4 _11328_ (.A(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__a221o_1 _11329_ (.A1(\rbzero.spi_registers.texadd3[19] ),
    .A2(_04494_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[19] ),
    .C1(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__o22a_1 _11330_ (.A1(\rbzero.spi_registers.texadd0[19] ),
    .A2(_04490_),
    .B1(_04493_),
    .B2(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(\rbzero.spi_registers.texadd1[17] ),
    .B(_04492_),
    .X(_04503_));
 sky130_fd_sc_hd__a221o_1 _11332_ (.A1(\rbzero.spi_registers.texadd3[17] ),
    .A2(_04494_),
    .B1(_04496_),
    .B2(\rbzero.spi_registers.texadd2[17] ),
    .C1(_04499_),
    .X(_04504_));
 sky130_fd_sc_hd__o22a_1 _11333_ (.A1(\rbzero.spi_registers.texadd0[17] ),
    .A2(_04490_),
    .B1(_04503_),
    .B2(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__nor2_4 _11334_ (.A(\rbzero.wall_hot[1] ),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04506_));
 sky130_fd_sc_hd__a22o_1 _11335_ (.A1(\rbzero.spi_registers.texadd2[14] ),
    .A2(_04496_),
    .B1(_04506_),
    .B2(\rbzero.spi_registers.texadd3[14] ),
    .X(_04507_));
 sky130_fd_sc_hd__a22o_1 _11336_ (.A1(\rbzero.spi_registers.texadd1[13] ),
    .A2(_04492_),
    .B1(_04506_),
    .B2(\rbzero.spi_registers.texadd3[13] ),
    .X(_04508_));
 sky130_fd_sc_hd__buf_2 _11337_ (.A(\rbzero.side_hot ),
    .X(_04509_));
 sky130_fd_sc_hd__buf_2 _11338_ (.A(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__buf_4 _11339_ (.A(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__and2_1 _11340_ (.A(\rbzero.spi_registers.texadd1[12] ),
    .B(_04492_),
    .X(_04512_));
 sky130_fd_sc_hd__a221o_1 _11341_ (.A1(\rbzero.spi_registers.texadd3[12] ),
    .A2(_04487_),
    .B1(_04496_),
    .B2(\rbzero.spi_registers.texadd2[12] ),
    .C1(_04499_),
    .X(_04513_));
 sky130_fd_sc_hd__o22a_1 _11342_ (.A1(\rbzero.spi_registers.texadd0[12] ),
    .A2(_04489_),
    .B1(_04512_),
    .B2(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__nand2_1 _11343_ (.A(_04511_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__and2_1 _11344_ (.A(\rbzero.spi_registers.texadd1[11] ),
    .B(_04492_),
    .X(_04516_));
 sky130_fd_sc_hd__a221o_1 _11345_ (.A1(\rbzero.spi_registers.texadd3[11] ),
    .A2(_04487_),
    .B1(_04496_),
    .B2(\rbzero.spi_registers.texadd2[11] ),
    .C1(_04499_),
    .X(_04517_));
 sky130_fd_sc_hd__o22a_1 _11346_ (.A1(\rbzero.spi_registers.texadd0[11] ),
    .A2(_04489_),
    .B1(_04516_),
    .B2(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(\rbzero.texu_hot[5] ),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__and2_1 _11348_ (.A(\rbzero.spi_registers.texadd1[10] ),
    .B(_04491_),
    .X(_04520_));
 sky130_fd_sc_hd__a221o_1 _11349_ (.A1(\rbzero.spi_registers.texadd3[10] ),
    .A2(_04487_),
    .B1(_04496_),
    .B2(\rbzero.spi_registers.texadd2[10] ),
    .C1(_04499_),
    .X(_04521_));
 sky130_fd_sc_hd__o22a_1 _11350_ (.A1(\rbzero.spi_registers.texadd0[10] ),
    .A2(_04489_),
    .B1(_04520_),
    .B2(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__nand2_1 _11351_ (.A(\rbzero.texu_hot[4] ),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__a22o_1 _11352_ (.A1(\rbzero.spi_registers.texadd3[9] ),
    .A2(_04487_),
    .B1(_04495_),
    .B2(\rbzero.spi_registers.texadd2[9] ),
    .X(_04524_));
 sky130_fd_sc_hd__a211o_1 _11353_ (.A1(\rbzero.spi_registers.texadd1[9] ),
    .A2(_04491_),
    .B1(_04524_),
    .C1(_04499_),
    .X(_04525_));
 sky130_fd_sc_hd__o21a_1 _11354_ (.A1(\rbzero.spi_registers.texadd0[9] ),
    .A2(_04489_),
    .B1(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__and2_1 _11355_ (.A(\rbzero.texu_hot[3] ),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__a22o_1 _11356_ (.A1(\rbzero.spi_registers.texadd3[8] ),
    .A2(_04487_),
    .B1(_04495_),
    .B2(\rbzero.spi_registers.texadd2[8] ),
    .X(_04528_));
 sky130_fd_sc_hd__a211o_1 _11357_ (.A1(\rbzero.spi_registers.texadd1[8] ),
    .A2(_04491_),
    .B1(_04528_),
    .C1(_04499_),
    .X(_04529_));
 sky130_fd_sc_hd__o21a_1 _11358_ (.A1(\rbzero.spi_registers.texadd0[8] ),
    .A2(_04489_),
    .B1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__nand2_1 _11359_ (.A(\rbzero.texu_hot[2] ),
    .B(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__or2_1 _11360_ (.A(\rbzero.texu_hot[2] ),
    .B(_04530_),
    .X(_04532_));
 sky130_fd_sc_hd__nand2_1 _11361_ (.A(_04531_),
    .B(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__a22o_1 _11362_ (.A1(\rbzero.spi_registers.texadd3[7] ),
    .A2(_04486_),
    .B1(_04495_),
    .B2(\rbzero.spi_registers.texadd2[7] ),
    .X(_04534_));
 sky130_fd_sc_hd__a211o_1 _11363_ (.A1(\rbzero.spi_registers.texadd1[7] ),
    .A2(_04491_),
    .B1(_04534_),
    .C1(_04498_),
    .X(_04535_));
 sky130_fd_sc_hd__o21a_1 _11364_ (.A1(\rbzero.spi_registers.texadd0[7] ),
    .A2(_04488_),
    .B1(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__a22o_1 _11365_ (.A1(\rbzero.spi_registers.texadd3[6] ),
    .A2(_04487_),
    .B1(_04495_),
    .B2(\rbzero.spi_registers.texadd2[6] ),
    .X(_04537_));
 sky130_fd_sc_hd__a211o_1 _11366_ (.A1(\rbzero.spi_registers.texadd1[6] ),
    .A2(_04491_),
    .B1(_04537_),
    .C1(_04498_),
    .X(_04538_));
 sky130_fd_sc_hd__o21a_1 _11367_ (.A1(\rbzero.spi_registers.texadd0[6] ),
    .A2(_04489_),
    .B1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__nand2_1 _11368_ (.A(\rbzero.texu_hot[0] ),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__xnor2_1 _11369_ (.A(\rbzero.texu_hot[1] ),
    .B(_04536_),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_1 _11370_ (.A(_04540_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__a21o_1 _11371_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_04536_),
    .B1(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__or2b_1 _11372_ (.A(_04533_),
    .B_N(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__nor2_1 _11373_ (.A(\rbzero.texu_hot[3] ),
    .B(_04526_),
    .Y(_04545_));
 sky130_fd_sc_hd__or2_1 _11374_ (.A(_04527_),
    .B(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__a21oi_1 _11375_ (.A1(_04531_),
    .A2(_04544_),
    .B1(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__or2_1 _11376_ (.A(\rbzero.texu_hot[4] ),
    .B(_04522_),
    .X(_04548_));
 sky130_fd_sc_hd__and2_1 _11377_ (.A(_04523_),
    .B(_04548_),
    .X(_04549_));
 sky130_fd_sc_hd__o21ai_1 _11378_ (.A1(_04527_),
    .A2(_04547_),
    .B1(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__or2_1 _11379_ (.A(\rbzero.texu_hot[5] ),
    .B(_04518_),
    .X(_04551_));
 sky130_fd_sc_hd__nand2_1 _11380_ (.A(_04519_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a21o_1 _11381_ (.A1(_04523_),
    .A2(_04550_),
    .B1(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__or2_1 _11382_ (.A(_04511_),
    .B(_04514_),
    .X(_04554_));
 sky130_fd_sc_hd__nand2_1 _11383_ (.A(_04515_),
    .B(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__a21o_1 _11384_ (.A1(_04519_),
    .A2(_04553_),
    .B1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__nor2_1 _11385_ (.A(\rbzero.spi_registers.texadd0[13] ),
    .B(_04489_),
    .Y(_04557_));
 sky130_fd_sc_hd__and2b_1 _11386_ (.A_N(\rbzero.spi_registers.texadd2[13] ),
    .B(_04496_),
    .X(_04558_));
 sky130_fd_sc_hd__a2111oi_2 _11387_ (.A1(_04515_),
    .A2(_04556_),
    .B1(_04557_),
    .C1(_04558_),
    .D1(_04508_),
    .Y(_04559_));
 sky130_fd_sc_hd__or2_1 _11388_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_04489_),
    .X(_04560_));
 sky130_fd_sc_hd__inv_2 _11389_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .Y(_04561_));
 sky130_fd_sc_hd__a21oi_1 _11390_ (.A1(_04561_),
    .A2(_04492_),
    .B1(_04507_),
    .Y(_04562_));
 sky130_fd_sc_hd__o211a_1 _11391_ (.A1(_04508_),
    .A2(_04559_),
    .B1(_04560_),
    .C1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__and2_1 _11392_ (.A(\rbzero.spi_registers.texadd1[15] ),
    .B(_04492_),
    .X(_04564_));
 sky130_fd_sc_hd__a221o_1 _11393_ (.A1(\rbzero.spi_registers.texadd3[15] ),
    .A2(_04487_),
    .B1(_04496_),
    .B2(\rbzero.spi_registers.texadd2[15] ),
    .C1(_04499_),
    .X(_04565_));
 sky130_fd_sc_hd__o22a_1 _11394_ (.A1(\rbzero.spi_registers.texadd0[15] ),
    .A2(_04489_),
    .B1(_04564_),
    .B2(_04565_),
    .X(_04566_));
 sky130_fd_sc_hd__o21a_1 _11395_ (.A1(_04507_),
    .A2(_04563_),
    .B1(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__a22o_1 _11396_ (.A1(\rbzero.spi_registers.texadd3[16] ),
    .A2(_04494_),
    .B1(_04496_),
    .B2(\rbzero.spi_registers.texadd2[16] ),
    .X(_04568_));
 sky130_fd_sc_hd__a211o_1 _11397_ (.A1(\rbzero.spi_registers.texadd1[16] ),
    .A2(_04492_),
    .B1(_04568_),
    .C1(_04499_),
    .X(_04569_));
 sky130_fd_sc_hd__o21a_1 _11398_ (.A1(\rbzero.spi_registers.texadd0[16] ),
    .A2(_04490_),
    .B1(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__and3_1 _11399_ (.A(_04505_),
    .B(_04567_),
    .C(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__a22o_1 _11400_ (.A1(\rbzero.spi_registers.texadd3[18] ),
    .A2(_04494_),
    .B1(_04496_),
    .B2(\rbzero.spi_registers.texadd2[18] ),
    .X(_04572_));
 sky130_fd_sc_hd__a211o_1 _11401_ (.A1(\rbzero.spi_registers.texadd1[18] ),
    .A2(_04492_),
    .B1(_04572_),
    .C1(_04499_),
    .X(_04573_));
 sky130_fd_sc_hd__o21a_1 _11402_ (.A1(\rbzero.spi_registers.texadd0[18] ),
    .A2(_04490_),
    .B1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__and2_1 _11403_ (.A(_04571_),
    .B(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__inv_4 _11404_ (.A(\gpout0.hpos[0] ),
    .Y(_04576_));
 sky130_fd_sc_hd__nor3_1 _11405_ (.A(_04576_),
    .B(_04571_),
    .C(_04574_),
    .Y(_04577_));
 sky130_fd_sc_hd__o22a_1 _11406_ (.A1(_04012_),
    .A2(_04502_),
    .B1(_04575_),
    .B2(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__clkinv_4 _11407_ (.A(\gpout0.hpos[1] ),
    .Y(_04579_));
 sky130_fd_sc_hd__o31ai_1 _11408_ (.A1(_04012_),
    .A2(_04502_),
    .A3(_04575_),
    .B1(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__and2_1 _11409_ (.A(_04567_),
    .B(_04570_),
    .X(_04581_));
 sky130_fd_sc_hd__nor3_1 _11410_ (.A(_04576_),
    .B(_04567_),
    .C(_04570_),
    .Y(_04582_));
 sky130_fd_sc_hd__o22a_1 _11411_ (.A1(_04012_),
    .A2(_04505_),
    .B1(_04581_),
    .B2(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__buf_4 _11412_ (.A(\gpout0.hpos[1] ),
    .X(_04584_));
 sky130_fd_sc_hd__clkbuf_4 _11413_ (.A(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__o31ai_1 _11414_ (.A1(_04012_),
    .A2(_04505_),
    .A3(_04581_),
    .B1(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__buf_4 _11415_ (.A(\gpout0.hpos[2] ),
    .X(_04587_));
 sky130_fd_sc_hd__o221a_1 _11416_ (.A1(_04578_),
    .A2(_04580_),
    .B1(_04583_),
    .B2(_04586_),
    .C1(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__or2_1 _11417_ (.A(\rbzero.spi_registers.texadd0[23] ),
    .B(_04490_),
    .X(_04589_));
 sky130_fd_sc_hd__clkbuf_4 _11418_ (.A(_04492_),
    .X(_04590_));
 sky130_fd_sc_hd__a22o_1 _11419_ (.A1(\rbzero.spi_registers.texadd3[23] ),
    .A2(_04494_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[23] ),
    .X(_04591_));
 sky130_fd_sc_hd__a211o_1 _11420_ (.A1(\rbzero.spi_registers.texadd1[23] ),
    .A2(_04590_),
    .B1(_04591_),
    .C1(_04500_),
    .X(_04592_));
 sky130_fd_sc_hd__a21oi_1 _11421_ (.A1(_04589_),
    .A2(_04592_),
    .B1(_04012_),
    .Y(_04593_));
 sky130_fd_sc_hd__o21a_1 _11422_ (.A1(\rbzero.spi_registers.texadd2[22] ),
    .A2(_04494_),
    .B1(\rbzero.wall_hot[0] ),
    .X(_04594_));
 sky130_fd_sc_hd__a221o_1 _11423_ (.A1(\rbzero.spi_registers.texadd3[22] ),
    .A2(_04494_),
    .B1(_04590_),
    .B2(\rbzero.spi_registers.texadd1[22] ),
    .C1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__o21ai_1 _11424_ (.A1(\rbzero.spi_registers.texadd0[22] ),
    .A2(_04490_),
    .B1(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__nand2_1 _11425_ (.A(_04011_),
    .B(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__a22o_1 _11426_ (.A1(\rbzero.spi_registers.texadd3[20] ),
    .A2(_04494_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[20] ),
    .X(_04598_));
 sky130_fd_sc_hd__a211o_1 _11427_ (.A1(\rbzero.spi_registers.texadd1[20] ),
    .A2(_04590_),
    .B1(_04598_),
    .C1(_04500_),
    .X(_04599_));
 sky130_fd_sc_hd__o21a_1 _11428_ (.A1(\rbzero.spi_registers.texadd0[20] ),
    .A2(_04490_),
    .B1(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__and3_1 _11429_ (.A(_04502_),
    .B(_04575_),
    .C(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__a22o_1 _11430_ (.A1(\rbzero.spi_registers.texadd3[21] ),
    .A2(_04494_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[21] ),
    .X(_04602_));
 sky130_fd_sc_hd__a211o_1 _11431_ (.A1(\rbzero.spi_registers.texadd1[21] ),
    .A2(_04590_),
    .B1(_04602_),
    .C1(_04500_),
    .X(_04603_));
 sky130_fd_sc_hd__o21a_1 _11432_ (.A1(\rbzero.spi_registers.texadd0[21] ),
    .A2(_04490_),
    .B1(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__nand2_1 _11433_ (.A(_04601_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__mux2_1 _11434_ (.A0(_04596_),
    .A1(_04597_),
    .S(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__or2_1 _11435_ (.A(_04593_),
    .B(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__a21oi_1 _11436_ (.A1(_04593_),
    .A2(_04606_),
    .B1(_04585_),
    .Y(_04608_));
 sky130_fd_sc_hd__a211oi_1 _11437_ (.A1(_04502_),
    .A2(_04575_),
    .B1(_04600_),
    .C1(_04576_),
    .Y(_04609_));
 sky130_fd_sc_hd__o22a_1 _11438_ (.A1(_04011_),
    .A2(_04604_),
    .B1(_04609_),
    .B2(_04601_),
    .X(_04610_));
 sky130_fd_sc_hd__or3_1 _11439_ (.A(_04011_),
    .B(_04601_),
    .C(_04604_),
    .X(_04611_));
 sky130_fd_sc_hd__and3b_1 _11440_ (.A_N(_04610_),
    .B(_04611_),
    .C(_04585_),
    .X(_04612_));
 sky130_fd_sc_hd__a211o_1 _11441_ (.A1(_04607_),
    .A2(_04608_),
    .B1(_04612_),
    .C1(_04587_),
    .X(_04613_));
 sky130_fd_sc_hd__nor4b_1 _11442_ (.A(_04481_),
    .B(_04485_),
    .C(_04588_),
    .D_N(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__inv_2 _11443_ (.A(\gpout0.hpos[2] ),
    .Y(_04615_));
 sky130_fd_sc_hd__nand2_2 _11444_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .Y(_04616_));
 sky130_fd_sc_hd__or2_4 _11445_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .X(_04617_));
 sky130_fd_sc_hd__a21oi_1 _11446_ (.A1(_04579_),
    .A2(_04012_),
    .B1(_04615_),
    .Y(_04618_));
 sky130_fd_sc_hd__a31o_1 _11447_ (.A1(_04615_),
    .A2(_04616_),
    .A3(_04617_),
    .B1(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__nand3_1 _11448_ (.A(_04552_),
    .B(_04523_),
    .C(_04550_),
    .Y(_04620_));
 sky130_fd_sc_hd__or3_1 _11449_ (.A(_04549_),
    .B(_04527_),
    .C(_04547_),
    .X(_04621_));
 sky130_fd_sc_hd__a31o_1 _11450_ (.A1(_04011_),
    .A2(_04550_),
    .A3(_04621_),
    .B1(_04585_),
    .X(_04622_));
 sky130_fd_sc_hd__a31o_1 _11451_ (.A1(_04576_),
    .A2(_04553_),
    .A3(_04620_),
    .B1(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__xnor2_1 _11452_ (.A(_04533_),
    .B(_04543_),
    .Y(_04624_));
 sky130_fd_sc_hd__and3_1 _11453_ (.A(_04531_),
    .B(_04544_),
    .C(_04546_),
    .X(_04625_));
 sky130_fd_sc_hd__o31a_1 _11454_ (.A1(_04011_),
    .A2(_04547_),
    .A3(_04625_),
    .B1(_04585_),
    .X(_04626_));
 sky130_fd_sc_hd__a21bo_1 _11455_ (.A1(_04011_),
    .A2(_04624_),
    .B1_N(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__a211o_1 _11456_ (.A1(_04560_),
    .A2(_04562_),
    .B1(_04508_),
    .C1(_04559_),
    .X(_04628_));
 sky130_fd_sc_hd__or3b_1 _11457_ (.A(_04585_),
    .B(_04563_),
    .C_N(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _11458_ (.A(_04585_),
    .B(_04556_),
    .Y(_04630_));
 sky130_fd_sc_hd__a31o_1 _11459_ (.A1(_04555_),
    .A2(_04519_),
    .A3(_04553_),
    .B1(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__nor3_1 _11460_ (.A(_04507_),
    .B(_04563_),
    .C(_04566_),
    .Y(_04632_));
 sky130_fd_sc_hd__o311a_1 _11461_ (.A1(_04508_),
    .A2(_04557_),
    .A3(_04558_),
    .B1(_04515_),
    .C1(_04556_),
    .X(_04633_));
 sky130_fd_sc_hd__or3_1 _11462_ (.A(_04579_),
    .B(_04559_),
    .C(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__o311a_1 _11463_ (.A1(_04585_),
    .A2(_04567_),
    .A3(_04632_),
    .B1(_04634_),
    .C1(_04576_),
    .X(_04635_));
 sky130_fd_sc_hd__a311oi_2 _11464_ (.A1(_04012_),
    .A2(_04629_),
    .A3(_04631_),
    .B1(_04635_),
    .C1(_04587_),
    .Y(_04636_));
 sky130_fd_sc_hd__a311o_1 _11465_ (.A1(_04587_),
    .A2(_04623_),
    .A3(_04627_),
    .B1(_04484_),
    .C1(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__or2_1 _11466_ (.A(\rbzero.texu_hot[0] ),
    .B(_04539_),
    .X(_04638_));
 sky130_fd_sc_hd__a31o_1 _11467_ (.A1(_04011_),
    .A2(_04540_),
    .A3(_04638_),
    .B1(_04585_),
    .X(_04639_));
 sky130_fd_sc_hd__or2_1 _11468_ (.A(_04010_),
    .B(_04542_),
    .X(_04640_));
 sky130_fd_sc_hd__a21oi_1 _11469_ (.A1(_04540_),
    .A2(_04541_),
    .B1(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__a22o_1 _11470_ (.A1(\rbzero.spi_registers.texadd1[5] ),
    .A2(_04590_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[5] ),
    .X(_04642_));
 sky130_fd_sc_hd__a221o_1 _11471_ (.A1(\rbzero.spi_registers.texadd0[5] ),
    .A2(_04500_),
    .B1(_04506_),
    .B2(\rbzero.spi_registers.texadd3[5] ),
    .C1(_04010_),
    .X(_04643_));
 sky130_fd_sc_hd__a221o_1 _11472_ (.A1(\rbzero.spi_registers.texadd0[4] ),
    .A2(_04500_),
    .B1(_04506_),
    .B2(\rbzero.spi_registers.texadd3[4] ),
    .C1(_04576_),
    .X(_04644_));
 sky130_fd_sc_hd__a22o_1 _11473_ (.A1(\rbzero.spi_registers.texadd1[4] ),
    .A2(_04590_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[4] ),
    .X(_04645_));
 sky130_fd_sc_hd__o22a_1 _11474_ (.A1(_04642_),
    .A2(_04643_),
    .B1(_04644_),
    .B2(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__o22a_1 _11475_ (.A1(_04639_),
    .A2(_04641_),
    .B1(_04646_),
    .B2(_04579_),
    .X(_04647_));
 sky130_fd_sc_hd__a22o_1 _11476_ (.A1(\rbzero.spi_registers.texadd2[1] ),
    .A2(_04497_),
    .B1(_04506_),
    .B2(\rbzero.spi_registers.texadd3[1] ),
    .X(_04648_));
 sky130_fd_sc_hd__a211o_1 _11477_ (.A1(\rbzero.spi_registers.texadd1[1] ),
    .A2(_04590_),
    .B1(_04648_),
    .C1(_04500_),
    .X(_04649_));
 sky130_fd_sc_hd__o211a_1 _11478_ (.A1(\rbzero.spi_registers.texadd0[1] ),
    .A2(_04490_),
    .B1(_04649_),
    .C1(_04576_),
    .X(_04650_));
 sky130_fd_sc_hd__a22o_1 _11479_ (.A1(\rbzero.spi_registers.texadd2[0] ),
    .A2(_04497_),
    .B1(_04506_),
    .B2(\rbzero.spi_registers.texadd3[0] ),
    .X(_04651_));
 sky130_fd_sc_hd__a211o_1 _11480_ (.A1(\rbzero.spi_registers.texadd1[0] ),
    .A2(_04590_),
    .B1(_04651_),
    .C1(_04500_),
    .X(_04652_));
 sky130_fd_sc_hd__o211a_1 _11481_ (.A1(\rbzero.spi_registers.texadd0[0] ),
    .A2(_04490_),
    .B1(_04652_),
    .C1(_04011_),
    .X(_04653_));
 sky130_fd_sc_hd__or3_1 _11482_ (.A(_04579_),
    .B(_04650_),
    .C(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__and2_1 _11483_ (.A(\rbzero.spi_registers.texadd3[3] ),
    .B(_04506_),
    .X(_04655_));
 sky130_fd_sc_hd__a221o_1 _11484_ (.A1(\rbzero.spi_registers.texadd1[3] ),
    .A2(_04590_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[3] ),
    .C1(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__a211o_1 _11485_ (.A1(\rbzero.spi_registers.texadd0[3] ),
    .A2(_04500_),
    .B1(_04617_),
    .C1(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__a211o_1 _11486_ (.A1(\rbzero.spi_registers.texadd0[2] ),
    .A2(_04500_),
    .B1(_04576_),
    .C1(_04584_),
    .X(_04658_));
 sky130_fd_sc_hd__a22o_1 _11487_ (.A1(\rbzero.spi_registers.texadd1[2] ),
    .A2(_04590_),
    .B1(_04497_),
    .B2(\rbzero.spi_registers.texadd2[2] ),
    .X(_04659_));
 sky130_fd_sc_hd__a211o_1 _11488_ (.A1(\rbzero.spi_registers.texadd3[2] ),
    .A2(_04506_),
    .B1(_04658_),
    .C1(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__and3_1 _11489_ (.A(_04587_),
    .B(_04657_),
    .C(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__a221o_1 _11490_ (.A1(_04615_),
    .A2(_04647_),
    .B1(_04654_),
    .B2(_04661_),
    .C1(_04482_),
    .X(_04662_));
 sky130_fd_sc_hd__and4b_1 _11491_ (.A_N(_04456_),
    .B(_04637_),
    .C(_04662_),
    .D(_04458_),
    .X(_04663_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(_04456_),
    .A2(_04619_),
    .B1(_04663_),
    .B2(_04485_),
    .X(_04664_));
 sky130_fd_sc_hd__o21ba_2 _11493_ (.A1(_04614_),
    .A2(_04664_),
    .B1_N(net73),
    .X(net74));
 sky130_fd_sc_hd__inv_2 _20689__4 (.A(clknet_1_1__leaf__03609_),
    .Y(net130));
 sky130_fd_sc_hd__nor2_4 _11495_ (.A(_04615_),
    .B(_04616_),
    .Y(_04665_));
 sky130_fd_sc_hd__and2_1 _11496_ (.A(\gpout0.hpos[3] ),
    .B(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__or2_1 _11497_ (.A(\gpout0.hpos[4] ),
    .B(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__o21a_1 _11498_ (.A1(\gpout0.hpos[5] ),
    .A2(_04667_),
    .B1(\gpout0.hpos[6] ),
    .X(_04668_));
 sky130_fd_sc_hd__and2_1 _11499_ (.A(\gpout0.hpos[7] ),
    .B(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__a21oi_2 _11500_ (.A1(_04016_),
    .A2(_04669_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04670_));
 sky130_fd_sc_hd__clkbuf_4 _11501_ (.A(\gpout0.vpos[7] ),
    .X(_04671_));
 sky130_fd_sc_hd__clkinv_4 _11502_ (.A(net3),
    .Y(_04672_));
 sky130_fd_sc_hd__or4_1 _11503_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.vpos[8] ),
    .C(_04671_),
    .D(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__inv_2 _11504_ (.A(\gpout0.vpos[1] ),
    .Y(_04674_));
 sky130_fd_sc_hd__buf_2 _11505_ (.A(\gpout0.vpos[2] ),
    .X(_04675_));
 sky130_fd_sc_hd__nor2_1 _11506_ (.A(_04675_),
    .B(\gpout0.vpos[0] ),
    .Y(_04676_));
 sky130_fd_sc_hd__nand2_2 _11507_ (.A(_04674_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__buf_4 _11508_ (.A(\gpout0.vpos[3] ),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_4 _11509_ (.A(\gpout0.vpos[5] ),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_4 _11510_ (.A(\gpout0.vpos[4] ),
    .X(_04680_));
 sky130_fd_sc_hd__or2_4 _11511_ (.A(_04679_),
    .B(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__or2_1 _11512_ (.A(_04678_),
    .B(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_4 _11513_ (.A(\gpout0.vpos[6] ),
    .X(_04683_));
 sky130_fd_sc_hd__o21a_1 _11514_ (.A1(_04677_),
    .A2(_04682_),
    .B1(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__nor3_4 _11515_ (.A(_04670_),
    .B(_04673_),
    .C(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__inv_2 _11516_ (.A(net2),
    .Y(_04686_));
 sky130_fd_sc_hd__and3_2 _11517_ (.A(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .C(_04472_),
    .X(_04687_));
 sky130_fd_sc_hd__a21oi_2 _11518_ (.A1(\rbzero.trace_state[0] ),
    .A2(_04687_),
    .B1(_04686_),
    .Y(_04688_));
 sky130_fd_sc_hd__or2_1 _11519_ (.A(\gpout0.hpos[2] ),
    .B(_04617_),
    .X(_04689_));
 sky130_fd_sc_hd__nor2_1 _11520_ (.A(_04482_),
    .B(_04483_),
    .Y(_04690_));
 sky130_fd_sc_hd__or2_1 _11521_ (.A(_04013_),
    .B(_04457_),
    .X(_04691_));
 sky130_fd_sc_hd__nor2_1 _11522_ (.A(_04452_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(_04690_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__o21a_1 _11524_ (.A1(_04689_),
    .A2(_04693_),
    .B1(_04016_),
    .X(_04694_));
 sky130_fd_sc_hd__or3b_1 _11525_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.hpos[9] ),
    .C_N(net1),
    .X(_04695_));
 sky130_fd_sc_hd__nor2_1 _11526_ (.A(\gpout0.vpos[7] ),
    .B(_04678_),
    .Y(_04696_));
 sky130_fd_sc_hd__or3b_1 _11527_ (.A(\gpout0.vpos[6] ),
    .B(_04681_),
    .C_N(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__o21a_1 _11528_ (.A1(_04677_),
    .A2(_04697_),
    .B1(\gpout0.vpos[8] ),
    .X(_04698_));
 sky130_fd_sc_hd__nor3_2 _11529_ (.A(_04694_),
    .B(_04695_),
    .C(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21oi_4 _11530_ (.A1(_04016_),
    .A2(_04691_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04700_));
 sky130_fd_sc_hd__mux2_1 _11531_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__buf_4 _11532_ (.A(\rbzero.row_render.side ),
    .X(_04702_));
 sky130_fd_sc_hd__nand2b_2 _11533_ (.A_N(\rbzero.row_render.wall[1] ),
    .B(\rbzero.row_render.wall[0] ),
    .Y(_04703_));
 sky130_fd_sc_hd__clkbuf_8 _11534_ (.A(net42),
    .X(_04704_));
 sky130_fd_sc_hd__o21ai_1 _11535_ (.A1(_04702_),
    .A2(_04703_),
    .B1(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__and2b_2 _11536_ (.A_N(\rbzero.row_render.wall[0] ),
    .B(\rbzero.row_render.wall[1] ),
    .X(_04706_));
 sky130_fd_sc_hd__nand2_1 _11537_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .Y(_04707_));
 sky130_fd_sc_hd__or2_1 _11538_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .X(_04708_));
 sky130_fd_sc_hd__nand3_1 _11539_ (.A(\rbzero.texV[6] ),
    .B(_04707_),
    .C(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__a21o_1 _11540_ (.A1(_04707_),
    .A2(_04708_),
    .B1(\rbzero.texV[6] ),
    .X(_04710_));
 sky130_fd_sc_hd__nand2_1 _11541_ (.A(_04709_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__and2_1 _11542_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .X(_04712_));
 sky130_fd_sc_hd__nor2_1 _11543_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .Y(_04713_));
 sky130_fd_sc_hd__nor2_1 _11544_ (.A(_04712_),
    .B(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__a21oi_2 _11545_ (.A1(\rbzero.texV[5] ),
    .A2(_04714_),
    .B1(_04712_),
    .Y(_04715_));
 sky130_fd_sc_hd__xnor2_1 _11546_ (.A(_04711_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_1 _11547_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .Y(_04717_));
 sky130_fd_sc_hd__or2_1 _11548_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .X(_04718_));
 sky130_fd_sc_hd__nand3_1 _11549_ (.A(\rbzero.texV[4] ),
    .B(_04717_),
    .C(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__xnor2_1 _11550_ (.A(\rbzero.texV[5] ),
    .B(_04714_),
    .Y(_04720_));
 sky130_fd_sc_hd__a21oi_1 _11551_ (.A1(_04717_),
    .A2(_04719_),
    .B1(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__a21o_1 _11552_ (.A1(_04717_),
    .A2(_04718_),
    .B1(\rbzero.texV[4] ),
    .X(_04722_));
 sky130_fd_sc_hd__nand2_1 _11553_ (.A(_04719_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__or2_1 _11554_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .X(_04724_));
 sky130_fd_sc_hd__nand2_1 _11555_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .Y(_04725_));
 sky130_fd_sc_hd__a21boi_1 _11556_ (.A1(\rbzero.texV[3] ),
    .A2(_04724_),
    .B1_N(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__or2_1 _11557_ (.A(_04723_),
    .B(_04726_),
    .X(_04727_));
 sky130_fd_sc_hd__xnor2_1 _11558_ (.A(_04723_),
    .B(_04726_),
    .Y(_04728_));
 sky130_fd_sc_hd__nand2_1 _11559_ (.A(_04725_),
    .B(_04724_),
    .Y(_04729_));
 sky130_fd_sc_hd__xor2_1 _11560_ (.A(\rbzero.texV[3] ),
    .B(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__o211a_1 _11561_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(\rbzero.texV[1] ),
    .B1(\rbzero.texV[0] ),
    .C1(\rbzero.traced_texVinit[0] ),
    .X(_04731_));
 sky130_fd_sc_hd__a221o_1 _11562_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(\rbzero.texV[1] ),
    .B2(\rbzero.traced_texVinit[1] ),
    .C1(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__o21ai_1 _11563_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__or2_1 _11564_ (.A(_04730_),
    .B(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__or2_2 _11565_ (.A(_04728_),
    .B(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__and3_1 _11566_ (.A(_04720_),
    .B(_04717_),
    .C(_04719_),
    .X(_04736_));
 sky130_fd_sc_hd__or2_1 _11567_ (.A(_04721_),
    .B(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__a21oi_2 _11568_ (.A1(_04727_),
    .A2(_04735_),
    .B1(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__nor2_1 _11569_ (.A(_04721_),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__nor2_1 _11570_ (.A(_04716_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__nand2_1 _11571_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_04741_));
 sky130_fd_sc_hd__xor2_1 _11572_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .X(_04742_));
 sky130_fd_sc_hd__xnor2_1 _11573_ (.A(_04741_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__or2_1 _11574_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .X(_04744_));
 sky130_fd_sc_hd__nand2_1 _11575_ (.A(_04741_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__or2_1 _11576_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .X(_04746_));
 sky130_fd_sc_hd__nand2_1 _11577_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .Y(_04747_));
 sky130_fd_sc_hd__a21boi_1 _11578_ (.A1(\rbzero.texV[8] ),
    .A2(_04746_),
    .B1_N(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__nor2_1 _11579_ (.A(_04745_),
    .B(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__nand2_1 _11580_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .Y(_04750_));
 sky130_fd_sc_hd__or2_1 _11581_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .X(_04751_));
 sky130_fd_sc_hd__nand3_1 _11582_ (.A(\rbzero.texV[7] ),
    .B(_04750_),
    .C(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _11583_ (.A(_04747_),
    .B(_04746_),
    .Y(_04753_));
 sky130_fd_sc_hd__xor2_1 _11584_ (.A(\rbzero.texV[8] ),
    .B(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__a21oi_1 _11585_ (.A1(_04750_),
    .A2(_04752_),
    .B1(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__and3_1 _11586_ (.A(_04754_),
    .B(_04750_),
    .C(_04752_),
    .X(_04756_));
 sky130_fd_sc_hd__a21o_1 _11587_ (.A1(_04750_),
    .A2(_04751_),
    .B1(\rbzero.texV[7] ),
    .X(_04757_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(_04752_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand3_2 _11589_ (.A(_04758_),
    .B(_04707_),
    .C(_04709_),
    .Y(_04759_));
 sky130_fd_sc_hd__o21bai_4 _11590_ (.A1(_04711_),
    .A2(_04715_),
    .B1_N(_04740_),
    .Y(_04760_));
 sky130_fd_sc_hd__a21oi_2 _11591_ (.A1(_04707_),
    .A2(_04709_),
    .B1(_04758_),
    .Y(_04761_));
 sky130_fd_sc_hd__a21oi_4 _11592_ (.A1(_04759_),
    .A2(_04760_),
    .B1(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__nor2_1 _11593_ (.A(_04756_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__nand2_1 _11594_ (.A(_04745_),
    .B(_04748_),
    .Y(_04764_));
 sky130_fd_sc_hd__o31a_1 _11595_ (.A1(_04749_),
    .A2(_04755_),
    .A3(_04763_),
    .B1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a21oi_1 _11596_ (.A1(_04743_),
    .A2(_04765_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04766_));
 sky130_fd_sc_hd__o21a_1 _11597_ (.A1(_04743_),
    .A2(_04765_),
    .B1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__buf_6 _11598_ (.A(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__and2_1 _11599_ (.A(_04716_),
    .B(_04739_),
    .X(_04769_));
 sky130_fd_sc_hd__nor3_4 _11600_ (.A(_04740_),
    .B(_04768_),
    .C(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__and3_1 _11601_ (.A(_04737_),
    .B(_04727_),
    .C(_04735_),
    .X(_04771_));
 sky130_fd_sc_hd__nor3_4 _11602_ (.A(_04738_),
    .B(_04768_),
    .C(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__buf_6 _11603_ (.A(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__a21oi_1 _11604_ (.A1(_04728_),
    .A2(_04734_),
    .B1(_04768_),
    .Y(_04774_));
 sky130_fd_sc_hd__and2_2 _11605_ (.A(_04735_),
    .B(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__buf_4 _11606_ (.A(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__clkbuf_8 _11607_ (.A(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__nor2_1 _11608_ (.A(\rbzero.row_render.texu[2] ),
    .B(\rbzero.row_render.texu[1] ),
    .Y(_04778_));
 sky130_fd_sc_hd__inv_2 _11609_ (.A(\rbzero.row_render.texu[3] ),
    .Y(_04779_));
 sky130_fd_sc_hd__a32o_1 _11610_ (.A1(_04770_),
    .A2(_04773_),
    .A3(_04777_),
    .B1(_04778_),
    .B2(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__inv_2 _11611_ (.A(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__or3_1 _11612_ (.A(_04740_),
    .B(_04768_),
    .C(_04769_),
    .X(_04782_));
 sky130_fd_sc_hd__buf_6 _11613_ (.A(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__or3_1 _11614_ (.A(_04738_),
    .B(_04768_),
    .C(_04771_),
    .X(_04784_));
 sky130_fd_sc_hd__buf_6 _11615_ (.A(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__buf_6 _11616_ (.A(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__nand2_2 _11617_ (.A(_04735_),
    .B(_04774_),
    .Y(_04787_));
 sky130_fd_sc_hd__buf_4 _11618_ (.A(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__buf_4 _11619_ (.A(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__and3_1 _11620_ (.A(_04783_),
    .B(_04786_),
    .C(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__a31o_1 _11621_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(\rbzero.row_render.texu[2] ),
    .A3(\rbzero.row_render.texu[1] ),
    .B1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__and4_1 _11622_ (.A(\rbzero.row_render.wall[0] ),
    .B(\rbzero.row_render.wall[1] ),
    .C(_04781_),
    .D(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__xnor2_1 _11623_ (.A(_04702_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__nor2_8 _11624_ (.A(_04772_),
    .B(_04776_),
    .Y(_04794_));
 sky130_fd_sc_hd__inv_2 _11625_ (.A(_04734_),
    .Y(_04795_));
 sky130_fd_sc_hd__and2_1 _11626_ (.A(_04730_),
    .B(_04733_),
    .X(_04796_));
 sky130_fd_sc_hd__nor3_4 _11627_ (.A(_04795_),
    .B(_04768_),
    .C(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__buf_4 _11628_ (.A(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__buf_4 _11629_ (.A(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__nor2_1 _11630_ (.A(\rbzero.row_render.texu[0] ),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__inv_2 _11631_ (.A(\rbzero.row_render.texu[4] ),
    .Y(_04801_));
 sky130_fd_sc_hd__a41o_1 _11632_ (.A1(_04801_),
    .A2(_04779_),
    .A3(\rbzero.row_render.texu[2] ),
    .A4(\rbzero.row_render.texu[1] ),
    .B1(_04770_),
    .X(_04802_));
 sky130_fd_sc_hd__a31o_1 _11633_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(\rbzero.row_render.texu[3] ),
    .A3(_04778_),
    .B1(_04783_),
    .X(_04803_));
 sky130_fd_sc_hd__and3b_1 _11634_ (.A_N(\rbzero.row_render.texu[0] ),
    .B(_04802_),
    .C(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__a21o_1 _11635_ (.A1(_04794_),
    .A2(_04800_),
    .B1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__or2_1 _11636_ (.A(\rbzero.row_render.side ),
    .B(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__buf_6 _11637_ (.A(_04794_),
    .X(_04807_));
 sky130_fd_sc_hd__or3_1 _11638_ (.A(_04795_),
    .B(_04767_),
    .C(_04796_),
    .X(_04808_));
 sky130_fd_sc_hd__buf_2 _11639_ (.A(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__buf_4 _11640_ (.A(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__buf_4 _11641_ (.A(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__buf_6 _11642_ (.A(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__clkbuf_8 _11643_ (.A(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__inv_2 _11644_ (.A(_04702_),
    .Y(_04814_));
 sky130_fd_sc_hd__a31o_1 _11645_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04807_),
    .A3(_04813_),
    .B1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__nand3_1 _11646_ (.A(_04706_),
    .B(_04806_),
    .C(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__o211a_1 _11647_ (.A1(_04706_),
    .A2(_04793_),
    .B1(_04816_),
    .C1(_04703_),
    .X(_04817_));
 sky130_fd_sc_hd__clkinv_4 _11648_ (.A(net42),
    .Y(_04818_));
 sky130_fd_sc_hd__or2_2 _11649_ (.A(_04756_),
    .B(_04755_),
    .X(_04819_));
 sky130_fd_sc_hd__xnor2_4 _11650_ (.A(_04762_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__nor2_8 _11651_ (.A(_04768_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__inv_2 _11652_ (.A(_04759_),
    .Y(_04822_));
 sky130_fd_sc_hd__nor2_2 _11653_ (.A(_04822_),
    .B(_04761_),
    .Y(_04823_));
 sky130_fd_sc_hd__xnor2_4 _11654_ (.A(_04760_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__nor2_8 _11655_ (.A(_04768_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__buf_6 _11656_ (.A(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__buf_6 _11657_ (.A(_04786_),
    .X(_04827_));
 sky130_fd_sc_hd__buf_6 _11658_ (.A(_04809_),
    .X(_04828_));
 sky130_fd_sc_hd__buf_4 _11659_ (.A(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__buf_4 _11660_ (.A(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__clkbuf_8 _11662_ (.A(_04809_),
    .X(_04832_));
 sky130_fd_sc_hd__buf_4 _11663_ (.A(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_8 _11665_ (.A(_04776_),
    .X(_04835_));
 sky130_fd_sc_hd__buf_6 _11666_ (.A(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__mux2_1 _11667_ (.A0(_04831_),
    .A1(_04834_),
    .S(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_4 _11668_ (.A(_04787_),
    .X(_04838_));
 sky130_fd_sc_hd__clkbuf_4 _11669_ (.A(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__buf_4 _11670_ (.A(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__buf_6 _11671_ (.A(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__buf_4 _11672_ (.A(_04829_),
    .X(_04842_));
 sky130_fd_sc_hd__mux2_1 _11673_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__buf_6 _11674_ (.A(_04776_),
    .X(_04844_));
 sky130_fd_sc_hd__mux2_1 _11675_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04832_),
    .X(_04845_));
 sky130_fd_sc_hd__or2_1 _11676_ (.A(_04844_),
    .B(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__buf_6 _11677_ (.A(_04773_),
    .X(_04847_));
 sky130_fd_sc_hd__o211a_1 _11678_ (.A1(_04841_),
    .A2(_04843_),
    .B1(_04846_),
    .C1(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__buf_6 _11679_ (.A(_04783_),
    .X(_04849_));
 sky130_fd_sc_hd__buf_6 _11680_ (.A(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__a211o_1 _11681_ (.A1(_04827_),
    .A2(_04837_),
    .B1(_04848_),
    .C1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__buf_6 _11682_ (.A(_04847_),
    .X(_04852_));
 sky130_fd_sc_hd__buf_4 _11683_ (.A(_04829_),
    .X(_04853_));
 sky130_fd_sc_hd__mux2_1 _11684_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04853_),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_4 _11686_ (.A(_04838_),
    .X(_04856_));
 sky130_fd_sc_hd__buf_4 _11687_ (.A(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_8 _11688_ (.A(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__mux2_1 _11689_ (.A0(_04854_),
    .A1(_04855_),
    .S(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__mux2_1 _11690_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04842_),
    .X(_04860_));
 sky130_fd_sc_hd__mux2_1 _11691_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_04853_),
    .X(_04861_));
 sky130_fd_sc_hd__buf_6 _11692_ (.A(_04772_),
    .X(_04862_));
 sky130_fd_sc_hd__nor2_4 _11693_ (.A(_04862_),
    .B(_04788_),
    .Y(_04863_));
 sky130_fd_sc_hd__buf_4 _11694_ (.A(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__buf_4 _11695_ (.A(_04770_),
    .X(_04865_));
 sky130_fd_sc_hd__a221o_1 _11696_ (.A1(_04807_),
    .A2(_04860_),
    .B1(_04861_),
    .B2(_04864_),
    .C1(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__a21o_1 _11697_ (.A1(_04852_),
    .A2(_04859_),
    .B1(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__buf_6 _11698_ (.A(_04770_),
    .X(_04868_));
 sky130_fd_sc_hd__mux2_1 _11699_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04832_),
    .X(_04869_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04832_),
    .X(_04870_));
 sky130_fd_sc_hd__mux2_1 _11701_ (.A0(_04869_),
    .A1(_04870_),
    .S(_04777_),
    .X(_04871_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04832_),
    .X(_04872_));
 sky130_fd_sc_hd__mux2_1 _11703_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04832_),
    .X(_04873_));
 sky130_fd_sc_hd__clkbuf_8 _11704_ (.A(_04788_),
    .X(_04874_));
 sky130_fd_sc_hd__mux2_1 _11705_ (.A0(_04872_),
    .A1(_04873_),
    .S(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(_04871_),
    .A1(_04875_),
    .S(_04827_),
    .X(_04876_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04842_),
    .X(_04877_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04829_),
    .X(_04878_));
 sky130_fd_sc_hd__or2_1 _11709_ (.A(_04844_),
    .B(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__o211a_1 _11710_ (.A1(_04841_),
    .A2(_04877_),
    .B1(_04879_),
    .C1(_04847_),
    .X(_04880_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04833_),
    .X(_04881_));
 sky130_fd_sc_hd__mux2_1 _11712_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04833_),
    .X(_04882_));
 sky130_fd_sc_hd__a221o_1 _11713_ (.A1(_04794_),
    .A2(_04881_),
    .B1(_04864_),
    .B2(_04882_),
    .C1(_04849_),
    .X(_04883_));
 sky130_fd_sc_hd__or2_2 _11714_ (.A(_04768_),
    .B(_04824_),
    .X(_04884_));
 sky130_fd_sc_hd__buf_6 _11715_ (.A(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__o221a_1 _11716_ (.A1(_04868_),
    .A2(_04876_),
    .B1(_04880_),
    .B2(_04883_),
    .C1(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__a31o_1 _11717_ (.A1(_04826_),
    .A2(_04851_),
    .A3(_04867_),
    .B1(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__buf_4 _11718_ (.A(_04853_),
    .X(_04888_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__buf_4 _11720_ (.A(_04844_),
    .X(_04890_));
 sky130_fd_sc_hd__mux2_1 _11721_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04853_),
    .X(_04891_));
 sky130_fd_sc_hd__or2_1 _11722_ (.A(_04890_),
    .B(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__o211a_1 _11723_ (.A1(_04841_),
    .A2(_04889_),
    .B1(_04892_),
    .C1(_04852_),
    .X(_04893_));
 sky130_fd_sc_hd__mux2_1 _11724_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04812_),
    .X(_04894_));
 sky130_fd_sc_hd__clkbuf_4 _11725_ (.A(_04842_),
    .X(_04895_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__a221o_1 _11727_ (.A1(_04807_),
    .A2(_04894_),
    .B1(_04896_),
    .B2(_04864_),
    .C1(_04850_),
    .X(_04897_));
 sky130_fd_sc_hd__nor2_4 _11728_ (.A(_04826_),
    .B(_04821_),
    .Y(_04898_));
 sky130_fd_sc_hd__mux2_1 _11729_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04842_),
    .X(_04899_));
 sky130_fd_sc_hd__or2_1 _11730_ (.A(_04890_),
    .B(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__mux2_1 _11731_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04853_),
    .X(_04901_));
 sky130_fd_sc_hd__o21a_1 _11732_ (.A1(_04841_),
    .A2(_04901_),
    .B1(_04847_),
    .X(_04902_));
 sky130_fd_sc_hd__mux2_1 _11733_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_04842_),
    .X(_04903_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04842_),
    .X(_04904_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(_04903_),
    .A1(_04904_),
    .S(_04858_),
    .X(_04905_));
 sky130_fd_sc_hd__a221o_1 _11736_ (.A1(_04900_),
    .A2(_04902_),
    .B1(_04905_),
    .B2(_04827_),
    .C1(_04868_),
    .X(_04906_));
 sky130_fd_sc_hd__o211a_1 _11737_ (.A1(_04893_),
    .A2(_04897_),
    .B1(_04898_),
    .C1(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__or2_4 _11738_ (.A(_04768_),
    .B(_04820_),
    .X(_04908_));
 sky130_fd_sc_hd__mux2_1 _11739_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04833_),
    .X(_04909_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04833_),
    .X(_04910_));
 sky130_fd_sc_hd__mux2_1 _11741_ (.A0(_04909_),
    .A1(_04910_),
    .S(_04836_),
    .X(_04911_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04830_),
    .X(_04912_));
 sky130_fd_sc_hd__mux2_1 _11743_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04832_),
    .X(_04913_));
 sky130_fd_sc_hd__or2_1 _11744_ (.A(_04844_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__o211a_1 _11745_ (.A1(_04841_),
    .A2(_04912_),
    .B1(_04914_),
    .C1(_04847_),
    .X(_04915_));
 sky130_fd_sc_hd__a211o_1 _11746_ (.A1(_04827_),
    .A2(_04911_),
    .B1(_04915_),
    .C1(_04850_),
    .X(_04916_));
 sky130_fd_sc_hd__mux2_1 _11747_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04842_),
    .X(_04917_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04842_),
    .X(_04918_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(_04917_),
    .A1(_04918_),
    .S(_04858_),
    .X(_04919_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04842_),
    .X(_04920_));
 sky130_fd_sc_hd__mux2_1 _11751_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04853_),
    .X(_04921_));
 sky130_fd_sc_hd__a221o_1 _11752_ (.A1(_04807_),
    .A2(_04920_),
    .B1(_04921_),
    .B2(_04864_),
    .C1(_04865_),
    .X(_04922_));
 sky130_fd_sc_hd__a21o_1 _11753_ (.A1(_04852_),
    .A2(_04919_),
    .B1(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__and4_1 _11754_ (.A(_04826_),
    .B(_04908_),
    .C(_04916_),
    .D(_04923_),
    .X(_04924_));
 sky130_fd_sc_hd__a211o_1 _11755_ (.A1(_04821_),
    .A2(_04887_),
    .B1(_04907_),
    .C1(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__a2bb2o_1 _11756_ (.A1_N(_04705_),
    .A2_N(_04817_),
    .B1(_04818_),
    .B2(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_8 _11757_ (.A(_04799_),
    .X(_04927_));
 sky130_fd_sc_hd__or3_1 _11758_ (.A(_04844_),
    .B(_04700_),
    .C(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__or4b_1 _11759_ (.A(_04825_),
    .B(_04821_),
    .C(_04928_),
    .D_N(_04790_),
    .X(_04929_));
 sky130_fd_sc_hd__inv_2 _11760_ (.A(\rbzero.row_render.size[2] ),
    .Y(_04930_));
 sky130_fd_sc_hd__nor2_1 _11761_ (.A(\rbzero.row_render.size[1] ),
    .B(\rbzero.row_render.size[0] ),
    .Y(_04931_));
 sky130_fd_sc_hd__nand2_1 _11762_ (.A(_04930_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__or2_1 _11763_ (.A(\rbzero.row_render.size[3] ),
    .B(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__or3_1 _11764_ (.A(\rbzero.row_render.size[5] ),
    .B(\rbzero.row_render.size[4] ),
    .C(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__and2_1 _11765_ (.A(\rbzero.row_render.size[6] ),
    .B(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__o21a_1 _11766_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_04935_),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04936_));
 sky130_fd_sc_hd__a21o_1 _11767_ (.A1(\rbzero.row_render.size[7] ),
    .A2(\rbzero.row_render.size[6] ),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_1 _11768_ (.A(\rbzero.row_render.size[9] ),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand3_1 _11769_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(\rbzero.row_render.size[6] ),
    .Y(_04939_));
 sky130_fd_sc_hd__and2_1 _11770_ (.A(_04937_),
    .B(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__xnor2_1 _11771_ (.A(\rbzero.row_render.size[7] ),
    .B(\rbzero.row_render.size[6] ),
    .Y(_04941_));
 sky130_fd_sc_hd__inv_2 _11772_ (.A(\rbzero.row_render.size[5] ),
    .Y(_04942_));
 sky130_fd_sc_hd__inv_2 _11773_ (.A(\rbzero.row_render.size[4] ),
    .Y(_04943_));
 sky130_fd_sc_hd__inv_2 _11774_ (.A(\rbzero.row_render.size[3] ),
    .Y(_04944_));
 sky130_fd_sc_hd__inv_2 _11775_ (.A(\rbzero.row_render.size[1] ),
    .Y(_04945_));
 sky130_fd_sc_hd__a211oi_1 _11776_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_04579_),
    .B1(_04576_),
    .C1(\rbzero.row_render.size[0] ),
    .Y(_04946_));
 sky130_fd_sc_hd__a221o_1 _11777_ (.A1(_04930_),
    .A2(\gpout0.hpos[2] ),
    .B1(_04584_),
    .B2(_04945_),
    .C1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__o221a_1 _11778_ (.A1(_04930_),
    .A2(\gpout0.hpos[2] ),
    .B1(_04453_),
    .B2(_04944_),
    .C1(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__a221o_1 _11779_ (.A1(_04944_),
    .A2(_04453_),
    .B1(\gpout0.hpos[4] ),
    .B2(_04943_),
    .C1(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__o221a_1 _11780_ (.A1(_04942_),
    .A2(\gpout0.hpos[5] ),
    .B1(_04483_),
    .B2(_04943_),
    .C1(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__a221o_1 _11781_ (.A1(\rbzero.row_render.size[6] ),
    .A2(\gpout0.hpos[6] ),
    .B1(_04451_),
    .B2(_04942_),
    .C1(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__o221a_1 _11782_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_04457_),
    .B1(_04941_),
    .B2(\gpout0.hpos[7] ),
    .C1(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__a221o_1 _11783_ (.A1(_04013_),
    .A2(_04941_),
    .B1(_04940_),
    .B2(_04016_),
    .C1(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__nand2_1 _11784_ (.A(\rbzero.row_render.size[9] ),
    .B(_04937_),
    .Y(_04954_));
 sky130_fd_sc_hd__a21o_1 _11785_ (.A1(\gpout0.hpos[9] ),
    .A2(_04954_),
    .B1(_04938_),
    .X(_04955_));
 sky130_fd_sc_hd__o211a_1 _11786_ (.A1(_04016_),
    .A2(_04940_),
    .B1(_04953_),
    .C1(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__nor3_1 _11787_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(_04935_),
    .Y(_04957_));
 sky130_fd_sc_hd__nor2_1 _11788_ (.A(_04936_),
    .B(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__xnor2_1 _11789_ (.A(\rbzero.row_render.size[7] ),
    .B(_04935_),
    .Y(_04959_));
 sky130_fd_sc_hd__nor2_1 _11790_ (.A(\rbzero.row_render.size[6] ),
    .B(_04934_),
    .Y(_04960_));
 sky130_fd_sc_hd__nor2_1 _11791_ (.A(_04935_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__o21ai_1 _11792_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_04933_),
    .B1(\rbzero.row_render.size[5] ),
    .Y(_04962_));
 sky130_fd_sc_hd__nand2_1 _11793_ (.A(_04934_),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__xnor2_1 _11794_ (.A(\rbzero.row_render.size[4] ),
    .B(_04933_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand2_1 _11795_ (.A(\rbzero.row_render.size[3] ),
    .B(_04932_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_1 _11796_ (.A(_04933_),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__or2_1 _11797_ (.A(_04930_),
    .B(_04931_),
    .X(_04967_));
 sky130_fd_sc_hd__nand2_1 _11798_ (.A(_04932_),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__or2_1 _11799_ (.A(\rbzero.row_render.size[0] ),
    .B(\gpout0.hpos[1] ),
    .X(_04969_));
 sky130_fd_sc_hd__a221o_1 _11800_ (.A1(\rbzero.row_render.size[2] ),
    .A2(\gpout0.hpos[2] ),
    .B1(\gpout0.hpos[1] ),
    .B2(\gpout0.hpos[0] ),
    .C1(_04931_),
    .X(_04970_));
 sky130_fd_sc_hd__a31o_1 _11801_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_04617_),
    .A3(_04969_),
    .B1(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__o221a_1 _11802_ (.A1(_04453_),
    .A2(_04966_),
    .B1(_04968_),
    .B2(\gpout0.hpos[2] ),
    .C1(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__a221o_1 _11803_ (.A1(_04453_),
    .A2(_04966_),
    .B1(_04964_),
    .B2(\gpout0.hpos[4] ),
    .C1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__o221a_1 _11804_ (.A1(\gpout0.hpos[4] ),
    .A2(_04964_),
    .B1(_04963_),
    .B2(\gpout0.hpos[5] ),
    .C1(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__a221o_1 _11805_ (.A1(_04451_),
    .A2(_04963_),
    .B1(_04961_),
    .B2(\gpout0.hpos[6] ),
    .C1(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__o221a_1 _11806_ (.A1(\gpout0.hpos[6] ),
    .A2(_04961_),
    .B1(_04959_),
    .B2(\gpout0.hpos[7] ),
    .C1(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__a221o_1 _11807_ (.A1(\gpout0.hpos[7] ),
    .A2(_04959_),
    .B1(_04958_),
    .B2(_04016_),
    .C1(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__xnor2_1 _11808_ (.A(\rbzero.row_render.size[9] ),
    .B(_04936_),
    .Y(_04978_));
 sky130_fd_sc_hd__o211a_1 _11809_ (.A1(_04016_),
    .A2(_04958_),
    .B1(_04977_),
    .C1(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__nor2_1 _11810_ (.A(\gpout0.hpos[9] ),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__a211o_1 _11811_ (.A1(\gpout0.hpos[9] ),
    .A2(_04938_),
    .B1(_04956_),
    .C1(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__or4b_4 _11812_ (.A(\rbzero.row_render.size[10] ),
    .B(\rbzero.row_render.size[9] ),
    .C(_04936_),
    .D_N(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__a21oi_1 _11813_ (.A1(_04929_),
    .A2(_04982_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04983_));
 sky130_fd_sc_hd__o211a_1 _11814_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_04788_),
    .B1(_04832_),
    .C1(\rbzero.floor_leak[0] ),
    .X(_04984_));
 sky130_fd_sc_hd__a221o_1 _11815_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_04786_),
    .B1(_04874_),
    .B2(\rbzero.floor_leak[1] ),
    .C1(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__o221a_1 _11816_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04783_),
    .B1(_04827_),
    .B2(\rbzero.floor_leak[2] ),
    .C1(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__a221o_1 _11817_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04849_),
    .B1(_04885_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__o221a_1 _11818_ (.A1(\rbzero.floor_leak[4] ),
    .A2(_04885_),
    .B1(_04908_),
    .B2(\rbzero.floor_leak[5] ),
    .C1(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__a211oi_4 _11819_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_04908_),
    .B1(_04983_),
    .C1(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(_04701_),
    .A1(_04926_),
    .S(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__xor2_1 _11821_ (.A(_04679_),
    .B(\rbzero.debug_overlay.playerY[2] ),
    .X(_04991_));
 sky130_fd_sc_hd__xor2_1 _11822_ (.A(_04678_),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .X(_04992_));
 sky130_fd_sc_hd__inv_2 _11823_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .Y(_04993_));
 sky130_fd_sc_hd__xnor2_1 _11824_ (.A(_04680_),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .Y(_04994_));
 sky130_fd_sc_hd__o221a_1 _11825_ (.A1(\gpout0.vpos[6] ),
    .A2(_04993_),
    .B1(\rbzero.debug_overlay.playerX[0] ),
    .B2(_04454_),
    .C1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__or3b_1 _11826_ (.A(_04991_),
    .B(_04992_),
    .C_N(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__inv_2 _11827_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .Y(_04997_));
 sky130_fd_sc_hd__inv_2 _11828_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .Y(_04998_));
 sky130_fd_sc_hd__inv_2 _11829_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .Y(_04999_));
 sky130_fd_sc_hd__inv_2 _11830_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .Y(_05000_));
 sky130_fd_sc_hd__clkinv_2 _11831_ (.A(\gpout0.vpos[7] ),
    .Y(_05001_));
 sky130_fd_sc_hd__inv_2 _11832_ (.A(\gpout0.hpos[5] ),
    .Y(_05002_));
 sky130_fd_sc_hd__clkbuf_4 _11833_ (.A(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__a22o_1 _11834_ (.A1(_05001_),
    .A2(\rbzero.debug_overlay.playerY[4] ),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .B2(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__a221o_1 _11835_ (.A1(\gpout0.vpos[6] ),
    .A2(_04993_),
    .B1(_05000_),
    .B2(_04451_),
    .C1(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__a221o_1 _11836_ (.A1(_04999_),
    .A2(_04457_),
    .B1(_04455_),
    .B2(\rbzero.debug_overlay.playerX[1] ),
    .C1(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__a221o_1 _11837_ (.A1(_04671_),
    .A2(_04997_),
    .B1(_04998_),
    .B2(_04483_),
    .C1(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__xor2_1 _11838_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_04013_),
    .X(_05008_));
 sky130_fd_sc_hd__a221o_1 _11839_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_04454_),
    .B1(_04481_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .C1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__or3_2 _11840_ (.A(_04996_),
    .B(_05007_),
    .C(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__and3_1 _11841_ (.A(_04677_),
    .B(_04689_),
    .C(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__clkinv_2 _11842_ (.A(_04679_),
    .Y(_05012_));
 sky130_fd_sc_hd__a22o_1 _11843_ (.A1(_05001_),
    .A2(\rbzero.map_overlay.i_mapdy[4] ),
    .B1(\rbzero.map_overlay.i_mapdy[2] ),
    .B2(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__inv_2 _11844_ (.A(\gpout0.vpos[6] ),
    .Y(_05014_));
 sky130_fd_sc_hd__inv_2 _11845_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .Y(_05015_));
 sky130_fd_sc_hd__clkbuf_4 _11846_ (.A(_04679_),
    .X(_05016_));
 sky130_fd_sc_hd__xor2_1 _11847_ (.A(_04680_),
    .B(\rbzero.map_overlay.i_mapdy[1] ),
    .X(_05017_));
 sky130_fd_sc_hd__a221o_1 _11848_ (.A1(_05014_),
    .A2(\rbzero.map_overlay.i_mapdy[3] ),
    .B1(_05015_),
    .B2(_05016_),
    .C1(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__inv_2 _11849_ (.A(\gpout0.vpos[3] ),
    .Y(_05019_));
 sky130_fd_sc_hd__or4_1 _11850_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_overlay.i_mapdy[2] ),
    .C(\rbzero.map_overlay.i_mapdy[1] ),
    .D(\rbzero.map_overlay.i_mapdy[0] ),
    .X(_05020_));
 sky130_fd_sc_hd__o21a_1 _11851_ (.A1(\rbzero.map_overlay.i_mapdy[5] ),
    .A2(_05020_),
    .B1(_05001_),
    .X(_05021_));
 sky130_fd_sc_hd__inv_2 _11852_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .Y(_05022_));
 sky130_fd_sc_hd__o22a_1 _11853_ (.A1(_05014_),
    .A2(\rbzero.map_overlay.i_mapdy[3] ),
    .B1(_05022_),
    .B2(_04678_),
    .X(_05023_));
 sky130_fd_sc_hd__o221a_1 _11854_ (.A1(_05019_),
    .A2(\rbzero.map_overlay.i_mapdy[0] ),
    .B1(_05021_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__or3b_1 _11855_ (.A(_05013_),
    .B(_05018_),
    .C_N(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__inv_2 _11856_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .Y(_05026_));
 sky130_fd_sc_hd__inv_2 _11857_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .Y(_05027_));
 sky130_fd_sc_hd__a22o_1 _11858_ (.A1(_05026_),
    .A2(_04013_),
    .B1(_04483_),
    .B2(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__xor2_1 _11859_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_04452_),
    .X(_05029_));
 sky130_fd_sc_hd__a22o_1 _11860_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04454_),
    .B1(_04455_),
    .B2(\rbzero.map_overlay.i_mapdx[1] ),
    .X(_05030_));
 sky130_fd_sc_hd__or4_1 _11861_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(\rbzero.map_overlay.i_mapdx[2] ),
    .C(\rbzero.map_overlay.i_mapdx[1] ),
    .D(\rbzero.map_overlay.i_mapdx[0] ),
    .X(_05031_));
 sky130_fd_sc_hd__o21a_1 _11862_ (.A1(\rbzero.map_overlay.i_mapdx[5] ),
    .A2(_05031_),
    .B1(_05026_),
    .X(_05032_));
 sky130_fd_sc_hd__xnor2_1 _11863_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_04457_),
    .Y(_05033_));
 sky130_fd_sc_hd__o221a_1 _11864_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04454_),
    .B1(_04013_),
    .B2(_05032_),
    .C1(_05033_),
    .X(_05034_));
 sky130_fd_sc_hd__or3b_1 _11865_ (.A(_05029_),
    .B(_05030_),
    .C_N(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__nor2_1 _11866_ (.A(_05028_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_1 _11867_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_04013_),
    .Y(_05037_));
 sky130_fd_sc_hd__or2_1 _11868_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_04013_),
    .X(_05038_));
 sky130_fd_sc_hd__inv_2 _11869_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .Y(_05039_));
 sky130_fd_sc_hd__xor2_1 _11870_ (.A(\gpout0.vpos[5] ),
    .B(\rbzero.map_overlay.i_othery[2] ),
    .X(_05040_));
 sky130_fd_sc_hd__a221o_1 _11871_ (.A1(\gpout0.vpos[7] ),
    .A2(_05039_),
    .B1(\rbzero.map_overlay.i_otherx[1] ),
    .B2(_04455_),
    .C1(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__xor2_1 _11872_ (.A(_04678_),
    .B(\rbzero.map_overlay.i_othery[0] ),
    .X(_05042_));
 sky130_fd_sc_hd__a211o_1 _11873_ (.A1(_05037_),
    .A2(_05038_),
    .B1(_05041_),
    .C1(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__inv_2 _11874_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .Y(_05044_));
 sky130_fd_sc_hd__xor2_1 _11875_ (.A(_04680_),
    .B(\rbzero.map_overlay.i_othery[1] ),
    .X(_05045_));
 sky130_fd_sc_hd__a221o_1 _11876_ (.A1(\rbzero.map_overlay.i_otherx[3] ),
    .A2(_04481_),
    .B1(_04451_),
    .B2(_05044_),
    .C1(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__inv_2 _11877_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .Y(_05047_));
 sky130_fd_sc_hd__xor2_1 _11878_ (.A(\gpout0.vpos[6] ),
    .B(\rbzero.map_overlay.i_othery[3] ),
    .X(_05048_));
 sky130_fd_sc_hd__a221o_1 _11879_ (.A1(_05001_),
    .A2(\rbzero.map_overlay.i_othery[4] ),
    .B1(_05047_),
    .B2(_04483_),
    .C1(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__inv_2 _11880_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .Y(_05050_));
 sky130_fd_sc_hd__xor2_1 _11881_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(_04453_),
    .X(_05051_));
 sky130_fd_sc_hd__a221o_1 _11882_ (.A1(_05050_),
    .A2(_04457_),
    .B1(_05003_),
    .B2(\rbzero.map_overlay.i_otherx[2] ),
    .C1(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__or4_1 _11883_ (.A(_05043_),
    .B(_05046_),
    .C(_05049_),
    .D(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__o21ai_1 _11884_ (.A1(_05025_),
    .A2(_05036_),
    .B1(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__inv_2 _11885_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .Y(_05055_));
 sky130_fd_sc_hd__inv_2 _11886_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .Y(_05056_));
 sky130_fd_sc_hd__a2bb2o_1 _11887_ (.A1_N(_04674_),
    .A2_N(\rbzero.debug_overlay.playerY[-2] ),
    .B1(_05056_),
    .B2(\gpout0.vpos[0] ),
    .X(_05057_));
 sky130_fd_sc_hd__a221o_1 _11888_ (.A1(_04674_),
    .A2(\rbzero.debug_overlay.playerY[-2] ),
    .B1(_05055_),
    .B2(_04584_),
    .C1(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__clkinv_2 _11889_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .Y(_05059_));
 sky130_fd_sc_hd__a2bb2o_1 _11890_ (.A1_N(\gpout0.vpos[0] ),
    .A2_N(_05056_),
    .B1(\rbzero.debug_overlay.playerX[-2] ),
    .B2(_04579_),
    .X(_05060_));
 sky130_fd_sc_hd__a221o_1 _11891_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_04615_),
    .B1(\gpout0.hpos[0] ),
    .B2(_05059_),
    .C1(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__inv_2 _11892_ (.A(\gpout0.vpos[2] ),
    .Y(_05062_));
 sky130_fd_sc_hd__o2bb2a_1 _11893_ (.A1_N(_05062_),
    .A2_N(\rbzero.debug_overlay.playerY[-1] ),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .B2(_04615_),
    .X(_05063_));
 sky130_fd_sc_hd__o221a_1 _11894_ (.A1(_05062_),
    .A2(\rbzero.debug_overlay.playerY[-1] ),
    .B1(_05059_),
    .B2(_04010_),
    .C1(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__or3b_1 _11895_ (.A(_05058_),
    .B(_05061_),
    .C_N(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__o21ai_1 _11896_ (.A1(_05010_),
    .A2(_05065_),
    .B1(_04699_),
    .Y(_05066_));
 sky130_fd_sc_hd__a21o_1 _11897_ (.A1(_05011_),
    .A2(_05054_),
    .B1(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__o21a_1 _11898_ (.A1(_04699_),
    .A2(_04990_),
    .B1(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__o22a_1 _11899_ (.A1(\rbzero.trace_state[0] ),
    .A2(_04686_),
    .B1(_04688_),
    .B2(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__nor2_1 _11900_ (.A(_04680_),
    .B(\gpout0.vpos[3] ),
    .Y(_05070_));
 sky130_fd_sc_hd__inv_2 _11901_ (.A(\gpout0.vpos[4] ),
    .Y(_05071_));
 sky130_fd_sc_hd__nor2_1 _11902_ (.A(_05071_),
    .B(_05019_),
    .Y(_05072_));
 sky130_fd_sc_hd__nor2_1 _11903_ (.A(_05070_),
    .B(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_2 _11904_ (.A(_05016_),
    .B(_04680_),
    .Y(_05074_));
 sky130_fd_sc_hd__inv_2 _11905_ (.A(_04677_),
    .Y(_05075_));
 sky130_fd_sc_hd__a311o_1 _11906_ (.A1(_04681_),
    .A2(_05073_),
    .A3(_05074_),
    .B1(_05075_),
    .C1(_04665_),
    .X(_05076_));
 sky130_fd_sc_hd__o21a_4 _11907_ (.A1(\gpout0.hpos[7] ),
    .A2(\gpout0.hpos[8] ),
    .B1(\gpout0.hpos[9] ),
    .X(_05077_));
 sky130_fd_sc_hd__and3_1 _11908_ (.A(\gpout0.vpos[7] ),
    .B(\gpout0.vpos[6] ),
    .C(_04679_),
    .X(_05078_));
 sky130_fd_sc_hd__a21o_4 _11909_ (.A1(\gpout0.vpos[8] ),
    .A2(_05078_),
    .B1(\gpout0.vpos[9] ),
    .X(_05079_));
 sky130_fd_sc_hd__a211oi_4 _11910_ (.A1(_04685_),
    .A2(_05076_),
    .B1(_05077_),
    .C1(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__o21a_4 _11911_ (.A1(_04685_),
    .A2(_05069_),
    .B1(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__buf_4 _11912_ (.A(net45),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_2 _11913_ (.A0(\reg_rgb[6] ),
    .A1(_05081_),
    .S(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__clkbuf_1 _11914_ (.A(_05083_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(\rbzero.color_sky[1] ),
    .A1(\rbzero.color_floor[1] ),
    .S(_04700_),
    .X(_05084_));
 sky130_fd_sc_hd__buf_6 _11916_ (.A(_04828_),
    .X(_05085_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__mux2_1 _11918_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_05085_),
    .X(_05087_));
 sky130_fd_sc_hd__mux2_1 _11919_ (.A0(_05086_),
    .A1(_05087_),
    .S(_04840_),
    .X(_05088_));
 sky130_fd_sc_hd__buf_6 _11920_ (.A(_04874_),
    .X(_05089_));
 sky130_fd_sc_hd__buf_4 _11921_ (.A(_04828_),
    .X(_05090_));
 sky130_fd_sc_hd__mux2_1 _11922_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__mux2_1 _11923_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_04828_),
    .X(_05092_));
 sky130_fd_sc_hd__or2_1 _11924_ (.A(_04835_),
    .B(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__o211a_1 _11925_ (.A1(_05089_),
    .A2(_05091_),
    .B1(_05093_),
    .C1(_04827_),
    .X(_05094_));
 sky130_fd_sc_hd__a211o_1 _11926_ (.A1(_04852_),
    .A2(_05088_),
    .B1(_05094_),
    .C1(_04849_),
    .X(_05095_));
 sky130_fd_sc_hd__mux2_1 _11927_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_05085_),
    .X(_05096_));
 sky130_fd_sc_hd__mux2_1 _11928_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_05085_),
    .X(_05097_));
 sky130_fd_sc_hd__mux2_1 _11929_ (.A0(_05096_),
    .A1(_05097_),
    .S(_04840_),
    .X(_05098_));
 sky130_fd_sc_hd__mux2_1 _11930_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_05090_),
    .X(_05099_));
 sky130_fd_sc_hd__mux2_1 _11931_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_04811_),
    .X(_05100_));
 sky130_fd_sc_hd__a22o_1 _11932_ (.A1(_04863_),
    .A2(_05099_),
    .B1(_05100_),
    .B2(_04794_),
    .X(_05101_));
 sky130_fd_sc_hd__a211o_1 _11933_ (.A1(_04847_),
    .A2(_05098_),
    .B1(_05101_),
    .C1(_04868_),
    .X(_05102_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04811_),
    .X(_05103_));
 sky130_fd_sc_hd__buf_4 _11935_ (.A(_04809_),
    .X(_05104_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__or2_1 _11937_ (.A(_04777_),
    .B(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__o211a_1 _11938_ (.A1(_05089_),
    .A2(_05103_),
    .B1(_05106_),
    .C1(_04847_),
    .X(_05107_));
 sky130_fd_sc_hd__mux2_1 _11939_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_05085_),
    .X(_05108_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_05090_),
    .X(_05109_));
 sky130_fd_sc_hd__a221o_1 _11941_ (.A1(_04794_),
    .A2(_05108_),
    .B1(_05109_),
    .B2(_04863_),
    .C1(_04770_),
    .X(_05110_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(_05104_),
    .X(_05111_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_05104_),
    .X(_05112_));
 sky130_fd_sc_hd__mux2_1 _11944_ (.A0(_05111_),
    .A1(_05112_),
    .S(_04835_),
    .X(_05113_));
 sky130_fd_sc_hd__mux2_1 _11945_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_04810_),
    .X(_05114_));
 sky130_fd_sc_hd__mux2_1 _11946_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_04809_),
    .X(_05115_));
 sky130_fd_sc_hd__or2_1 _11947_ (.A(_04776_),
    .B(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__o211a_1 _11948_ (.A1(_04874_),
    .A2(_05114_),
    .B1(_05116_),
    .C1(_04773_),
    .X(_05117_));
 sky130_fd_sc_hd__a211o_1 _11949_ (.A1(_04827_),
    .A2(_05113_),
    .B1(_05117_),
    .C1(_04849_),
    .X(_05118_));
 sky130_fd_sc_hd__o211a_1 _11950_ (.A1(_05107_),
    .A2(_05110_),
    .B1(_04885_),
    .C1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a31o_1 _11951_ (.A1(_04826_),
    .A2(_05095_),
    .A3(_05102_),
    .B1(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__buf_4 _11952_ (.A(_05085_),
    .X(_05121_));
 sky130_fd_sc_hd__clkbuf_4 _11953_ (.A(_04797_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_4 _11954_ (.A(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__or2_1 _11955_ (.A(\rbzero.tex_r1[26] ),
    .B(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__o211a_1 _11956_ (.A1(\rbzero.tex_r1[27] ),
    .A2(_05121_),
    .B1(_05124_),
    .C1(_04844_),
    .X(_05125_));
 sky130_fd_sc_hd__a31o_1 _11957_ (.A1(\rbzero.tex_r1[25] ),
    .A2(_04856_),
    .A3(_05123_),
    .B1(_04862_),
    .X(_05126_));
 sky130_fd_sc_hd__a31o_1 _11958_ (.A1(\rbzero.tex_r1[24] ),
    .A2(_04857_),
    .A3(_05121_),
    .B1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__or2_1 _11959_ (.A(\rbzero.tex_r1[30] ),
    .B(_05123_),
    .X(_05128_));
 sky130_fd_sc_hd__buf_4 _11960_ (.A(_04775_),
    .X(_05129_));
 sky130_fd_sc_hd__buf_4 _11961_ (.A(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__o211a_1 _11962_ (.A1(\rbzero.tex_r1[31] ),
    .A2(_05121_),
    .B1(_05128_),
    .C1(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__buf_4 _11963_ (.A(_04811_),
    .X(_05132_));
 sky130_fd_sc_hd__a31o_1 _11964_ (.A1(\rbzero.tex_r1[29] ),
    .A2(_04856_),
    .A3(_04799_),
    .B1(_04785_),
    .X(_05133_));
 sky130_fd_sc_hd__a31o_1 _11965_ (.A1(\rbzero.tex_r1[28] ),
    .A2(_04857_),
    .A3(_05132_),
    .B1(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__o221a_1 _11966_ (.A1(_05125_),
    .A2(_05127_),
    .B1(_05131_),
    .B2(_05134_),
    .C1(_04865_),
    .X(_05135_));
 sky130_fd_sc_hd__buf_4 _11967_ (.A(_05090_),
    .X(_05136_));
 sky130_fd_sc_hd__or2_1 _11968_ (.A(\rbzero.tex_r1[22] ),
    .B(_04799_),
    .X(_05137_));
 sky130_fd_sc_hd__o211a_1 _11969_ (.A1(\rbzero.tex_r1[23] ),
    .A2(_05136_),
    .B1(_05137_),
    .C1(_05130_),
    .X(_05138_));
 sky130_fd_sc_hd__buf_4 _11970_ (.A(_04839_),
    .X(_05139_));
 sky130_fd_sc_hd__a31o_1 _11971_ (.A1(\rbzero.tex_r1[21] ),
    .A2(_04856_),
    .A3(_04799_),
    .B1(_04786_),
    .X(_05140_));
 sky130_fd_sc_hd__a31o_1 _11972_ (.A1(\rbzero.tex_r1[20] ),
    .A2(_05139_),
    .A3(_05132_),
    .B1(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__or2_1 _11973_ (.A(\rbzero.tex_r1[18] ),
    .B(_04799_),
    .X(_05142_));
 sky130_fd_sc_hd__o211a_1 _11974_ (.A1(\rbzero.tex_r1[19] ),
    .A2(_05132_),
    .B1(_05142_),
    .C1(_05130_),
    .X(_05143_));
 sky130_fd_sc_hd__clkbuf_4 _11975_ (.A(_04797_),
    .X(_05144_));
 sky130_fd_sc_hd__buf_4 _11976_ (.A(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__a31o_1 _11977_ (.A1(\rbzero.tex_r1[17] ),
    .A2(_04856_),
    .A3(_05145_),
    .B1(_04862_),
    .X(_05146_));
 sky130_fd_sc_hd__a31o_1 _11978_ (.A1(\rbzero.tex_r1[16] ),
    .A2(_05139_),
    .A3(_04812_),
    .B1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__o221a_1 _11979_ (.A1(_05138_),
    .A2(_05141_),
    .B1(_05143_),
    .B2(_05147_),
    .C1(_04849_),
    .X(_05148_));
 sky130_fd_sc_hd__or4_1 _11980_ (.A(_04885_),
    .B(_04821_),
    .C(_05135_),
    .D(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__mux2_1 _11981_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_05121_),
    .X(_05150_));
 sky130_fd_sc_hd__mux2_1 _11982_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04853_),
    .X(_05151_));
 sky130_fd_sc_hd__mux2_1 _11983_ (.A0(_05150_),
    .A1(_05151_),
    .S(_04890_),
    .X(_05152_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[0] ),
    .S(_05121_),
    .X(_05153_));
 sky130_fd_sc_hd__mux2_1 _11985_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_05132_),
    .X(_05154_));
 sky130_fd_sc_hd__a221o_1 _11986_ (.A1(_04807_),
    .A2(_05153_),
    .B1(_05154_),
    .B2(_04864_),
    .C1(_04865_),
    .X(_05155_));
 sky130_fd_sc_hd__a21oi_1 _11987_ (.A1(_04852_),
    .A2(_05152_),
    .B1(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_05136_),
    .X(_05157_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_05121_),
    .X(_05158_));
 sky130_fd_sc_hd__mux2_1 _11990_ (.A0(_05157_),
    .A1(_05158_),
    .S(_04841_),
    .X(_05159_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_05136_),
    .X(_05160_));
 sky130_fd_sc_hd__mux2_1 _11992_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_05132_),
    .X(_05161_));
 sky130_fd_sc_hd__a221o_1 _11993_ (.A1(_04807_),
    .A2(_05160_),
    .B1(_05161_),
    .B2(_04864_),
    .C1(_04849_),
    .X(_05162_));
 sky130_fd_sc_hd__a21oi_1 _11994_ (.A1(_04852_),
    .A2(_05159_),
    .B1(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__o21ai_1 _11995_ (.A1(_05156_),
    .A2(_05163_),
    .B1(_04898_),
    .Y(_05164_));
 sky130_fd_sc_hd__o2111a_1 _11996_ (.A1(_04908_),
    .A2(_05120_),
    .B1(_05149_),
    .C1(_05164_),
    .D1(_04818_),
    .X(_05165_));
 sky130_fd_sc_hd__xnor2_1 _11997_ (.A(_04801_),
    .B(_04826_),
    .Y(_05166_));
 sky130_fd_sc_hd__a21boi_1 _11998_ (.A1(_04702_),
    .A2(_04805_),
    .B1_N(_04706_),
    .Y(_05167_));
 sky130_fd_sc_hd__a21oi_1 _11999_ (.A1(_04814_),
    .A2(_04792_),
    .B1(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__o211a_1 _12000_ (.A1(_04703_),
    .A2(_05166_),
    .B1(_05168_),
    .C1(_04704_),
    .X(_05169_));
 sky130_fd_sc_hd__or3b_1 _12001_ (.A(_05165_),
    .B(_05169_),
    .C_N(_04989_),
    .X(_05170_));
 sky130_fd_sc_hd__o21a_1 _12002_ (.A1(_04989_),
    .A2(_05084_),
    .B1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nor2_2 _12003_ (.A(_04481_),
    .B(_05002_),
    .Y(_05172_));
 sky130_fd_sc_hd__and3_1 _12004_ (.A(_04013_),
    .B(_05172_),
    .C(_04456_),
    .X(_05173_));
 sky130_fd_sc_hd__nand2_1 _12005_ (.A(_04679_),
    .B(_04451_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_1 _12006_ (.A(_05072_),
    .B(_05078_),
    .Y(_05175_));
 sky130_fd_sc_hd__o31ai_1 _12007_ (.A1(_04455_),
    .A2(_05073_),
    .A3(_05174_),
    .B1(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__nor2_1 _12008_ (.A(_05012_),
    .B(_05003_),
    .Y(_05177_));
 sky130_fd_sc_hd__nor2_1 _12009_ (.A(_04679_),
    .B(_04451_),
    .Y(_05178_));
 sky130_fd_sc_hd__o211a_1 _12010_ (.A1(_05177_),
    .A2(_05178_),
    .B1(_05019_),
    .C1(_04454_),
    .X(_05179_));
 sky130_fd_sc_hd__or3b_1 _12011_ (.A(_05176_),
    .B(_05179_),
    .C_N(_04697_),
    .X(_05180_));
 sky130_fd_sc_hd__a22o_1 _12012_ (.A1(_04678_),
    .A2(_04453_),
    .B1(_04455_),
    .B2(_05071_),
    .X(_05181_));
 sky130_fd_sc_hd__or3_1 _12013_ (.A(\gpout0.vpos[6] ),
    .B(_04457_),
    .C(_05178_),
    .X(_05182_));
 sky130_fd_sc_hd__a22o_1 _12014_ (.A1(_05019_),
    .A2(_04454_),
    .B1(_04483_),
    .B2(_04680_),
    .X(_05183_));
 sky130_fd_sc_hd__or4b_1 _12015_ (.A(_05181_),
    .B(_05182_),
    .C(_05183_),
    .D_N(_05174_),
    .X(_05184_));
 sky130_fd_sc_hd__or4bb_1 _12016_ (.A(_05173_),
    .B(_05180_),
    .C_N(_05184_),
    .D_N(_04693_),
    .X(_05185_));
 sky130_fd_sc_hd__clkbuf_4 _12017_ (.A(_04680_),
    .X(_05186_));
 sky130_fd_sc_hd__and4_1 _12018_ (.A(_05186_),
    .B(_04458_),
    .C(_04690_),
    .D(_05178_),
    .X(_05187_));
 sky130_fd_sc_hd__a22o_1 _12019_ (.A1(_04679_),
    .A2(_04482_),
    .B1(_04457_),
    .B2(_04680_),
    .X(_05188_));
 sky130_fd_sc_hd__xor2_1 _12020_ (.A(_04678_),
    .B(_04483_),
    .X(_05189_));
 sky130_fd_sc_hd__xor2_1 _12021_ (.A(\gpout0.vpos[6] ),
    .B(_04452_),
    .X(_05190_));
 sky130_fd_sc_hd__o22a_1 _12022_ (.A1(_04679_),
    .A2(_04453_),
    .B1(_04457_),
    .B2(_04680_),
    .X(_05191_));
 sky130_fd_sc_hd__and4b_1 _12023_ (.A_N(_05188_),
    .B(_05189_),
    .C(_05190_),
    .D(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__a41o_1 _12024_ (.A1(_04683_),
    .A2(_04093_),
    .A3(_04696_),
    .A4(_05187_),
    .B1(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__o21ai_1 _12025_ (.A1(_05028_),
    .A2(_05035_),
    .B1(_05053_),
    .Y(_05194_));
 sky130_fd_sc_hd__a31o_1 _12026_ (.A1(_05025_),
    .A2(_05185_),
    .A3(_05193_),
    .B1(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__a21o_1 _12027_ (.A1(_05011_),
    .A2(_05195_),
    .B1(_05066_),
    .X(_05196_));
 sky130_fd_sc_hd__o21a_1 _12028_ (.A1(_04699_),
    .A2(_05171_),
    .B1(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__o22a_1 _12029_ (.A1(_04472_),
    .A2(_04686_),
    .B1(_04688_),
    .B2(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__nor2_1 _12030_ (.A(_04453_),
    .B(_04665_),
    .Y(_05199_));
 sky130_fd_sc_hd__or2_2 _12031_ (.A(_04666_),
    .B(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__nor2_1 _12032_ (.A(\gpout0.hpos[7] ),
    .B(_04668_),
    .Y(_05201_));
 sky130_fd_sc_hd__or2_1 _12033_ (.A(_04669_),
    .B(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__nand2_2 _12034_ (.A(_04460_),
    .B(_04665_),
    .Y(_05203_));
 sky130_fd_sc_hd__xnor2_4 _12035_ (.A(_04481_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__or3_1 _12036_ (.A(\gpout0.hpos[6] ),
    .B(\gpout0.hpos[5] ),
    .C(_04667_),
    .X(_05205_));
 sky130_fd_sc_hd__inv_2 _12037_ (.A(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__o22a_1 _12038_ (.A1(\gpout0.hpos[4] ),
    .A2(_05200_),
    .B1(_05206_),
    .B2(_04668_),
    .X(_05207_));
 sky130_fd_sc_hd__and3b_1 _12039_ (.A_N(_05202_),
    .B(_05204_),
    .C(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__or3_1 _12040_ (.A(_04670_),
    .B(_05077_),
    .C(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__nor2_1 _12041_ (.A(_05200_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__and2_1 _12042_ (.A(_04455_),
    .B(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__or3_1 _12043_ (.A(_05172_),
    .B(_05201_),
    .C(_05207_),
    .X(_05212_));
 sky130_fd_sc_hd__and2b_1 _12044_ (.A_N(_04669_),
    .B(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__xnor2_1 _12045_ (.A(_04016_),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__clkinv_2 _12046_ (.A(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__mux2_1 _12047_ (.A0(_05215_),
    .A1(_04016_),
    .S(_05208_),
    .X(_05216_));
 sky130_fd_sc_hd__and2_1 _12048_ (.A(_05204_),
    .B(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__and3_2 _12049_ (.A(_04451_),
    .B(_05211_),
    .C(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__nor2_1 _12050_ (.A(_04666_),
    .B(_05199_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand2_1 _12051_ (.A(_04456_),
    .B(_04665_),
    .Y(_05220_));
 sky130_fd_sc_hd__nand2_1 _12052_ (.A(_04667_),
    .B(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__nor3_2 _12053_ (.A(_05219_),
    .B(_05221_),
    .C(_05209_),
    .Y(_05222_));
 sky130_fd_sc_hd__and3_2 _12054_ (.A(_04451_),
    .B(_05222_),
    .C(_05217_),
    .X(_05223_));
 sky130_fd_sc_hd__nand2_1 _12055_ (.A(_05003_),
    .B(_05220_),
    .Y(_05224_));
 sky130_fd_sc_hd__nand2_1 _12056_ (.A(_05203_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__and3_1 _12057_ (.A(_04483_),
    .B(_05225_),
    .C(_05210_),
    .X(_05226_));
 sky130_fd_sc_hd__inv_2 _12058_ (.A(_05204_),
    .Y(_05227_));
 sky130_fd_sc_hd__mux2_1 _12059_ (.A0(_05172_),
    .A1(_05227_),
    .S(_05207_),
    .X(_05228_));
 sky130_fd_sc_hd__xnor2_2 _12060_ (.A(_05202_),
    .B(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__or2_1 _12061_ (.A(_05229_),
    .B(_05214_),
    .X(_05230_));
 sky130_fd_sc_hd__nor2_1 _12062_ (.A(_05204_),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__and2_2 _12063_ (.A(_05226_),
    .B(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(_05204_),
    .B(_05214_),
    .X(_05233_));
 sky130_fd_sc_hd__and3b_2 _12065_ (.A_N(_05233_),
    .B(_05003_),
    .C(_05211_),
    .X(_05234_));
 sky130_fd_sc_hd__inv_2 _12066_ (.A(_05230_),
    .Y(_05235_));
 sky130_fd_sc_hd__and3_2 _12067_ (.A(_05172_),
    .B(_05211_),
    .C(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__a22o_1 _12068_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_05234_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.playerY[-9] ),
    .X(_05237_));
 sky130_fd_sc_hd__and2_1 _12069_ (.A(_05203_),
    .B(_05224_),
    .X(_05238_));
 sky130_fd_sc_hd__and3_1 _12070_ (.A(_04483_),
    .B(_05238_),
    .C(_05210_),
    .X(_05239_));
 sky130_fd_sc_hd__and3_2 _12071_ (.A(_05204_),
    .B(_05216_),
    .C(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__or3b_1 _12072_ (.A(_05219_),
    .B(_05209_),
    .C_N(_05221_),
    .X(_05241_));
 sky130_fd_sc_hd__or2_1 _12073_ (.A(_05238_),
    .B(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__nor2_4 _12074_ (.A(_05242_),
    .B(_05233_),
    .Y(_05243_));
 sky130_fd_sc_hd__and2_1 _12075_ (.A(_05229_),
    .B(_05239_),
    .X(_05244_));
 sky130_fd_sc_hd__a211o_1 _12076_ (.A1(\rbzero.debug_overlay.playerY[5] ),
    .A2(_05244_),
    .B1(_04681_),
    .C1(_05019_),
    .X(_05245_));
 sky130_fd_sc_hd__a221o_1 _12077_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_05240_),
    .B1(_05243_),
    .B2(\rbzero.debug_overlay.playerY[-4] ),
    .C1(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__a211o_1 _12078_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_05232_),
    .B1(_05237_),
    .C1(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__a221o_1 _12079_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_05218_),
    .B1(_05223_),
    .B2(\rbzero.debug_overlay.playerY[-2] ),
    .C1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__and3_1 _12080_ (.A(_05204_),
    .B(_05226_),
    .C(_05216_),
    .X(_05249_));
 sky130_fd_sc_hd__nor2_1 _12081_ (.A(_05225_),
    .B(_05241_),
    .Y(_05250_));
 sky130_fd_sc_hd__and2_1 _12082_ (.A(\gpout0.hpos[6] ),
    .B(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__and2_2 _12083_ (.A(_05251_),
    .B(_05235_),
    .X(_05252_));
 sky130_fd_sc_hd__and3_2 _12084_ (.A(_05204_),
    .B(_05250_),
    .C(_05216_),
    .X(_05253_));
 sky130_fd_sc_hd__a22o_1 _12085_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(_05252_),
    .B1(_05253_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .X(_05254_));
 sky130_fd_sc_hd__and3_1 _12086_ (.A(_05003_),
    .B(_05222_),
    .C(_05217_),
    .X(_05255_));
 sky130_fd_sc_hd__and3_1 _12087_ (.A(_05003_),
    .B(_05211_),
    .C(_05217_),
    .X(_05256_));
 sky130_fd_sc_hd__and3b_1 _12088_ (.A_N(_05242_),
    .B(_05204_),
    .C(_05216_),
    .X(_05257_));
 sky130_fd_sc_hd__and3_2 _12089_ (.A(_05003_),
    .B(_05222_),
    .C(_05231_),
    .X(_05258_));
 sky130_fd_sc_hd__a22o_1 _12090_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_05257_),
    .B1(_05258_),
    .B2(\rbzero.debug_overlay.playerY[-6] ),
    .X(_05259_));
 sky130_fd_sc_hd__a221o_1 _12091_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_05255_),
    .B1(_05256_),
    .B2(\rbzero.debug_overlay.playerY[3] ),
    .C1(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__a211o_1 _12092_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_05249_),
    .B1(_05254_),
    .C1(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__o22a_1 _12093_ (.A1(_04457_),
    .A2(_04451_),
    .B1(_05222_),
    .B2(_05251_),
    .X(_05262_));
 sky130_fd_sc_hd__a22o_1 _12094_ (.A1(_05172_),
    .A2(_05211_),
    .B1(_05226_),
    .B2(_05227_),
    .X(_05263_));
 sky130_fd_sc_hd__o31a_1 _12095_ (.A1(_05262_),
    .A2(_05263_),
    .A3(_05239_),
    .B1(_05229_),
    .X(_05264_));
 sky130_fd_sc_hd__or4_1 _12096_ (.A(_05249_),
    .B(_05257_),
    .C(_05255_),
    .D(_05256_),
    .X(_05265_));
 sky130_fd_sc_hd__or2_2 _12097_ (.A(_05264_),
    .B(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__a22o_1 _12098_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_05240_),
    .B1(_05253_),
    .B2(\rbzero.debug_overlay.facingX[0] ),
    .X(_05267_));
 sky130_fd_sc_hd__a21o_1 _12099_ (.A1(\rbzero.debug_overlay.facingX[-6] ),
    .A2(_05258_),
    .B1(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__a22o_1 _12100_ (.A1(\rbzero.debug_overlay.facingX[-7] ),
    .A2(_05232_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.facingX[-9] ),
    .X(_05269_));
 sky130_fd_sc_hd__a221o_1 _12101_ (.A1(\rbzero.debug_overlay.facingX[-8] ),
    .A2(_05252_),
    .B1(_05243_),
    .B2(\rbzero.debug_overlay.facingX[-4] ),
    .C1(_05071_),
    .X(_05270_));
 sky130_fd_sc_hd__a211o_1 _12102_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_05234_),
    .B1(_05269_),
    .C1(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__a221o_1 _12103_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(_05218_),
    .B1(_05223_),
    .B2(\rbzero.debug_overlay.facingX[-2] ),
    .C1(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__a211o_1 _12104_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_05266_),
    .B1(_05268_),
    .C1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__and3_1 _12105_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_05251_),
    .C(_05235_),
    .X(_05274_));
 sky130_fd_sc_hd__a221o_1 _12106_ (.A1(\rbzero.debug_overlay.facingY[-1] ),
    .A2(_05218_),
    .B1(_05223_),
    .B2(\rbzero.debug_overlay.facingY[-2] ),
    .C1(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__nand2_1 _12107_ (.A(_04679_),
    .B(_05070_),
    .Y(_05276_));
 sky130_fd_sc_hd__a221o_1 _12108_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_05234_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .C1(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__a221o_1 _12109_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_05253_),
    .B1(_05243_),
    .B2(\rbzero.debug_overlay.facingY[-4] ),
    .C1(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__a22o_1 _12110_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_05258_),
    .B1(_05232_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .X(_05279_));
 sky130_fd_sc_hd__a221o_1 _12111_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_05266_),
    .B1(_05240_),
    .B2(\rbzero.debug_overlay.facingY[-3] ),
    .C1(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__a22o_1 _12112_ (.A1(\rbzero.debug_overlay.vplaneY[-3] ),
    .A2(_05240_),
    .B1(_05252_),
    .B2(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_05281_));
 sky130_fd_sc_hd__clkbuf_4 _12113_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_05282_));
 sky130_fd_sc_hd__a22o_1 _12114_ (.A1(\rbzero.debug_overlay.vplaneY[-5] ),
    .A2(_05234_),
    .B1(_05243_),
    .B2(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_05283_));
 sky130_fd_sc_hd__a221o_1 _12115_ (.A1(\rbzero.debug_overlay.vplaneY[-7] ),
    .A2(_05232_),
    .B1(_05253_),
    .B2(\rbzero.debug_overlay.vplaneY[0] ),
    .C1(_05019_),
    .X(_05284_));
 sky130_fd_sc_hd__a211o_1 _12116_ (.A1(_05282_),
    .A2(_05236_),
    .B1(_05283_),
    .C1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__a221o_1 _12117_ (.A1(\rbzero.debug_overlay.vplaneY[-1] ),
    .A2(_05218_),
    .B1(_05223_),
    .B2(\rbzero.debug_overlay.vplaneY[-2] ),
    .C1(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__a211o_1 _12118_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(_05258_),
    .B1(_05281_),
    .C1(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__a21oi_1 _12119_ (.A1(\rbzero.debug_overlay.vplaneY[10] ),
    .A2(_05266_),
    .B1(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__a22o_1 _12120_ (.A1(\rbzero.debug_overlay.vplaneX[-3] ),
    .A2(_05240_),
    .B1(_05253_),
    .B2(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_05289_));
 sky130_fd_sc_hd__clkbuf_4 _12121_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_4 _12122_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_4 _12123_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_05292_));
 sky130_fd_sc_hd__a22o_1 _12124_ (.A1(_05291_),
    .A2(_05234_),
    .B1(_05243_),
    .B2(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__a221o_1 _12125_ (.A1(\rbzero.debug_overlay.vplaneX[-8] ),
    .A2(_05252_),
    .B1(_05232_),
    .B2(\rbzero.debug_overlay.vplaneX[-7] ),
    .C1(\gpout0.vpos[3] ),
    .X(_05294_));
 sky130_fd_sc_hd__a211o_1 _12126_ (.A1(_05290_),
    .A2(_05236_),
    .B1(_05293_),
    .C1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__a221o_1 _12127_ (.A1(\rbzero.debug_overlay.vplaneX[-1] ),
    .A2(_05218_),
    .B1(_05223_),
    .B2(\rbzero.debug_overlay.vplaneX[-2] ),
    .C1(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__a211o_1 _12128_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(_05258_),
    .B1(_05289_),
    .C1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__a21oi_1 _12129_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_05266_),
    .B1(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__o31ai_1 _12130_ (.A1(_05074_),
    .A2(_05288_),
    .A3(_05298_),
    .B1(_05276_),
    .Y(_05299_));
 sky130_fd_sc_hd__o31a_1 _12131_ (.A1(_05275_),
    .A2(_05278_),
    .A3(_05280_),
    .B1(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__a31o_1 _12132_ (.A1(_05012_),
    .A2(_04678_),
    .A3(_05273_),
    .B1(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__o21ai_1 _12133_ (.A1(_05248_),
    .A2(_05261_),
    .B1(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__a22o_1 _12134_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(_05252_),
    .B1(_05232_),
    .B2(\rbzero.debug_overlay.playerX[-7] ),
    .X(_05303_));
 sky130_fd_sc_hd__a221o_1 _12135_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_05258_),
    .B1(_05218_),
    .B2(\rbzero.debug_overlay.playerX[-1] ),
    .C1(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__a221o_1 _12136_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_05244_),
    .B1(_05236_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_04682_),
    .X(_05305_));
 sky130_fd_sc_hd__a221o_1 _12137_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_05234_),
    .B1(_05243_),
    .B2(\rbzero.debug_overlay.playerX[-4] ),
    .C1(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__a22o_1 _12138_ (.A1(\rbzero.debug_overlay.playerX[-3] ),
    .A2(_05240_),
    .B1(_05253_),
    .B2(\rbzero.debug_overlay.playerX[0] ),
    .X(_05307_));
 sky130_fd_sc_hd__a221o_1 _12139_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_05249_),
    .B1(_05255_),
    .B2(\rbzero.debug_overlay.playerX[2] ),
    .C1(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__a221o_1 _12140_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_05257_),
    .B1(_05256_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .C1(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__a211o_1 _12141_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_05223_),
    .B1(_05306_),
    .C1(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__o2bb2a_1 _12142_ (.A1_N(_04682_),
    .A2_N(_05302_),
    .B1(_05304_),
    .B2(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__or3b_1 _12143_ (.A(_04665_),
    .B(_05075_),
    .C_N(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__or3b_1 _12144_ (.A(_04458_),
    .B(_05003_),
    .C_N(_04690_),
    .X(_05313_));
 sky130_fd_sc_hd__o31a_1 _12145_ (.A1(_04461_),
    .A2(_05200_),
    .A3(_05313_),
    .B1(_04685_),
    .X(_05314_));
 sky130_fd_sc_hd__a211oi_4 _12146_ (.A1(_05312_),
    .A2(_05314_),
    .B1(_05077_),
    .C1(_05079_),
    .Y(_05315_));
 sky130_fd_sc_hd__o21ai_1 _12147_ (.A1(_04685_),
    .A2(_05198_),
    .B1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__inv_2 _12148_ (.A(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__mux2_2 _12149_ (.A0(\reg_rgb[7] ),
    .A1(_05317_),
    .S(_05082_),
    .X(_05318_));
 sky130_fd_sc_hd__clkbuf_1 _12150_ (.A(_05318_),
    .X(net71));
 sky130_fd_sc_hd__or3_2 _12151_ (.A(_04694_),
    .B(_04695_),
    .C(_04698_),
    .X(_05319_));
 sky130_fd_sc_hd__o21ba_1 _12152_ (.A1(_05319_),
    .A2(_05010_),
    .B1_N(_04688_),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _12153_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_04700_),
    .X(_05321_));
 sky130_fd_sc_hd__inv_2 _12154_ (.A(_04705_),
    .Y(_05322_));
 sky130_fd_sc_hd__and3_1 _12155_ (.A(_04847_),
    .B(_04836_),
    .C(_04927_),
    .X(_05323_));
 sky130_fd_sc_hd__a31oi_1 _12156_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04807_),
    .A3(_04813_),
    .B1(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__o21ai_1 _12157_ (.A1(_04804_),
    .A2(_05324_),
    .B1(_04702_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_1 _12158_ (.A(_04702_),
    .B(\rbzero.row_render.wall[0] ),
    .Y(_05326_));
 sky130_fd_sc_hd__o21ai_1 _12159_ (.A1(_04781_),
    .A2(_05326_),
    .B1(_04703_),
    .Y(_05327_));
 sky130_fd_sc_hd__a31o_1 _12160_ (.A1(_04706_),
    .A2(_04806_),
    .A3(_05325_),
    .B1(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04829_),
    .X(_05329_));
 sky130_fd_sc_hd__mux2_1 _12162_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04828_),
    .X(_05330_));
 sky130_fd_sc_hd__or2_1 _12163_ (.A(_05129_),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__buf_6 _12164_ (.A(_04862_),
    .X(_05332_));
 sky130_fd_sc_hd__o211a_1 _12165_ (.A1(_04840_),
    .A2(_05329_),
    .B1(_05331_),
    .C1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__mux2_1 _12166_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04829_),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04828_),
    .X(_05335_));
 sky130_fd_sc_hd__or2_1 _12168_ (.A(_04839_),
    .B(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__o211a_1 _12169_ (.A1(_05130_),
    .A2(_05334_),
    .B1(_05336_),
    .C1(_04827_),
    .X(_05337_));
 sky130_fd_sc_hd__mux2_1 _12170_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04811_),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_05104_),
    .X(_05339_));
 sky130_fd_sc_hd__or2_1 _12172_ (.A(_04777_),
    .B(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__o211a_1 _12173_ (.A1(_05089_),
    .A2(_05338_),
    .B1(_05340_),
    .C1(_04847_),
    .X(_05341_));
 sky130_fd_sc_hd__mux2_1 _12174_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_05085_),
    .X(_05342_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_05090_),
    .X(_05343_));
 sky130_fd_sc_hd__a221o_1 _12176_ (.A1(_04863_),
    .A2(_05342_),
    .B1(_05343_),
    .B2(_04794_),
    .C1(_04783_),
    .X(_05344_));
 sky130_fd_sc_hd__o32a_1 _12177_ (.A1(_04865_),
    .A2(_05333_),
    .A3(_05337_),
    .B1(_05341_),
    .B2(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__mux2_1 _12178_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_05104_),
    .X(_05346_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_05104_),
    .X(_05347_));
 sky130_fd_sc_hd__mux2_1 _12180_ (.A0(_05346_),
    .A1(_05347_),
    .S(_04835_),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_05104_),
    .X(_05349_));
 sky130_fd_sc_hd__mux2_1 _12182_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04809_),
    .X(_05350_));
 sky130_fd_sc_hd__or2_1 _12183_ (.A(_04776_),
    .B(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__o211a_1 _12184_ (.A1(_04874_),
    .A2(_05349_),
    .B1(_05351_),
    .C1(_04773_),
    .X(_05352_));
 sky130_fd_sc_hd__a211o_1 _12185_ (.A1(_04827_),
    .A2(_05348_),
    .B1(_05352_),
    .C1(_04783_),
    .X(_05353_));
 sky130_fd_sc_hd__mux2_1 _12186_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04810_),
    .X(_05354_));
 sky130_fd_sc_hd__mux2_1 _12187_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_04810_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _12188_ (.A0(_05354_),
    .A1(_05355_),
    .S(_04874_),
    .X(_05356_));
 sky130_fd_sc_hd__mux2_1 _12189_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04810_),
    .X(_05357_));
 sky130_fd_sc_hd__mux2_1 _12190_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_04832_),
    .X(_05358_));
 sky130_fd_sc_hd__a221o_1 _12191_ (.A1(_04794_),
    .A2(_05357_),
    .B1(_05358_),
    .B2(_04863_),
    .C1(_04770_),
    .X(_05359_));
 sky130_fd_sc_hd__a21o_1 _12192_ (.A1(_04847_),
    .A2(_05356_),
    .B1(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__a21o_1 _12193_ (.A1(_05353_),
    .A2(_05360_),
    .B1(_04885_),
    .X(_05361_));
 sky130_fd_sc_hd__o211a_1 _12194_ (.A1(_04826_),
    .A2(_05345_),
    .B1(_05361_),
    .C1(_04821_),
    .X(_05362_));
 sky130_fd_sc_hd__mux2_1 _12195_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_05121_),
    .X(_05363_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_05132_),
    .X(_05364_));
 sky130_fd_sc_hd__mux2_1 _12197_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_05085_),
    .X(_05365_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04828_),
    .X(_05366_));
 sky130_fd_sc_hd__or2_1 _12199_ (.A(_04835_),
    .B(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__o211a_1 _12200_ (.A1(_05089_),
    .A2(_05365_),
    .B1(_05367_),
    .C1(_05332_),
    .X(_05368_));
 sky130_fd_sc_hd__a221o_1 _12201_ (.A1(_04807_),
    .A2(_05363_),
    .B1(_05364_),
    .B2(_04864_),
    .C1(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__buf_4 _12202_ (.A(_04832_),
    .X(_05370_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _12204_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_05370_),
    .X(_05372_));
 sky130_fd_sc_hd__mux2_1 _12205_ (.A0(_05371_),
    .A1(_05372_),
    .S(_05089_),
    .X(_05373_));
 sky130_fd_sc_hd__mux2_1 _12206_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04811_),
    .X(_05374_));
 sky130_fd_sc_hd__mux2_1 _12207_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_05370_),
    .X(_05375_));
 sky130_fd_sc_hd__a221o_1 _12208_ (.A1(_04794_),
    .A2(_05374_),
    .B1(_05375_),
    .B2(_04864_),
    .C1(_04783_),
    .X(_05376_));
 sky130_fd_sc_hd__a21o_1 _12209_ (.A1(_04852_),
    .A2(_05373_),
    .B1(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__o211a_1 _12210_ (.A1(_04868_),
    .A2(_05369_),
    .B1(_05377_),
    .C1(_04898_),
    .X(_05378_));
 sky130_fd_sc_hd__mux2_1 _12211_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_05136_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _12212_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_04812_),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_05090_),
    .X(_05381_));
 sky130_fd_sc_hd__mux2_1 _12214_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04828_),
    .X(_05382_));
 sky130_fd_sc_hd__or2_1 _12215_ (.A(_04835_),
    .B(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__o211a_1 _12216_ (.A1(_05089_),
    .A2(_05381_),
    .B1(_05383_),
    .C1(_05332_),
    .X(_05384_));
 sky130_fd_sc_hd__a221o_1 _12217_ (.A1(_04807_),
    .A2(_05379_),
    .B1(_05380_),
    .B2(_04864_),
    .C1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__mux2_1 _12218_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_05370_),
    .X(_05386_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_05370_),
    .X(_05387_));
 sky130_fd_sc_hd__mux2_1 _12220_ (.A0(_05386_),
    .A1(_05387_),
    .S(_05089_),
    .X(_05388_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_05370_),
    .X(_05389_));
 sky130_fd_sc_hd__mux2_1 _12222_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_05370_),
    .X(_05390_));
 sky130_fd_sc_hd__a221o_1 _12223_ (.A1(_04794_),
    .A2(_05389_),
    .B1(_05390_),
    .B2(_04864_),
    .C1(_04770_),
    .X(_05391_));
 sky130_fd_sc_hd__a21o_1 _12224_ (.A1(_04852_),
    .A2(_05388_),
    .B1(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__o2111a_1 _12225_ (.A1(_04850_),
    .A2(_05385_),
    .B1(_05392_),
    .C1(_04908_),
    .D1(_04826_),
    .X(_05393_));
 sky130_fd_sc_hd__o31a_1 _12226_ (.A1(_05362_),
    .A2(_05378_),
    .A3(_05393_),
    .B1(_04818_),
    .X(_05394_));
 sky130_fd_sc_hd__a21o_1 _12227_ (.A1(_05322_),
    .A2(_05328_),
    .B1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__mux2_1 _12228_ (.A0(_05321_),
    .A1(_05395_),
    .S(_04989_),
    .X(_05396_));
 sky130_fd_sc_hd__nand2_1 _12229_ (.A(_05319_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__o2bb2a_1 _12230_ (.A1_N(_05320_),
    .A2_N(_05397_),
    .B1(_04686_),
    .B2(\rbzero.trace_state[2] ),
    .X(_05398_));
 sky130_fd_sc_hd__o21a_4 _12231_ (.A1(_04685_),
    .A2(_05398_),
    .B1(_05080_),
    .X(_05399_));
 sky130_fd_sc_hd__mux2_2 _12232_ (.A0(\reg_rgb[14] ),
    .A1(_05399_),
    .S(_05082_),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_1 _12233_ (.A(_05400_),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_04700_),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_4 _12235_ (.A(_05121_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_4 _12236_ (.A(_05123_),
    .X(_05403_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(\rbzero.tex_g1[62] ),
    .B(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__o211a_1 _12238_ (.A1(\rbzero.tex_g1[63] ),
    .A2(_05402_),
    .B1(_05404_),
    .C1(_04890_),
    .X(_05405_));
 sky130_fd_sc_hd__clkbuf_4 _12239_ (.A(_04856_),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_4 _12240_ (.A(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_4 _12241_ (.A(_05144_),
    .X(_05408_));
 sky130_fd_sc_hd__buf_6 _12242_ (.A(_04785_),
    .X(_05409_));
 sky130_fd_sc_hd__a31o_1 _12243_ (.A1(\rbzero.tex_g1[61] ),
    .A2(_05406_),
    .A3(_05408_),
    .B1(_05409_),
    .X(_05410_));
 sky130_fd_sc_hd__a31o_1 _12244_ (.A1(\rbzero.tex_g1[60] ),
    .A2(_05407_),
    .A3(_05402_),
    .B1(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__or2_1 _12245_ (.A(\rbzero.tex_g1[58] ),
    .B(_05408_),
    .X(_05412_));
 sky130_fd_sc_hd__o211a_1 _12246_ (.A1(\rbzero.tex_g1[59] ),
    .A2(_05402_),
    .B1(_05412_),
    .C1(_04890_),
    .X(_05413_));
 sky130_fd_sc_hd__a31o_1 _12247_ (.A1(\rbzero.tex_g1[57] ),
    .A2(_04857_),
    .A3(_05408_),
    .B1(_05332_),
    .X(_05414_));
 sky130_fd_sc_hd__a31o_1 _12248_ (.A1(\rbzero.tex_g1[56] ),
    .A2(_04858_),
    .A3(_05402_),
    .B1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__o221a_1 _12249_ (.A1(_05405_),
    .A2(_05411_),
    .B1(_05413_),
    .B2(_05415_),
    .C1(_04868_),
    .X(_05416_));
 sky130_fd_sc_hd__or2_1 _12250_ (.A(\rbzero.tex_g1[54] ),
    .B(_05408_),
    .X(_05417_));
 sky130_fd_sc_hd__o211a_1 _12251_ (.A1(\rbzero.tex_g1[55] ),
    .A2(_05402_),
    .B1(_05417_),
    .C1(_04890_),
    .X(_05418_));
 sky130_fd_sc_hd__a31o_1 _12252_ (.A1(\rbzero.tex_g1[53] ),
    .A2(_04857_),
    .A3(_05408_),
    .B1(_05409_),
    .X(_05419_));
 sky130_fd_sc_hd__a31o_1 _12253_ (.A1(\rbzero.tex_g1[52] ),
    .A2(_04858_),
    .A3(_05402_),
    .B1(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__or2_1 _12254_ (.A(\rbzero.tex_g1[50] ),
    .B(_05408_),
    .X(_05421_));
 sky130_fd_sc_hd__o211a_1 _12255_ (.A1(\rbzero.tex_g1[51] ),
    .A2(_05402_),
    .B1(_05421_),
    .C1(_04890_),
    .X(_05422_));
 sky130_fd_sc_hd__a31o_1 _12256_ (.A1(\rbzero.tex_g1[49] ),
    .A2(_04857_),
    .A3(_05408_),
    .B1(_05332_),
    .X(_05423_));
 sky130_fd_sc_hd__a31o_1 _12257_ (.A1(\rbzero.tex_g1[48] ),
    .A2(_04858_),
    .A3(_04813_),
    .B1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__o221a_1 _12258_ (.A1(_05418_),
    .A2(_05420_),
    .B1(_05422_),
    .B2(_05424_),
    .C1(_04850_),
    .X(_05425_));
 sky130_fd_sc_hd__or2_1 _12259_ (.A(\rbzero.tex_g1[38] ),
    .B(_05145_),
    .X(_05426_));
 sky130_fd_sc_hd__o211a_1 _12260_ (.A1(\rbzero.tex_g1[39] ),
    .A2(_04812_),
    .B1(_05426_),
    .C1(_04836_),
    .X(_05427_));
 sky130_fd_sc_hd__a31o_1 _12261_ (.A1(\rbzero.tex_g1[37] ),
    .A2(_04840_),
    .A3(_04927_),
    .B1(_04827_),
    .X(_05428_));
 sky130_fd_sc_hd__a311o_1 _12262_ (.A1(\rbzero.tex_g1[36] ),
    .A2(_04841_),
    .A3(_04813_),
    .B1(_05427_),
    .C1(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__or2_1 _12263_ (.A(\rbzero.tex_g1[34] ),
    .B(_04799_),
    .X(_05430_));
 sky130_fd_sc_hd__o211a_1 _12264_ (.A1(\rbzero.tex_g1[35] ),
    .A2(_04812_),
    .B1(_05430_),
    .C1(_04836_),
    .X(_05431_));
 sky130_fd_sc_hd__a31o_1 _12265_ (.A1(\rbzero.tex_g1[33] ),
    .A2(_04840_),
    .A3(_04927_),
    .B1(_05332_),
    .X(_05432_));
 sky130_fd_sc_hd__a311o_1 _12266_ (.A1(\rbzero.tex_g1[32] ),
    .A2(_04841_),
    .A3(_04813_),
    .B1(_05431_),
    .C1(_05432_),
    .X(_05433_));
 sky130_fd_sc_hd__or2_1 _12267_ (.A(\rbzero.tex_g1[46] ),
    .B(_04798_),
    .X(_05434_));
 sky130_fd_sc_hd__o211a_1 _12268_ (.A1(\rbzero.tex_g1[47] ),
    .A2(_04811_),
    .B1(_05434_),
    .C1(_04835_),
    .X(_05435_));
 sky130_fd_sc_hd__a31o_1 _12269_ (.A1(\rbzero.tex_g1[45] ),
    .A2(_04839_),
    .A3(_05145_),
    .B1(_04786_),
    .X(_05436_));
 sky130_fd_sc_hd__a311o_1 _12270_ (.A1(\rbzero.tex_g1[44] ),
    .A2(_04840_),
    .A3(_04812_),
    .B1(_05435_),
    .C1(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__or2_1 _12271_ (.A(\rbzero.tex_g1[42] ),
    .B(_04798_),
    .X(_05438_));
 sky130_fd_sc_hd__o211a_1 _12272_ (.A1(\rbzero.tex_g1[43] ),
    .A2(_04811_),
    .B1(_05438_),
    .C1(_04835_),
    .X(_05439_));
 sky130_fd_sc_hd__a31o_1 _12273_ (.A1(\rbzero.tex_g1[41] ),
    .A2(_04839_),
    .A3(_05145_),
    .B1(_04862_),
    .X(_05440_));
 sky130_fd_sc_hd__a311o_1 _12274_ (.A1(\rbzero.tex_g1[40] ),
    .A2(_04840_),
    .A3(_04812_),
    .B1(_05439_),
    .C1(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__a31o_1 _12275_ (.A1(_04865_),
    .A2(_05437_),
    .A3(_05441_),
    .B1(_04826_),
    .X(_05442_));
 sky130_fd_sc_hd__a31o_1 _12276_ (.A1(_04850_),
    .A2(_05429_),
    .A3(_05433_),
    .B1(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__o311a_1 _12277_ (.A1(_04885_),
    .A2(_05416_),
    .A3(_05425_),
    .B1(_04821_),
    .C1(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__or2_1 _12278_ (.A(\rbzero.tex_g1[6] ),
    .B(_04799_),
    .X(_05445_));
 sky130_fd_sc_hd__o211a_1 _12279_ (.A1(\rbzero.tex_g1[7] ),
    .A2(_05136_),
    .B1(_05445_),
    .C1(_05130_),
    .X(_05446_));
 sky130_fd_sc_hd__a31o_1 _12280_ (.A1(\rbzero.tex_g1[5] ),
    .A2(_05139_),
    .A3(_04927_),
    .B1(_05409_),
    .X(_05447_));
 sky130_fd_sc_hd__a311o_1 _12281_ (.A1(\rbzero.tex_g1[4] ),
    .A2(_04841_),
    .A3(_04813_),
    .B1(_05446_),
    .C1(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__or2_1 _12282_ (.A(\rbzero.tex_g1[2] ),
    .B(_05123_),
    .X(_05449_));
 sky130_fd_sc_hd__o211a_1 _12283_ (.A1(\rbzero.tex_g1[3] ),
    .A2(_05136_),
    .B1(_05449_),
    .C1(_05130_),
    .X(_05450_));
 sky130_fd_sc_hd__a31o_1 _12284_ (.A1(\rbzero.tex_g1[1] ),
    .A2(_05139_),
    .A3(_04927_),
    .B1(_05332_),
    .X(_05451_));
 sky130_fd_sc_hd__a311o_1 _12285_ (.A1(\rbzero.tex_g1[0] ),
    .A2(_04858_),
    .A3(_04813_),
    .B1(_05450_),
    .C1(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__or2_1 _12286_ (.A(\rbzero.tex_g1[14] ),
    .B(_04798_),
    .X(_05453_));
 sky130_fd_sc_hd__o211a_1 _12287_ (.A1(\rbzero.tex_g1[15] ),
    .A2(_05090_),
    .B1(_05453_),
    .C1(_05129_),
    .X(_05454_));
 sky130_fd_sc_hd__a31o_1 _12288_ (.A1(\rbzero.tex_g1[13] ),
    .A2(_04839_),
    .A3(_05145_),
    .B1(_04786_),
    .X(_05455_));
 sky130_fd_sc_hd__a311o_1 _12289_ (.A1(\rbzero.tex_g1[12] ),
    .A2(_05139_),
    .A3(_05132_),
    .B1(_05454_),
    .C1(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__or2_1 _12290_ (.A(\rbzero.tex_g1[10] ),
    .B(_04798_),
    .X(_05457_));
 sky130_fd_sc_hd__o211a_1 _12291_ (.A1(\rbzero.tex_g1[11] ),
    .A2(_05090_),
    .B1(_05457_),
    .C1(_05129_),
    .X(_05458_));
 sky130_fd_sc_hd__a31o_1 _12292_ (.A1(\rbzero.tex_g1[9] ),
    .A2(_04839_),
    .A3(_05145_),
    .B1(_04862_),
    .X(_05459_));
 sky130_fd_sc_hd__a311o_1 _12293_ (.A1(\rbzero.tex_g1[8] ),
    .A2(_04857_),
    .A3(_05132_),
    .B1(_05458_),
    .C1(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__a31o_1 _12294_ (.A1(_04865_),
    .A2(_05456_),
    .A3(_05460_),
    .B1(_04825_),
    .X(_05461_));
 sky130_fd_sc_hd__a31o_1 _12295_ (.A1(_04850_),
    .A2(_05448_),
    .A3(_05452_),
    .B1(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__or2_1 _12296_ (.A(\rbzero.tex_g1[22] ),
    .B(_05123_),
    .X(_05463_));
 sky130_fd_sc_hd__o211a_1 _12297_ (.A1(\rbzero.tex_g1[23] ),
    .A2(_05136_),
    .B1(_05463_),
    .C1(_05130_),
    .X(_05464_));
 sky130_fd_sc_hd__a31o_1 _12298_ (.A1(\rbzero.tex_g1[21] ),
    .A2(_05139_),
    .A3(_04927_),
    .B1(_05409_),
    .X(_05465_));
 sky130_fd_sc_hd__a311o_1 _12299_ (.A1(\rbzero.tex_g1[20] ),
    .A2(_04841_),
    .A3(_04813_),
    .B1(_05464_),
    .C1(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__or2_1 _12300_ (.A(\rbzero.tex_g1[18] ),
    .B(_05123_),
    .X(_05467_));
 sky130_fd_sc_hd__o211a_1 _12301_ (.A1(\rbzero.tex_g1[19] ),
    .A2(_05136_),
    .B1(_05467_),
    .C1(_05130_),
    .X(_05468_));
 sky130_fd_sc_hd__a31o_1 _12302_ (.A1(\rbzero.tex_g1[17] ),
    .A2(_05139_),
    .A3(_04927_),
    .B1(_05332_),
    .X(_05469_));
 sky130_fd_sc_hd__a311o_1 _12303_ (.A1(\rbzero.tex_g1[16] ),
    .A2(_04858_),
    .A3(_04813_),
    .B1(_05468_),
    .C1(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__or2_1 _12304_ (.A(\rbzero.tex_g1[30] ),
    .B(_04798_),
    .X(_05471_));
 sky130_fd_sc_hd__o211a_1 _12305_ (.A1(\rbzero.tex_g1[31] ),
    .A2(_05090_),
    .B1(_05471_),
    .C1(_05129_),
    .X(_05472_));
 sky130_fd_sc_hd__a31o_1 _12306_ (.A1(\rbzero.tex_g1[29] ),
    .A2(_04839_),
    .A3(_05145_),
    .B1(_04786_),
    .X(_05473_));
 sky130_fd_sc_hd__a311o_1 _12307_ (.A1(\rbzero.tex_g1[28] ),
    .A2(_05139_),
    .A3(_05132_),
    .B1(_05472_),
    .C1(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__or2_1 _12308_ (.A(\rbzero.tex_g1[26] ),
    .B(_04798_),
    .X(_05475_));
 sky130_fd_sc_hd__o211a_1 _12309_ (.A1(\rbzero.tex_g1[27] ),
    .A2(_05090_),
    .B1(_05475_),
    .C1(_05129_),
    .X(_05476_));
 sky130_fd_sc_hd__a31o_1 _12310_ (.A1(\rbzero.tex_g1[25] ),
    .A2(_04839_),
    .A3(_05145_),
    .B1(_04862_),
    .X(_05477_));
 sky130_fd_sc_hd__a311o_1 _12311_ (.A1(\rbzero.tex_g1[24] ),
    .A2(_04857_),
    .A3(_05132_),
    .B1(_05476_),
    .C1(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__a31o_1 _12312_ (.A1(_04865_),
    .A2(_05474_),
    .A3(_05478_),
    .B1(_04884_),
    .X(_05479_));
 sky130_fd_sc_hd__a31o_1 _12313_ (.A1(_04850_),
    .A2(_05466_),
    .A3(_05470_),
    .B1(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__a31o_1 _12314_ (.A1(_04908_),
    .A2(_05462_),
    .A3(_05480_),
    .B1(_04704_),
    .X(_05481_));
 sky130_fd_sc_hd__a21oi_1 _12315_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_04852_),
    .B1(_04703_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21a_1 _12316_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_04852_),
    .B1(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__a311oi_4 _12317_ (.A1(_04702_),
    .A2(_04706_),
    .A3(_04805_),
    .B1(_05483_),
    .C1(_04818_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21ba_1 _12318_ (.A1(_05444_),
    .A2(_05481_),
    .B1_N(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _12319_ (.A0(_05401_),
    .A1(_05485_),
    .S(_04989_),
    .X(_05486_));
 sky130_fd_sc_hd__inv_2 _12320_ (.A(_05193_),
    .Y(_05487_));
 sky130_fd_sc_hd__and2b_1 _12321_ (.A_N(_05194_),
    .B(_05025_),
    .X(_05488_));
 sky130_fd_sc_hd__a41o_1 _12322_ (.A1(_05011_),
    .A2(_05185_),
    .A3(_05487_),
    .A4(_05488_),
    .B1(_05066_),
    .X(_05489_));
 sky130_fd_sc_hd__o21a_1 _12323_ (.A1(_04699_),
    .A2(_05486_),
    .B1(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__o22a_1 _12324_ (.A1(\rbzero.trace_state[3] ),
    .A2(_04686_),
    .B1(_04688_),
    .B2(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__o21a_4 _12325_ (.A1(_04685_),
    .A2(_05491_),
    .B1(_05315_),
    .X(_05492_));
 sky130_fd_sc_hd__mux2_2 _12326_ (.A0(\reg_rgb[15] ),
    .A1(_05492_),
    .S(_05082_),
    .X(_05493_));
 sky130_fd_sc_hd__clkbuf_1 _12327_ (.A(_05493_),
    .X(net67));
 sky130_fd_sc_hd__nand2_1 _12328_ (.A(_04677_),
    .B(_04689_),
    .Y(_05494_));
 sky130_fd_sc_hd__o21a_1 _12329_ (.A1(_05185_),
    .A2(_05193_),
    .B1(_05488_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_04700_),
    .X(_05496_));
 sky130_fd_sc_hd__o21a_1 _12331_ (.A1(_04806_),
    .A2(_05323_),
    .B1(_05167_),
    .X(_05497_));
 sky130_fd_sc_hd__a311o_1 _12332_ (.A1(_04814_),
    .A2(\rbzero.row_render.wall[0] ),
    .A3(_04781_),
    .B1(_05327_),
    .C1(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__or2_1 _12333_ (.A(\rbzero.tex_b0[58] ),
    .B(_05144_),
    .X(_05499_));
 sky130_fd_sc_hd__o211a_1 _12334_ (.A1(\rbzero.tex_b0[59] ),
    .A2(_04833_),
    .B1(_05499_),
    .C1(_04777_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_4 _12335_ (.A(_05122_),
    .X(_05501_));
 sky130_fd_sc_hd__a31o_1 _12336_ (.A1(\rbzero.tex_b0[57] ),
    .A2(_04788_),
    .A3(_05501_),
    .B1(_04772_),
    .X(_05502_));
 sky130_fd_sc_hd__a31o_1 _12337_ (.A1(\rbzero.tex_b0[56] ),
    .A2(_04874_),
    .A3(_04833_),
    .B1(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__or2_1 _12338_ (.A(\rbzero.tex_b0[62] ),
    .B(_05144_),
    .X(_05504_));
 sky130_fd_sc_hd__o211a_1 _12339_ (.A1(\rbzero.tex_b0[63] ),
    .A2(_04833_),
    .B1(_05504_),
    .C1(_04777_),
    .X(_05505_));
 sky130_fd_sc_hd__a31o_1 _12340_ (.A1(\rbzero.tex_b0[61] ),
    .A2(_04788_),
    .A3(_05501_),
    .B1(_04785_),
    .X(_05506_));
 sky130_fd_sc_hd__a31o_1 _12341_ (.A1(\rbzero.tex_b0[60] ),
    .A2(_04789_),
    .A3(_04830_),
    .B1(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__o221a_1 _12342_ (.A1(_05500_),
    .A2(_05503_),
    .B1(_05505_),
    .B2(_05507_),
    .C1(_04865_),
    .X(_05508_));
 sky130_fd_sc_hd__or2_1 _12343_ (.A(\rbzero.tex_b0[54] ),
    .B(_05501_),
    .X(_05509_));
 sky130_fd_sc_hd__o211a_1 _12344_ (.A1(\rbzero.tex_b0[55] ),
    .A2(_04833_),
    .B1(_05509_),
    .C1(_04777_),
    .X(_05510_));
 sky130_fd_sc_hd__a31o_1 _12345_ (.A1(\rbzero.tex_b0[53] ),
    .A2(_04788_),
    .A3(_05501_),
    .B1(_04785_),
    .X(_05511_));
 sky130_fd_sc_hd__a31o_1 _12346_ (.A1(\rbzero.tex_b0[52] ),
    .A2(_04789_),
    .A3(_04830_),
    .B1(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__or2_1 _12347_ (.A(\rbzero.tex_b0[50] ),
    .B(_05501_),
    .X(_05513_));
 sky130_fd_sc_hd__o211a_1 _12348_ (.A1(\rbzero.tex_b0[51] ),
    .A2(_04830_),
    .B1(_05513_),
    .C1(_04844_),
    .X(_05514_));
 sky130_fd_sc_hd__a31o_1 _12349_ (.A1(\rbzero.tex_b0[49] ),
    .A2(_04788_),
    .A3(_05501_),
    .B1(_04862_),
    .X(_05515_));
 sky130_fd_sc_hd__a31o_1 _12350_ (.A1(\rbzero.tex_b0[48] ),
    .A2(_04789_),
    .A3(_04830_),
    .B1(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__o221a_1 _12351_ (.A1(_05510_),
    .A2(_05512_),
    .B1(_05514_),
    .B2(_05516_),
    .C1(_04849_),
    .X(_05517_));
 sky130_fd_sc_hd__or2_1 _12352_ (.A(\rbzero.tex_b0[42] ),
    .B(_05122_),
    .X(_05518_));
 sky130_fd_sc_hd__o211a_1 _12353_ (.A1(\rbzero.tex_b0[43] ),
    .A2(_04829_),
    .B1(_05518_),
    .C1(_05129_),
    .X(_05519_));
 sky130_fd_sc_hd__a31o_1 _12354_ (.A1(\rbzero.tex_b0[41] ),
    .A2(_04856_),
    .A3(_04799_),
    .B1(_04862_),
    .X(_05520_));
 sky130_fd_sc_hd__a311o_1 _12355_ (.A1(\rbzero.tex_b0[40] ),
    .A2(_05406_),
    .A3(_04853_),
    .B1(_05519_),
    .C1(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__or2_1 _12356_ (.A(\rbzero.tex_b0[46] ),
    .B(_05122_),
    .X(_05522_));
 sky130_fd_sc_hd__o211a_1 _12357_ (.A1(\rbzero.tex_b0[47] ),
    .A2(_04829_),
    .B1(_05522_),
    .C1(_05129_),
    .X(_05523_));
 sky130_fd_sc_hd__a31o_1 _12358_ (.A1(\rbzero.tex_b0[45] ),
    .A2(_04856_),
    .A3(_05123_),
    .B1(_04785_),
    .X(_05524_));
 sky130_fd_sc_hd__a311o_1 _12359_ (.A1(\rbzero.tex_b0[44] ),
    .A2(_05406_),
    .A3(_04853_),
    .B1(_05523_),
    .C1(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__or2_1 _12360_ (.A(\rbzero.tex_b0[38] ),
    .B(_04797_),
    .X(_05526_));
 sky130_fd_sc_hd__o211a_1 _12361_ (.A1(\rbzero.tex_b0[39] ),
    .A2(_04828_),
    .B1(_05526_),
    .C1(_04775_),
    .X(_05527_));
 sky130_fd_sc_hd__a31o_1 _12362_ (.A1(\rbzero.tex_b0[37] ),
    .A2(_04838_),
    .A3(_04798_),
    .B1(_04785_),
    .X(_05528_));
 sky130_fd_sc_hd__a311o_1 _12363_ (.A1(\rbzero.tex_b0[36] ),
    .A2(_04788_),
    .A3(_04829_),
    .B1(_05527_),
    .C1(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__or2_1 _12364_ (.A(\rbzero.tex_b0[34] ),
    .B(_04797_),
    .X(_05530_));
 sky130_fd_sc_hd__o211a_1 _12365_ (.A1(\rbzero.tex_b0[35] ),
    .A2(_04828_),
    .B1(_05530_),
    .C1(_04775_),
    .X(_05531_));
 sky130_fd_sc_hd__a31o_1 _12366_ (.A1(\rbzero.tex_b0[33] ),
    .A2(_04838_),
    .A3(_04798_),
    .B1(_04772_),
    .X(_05532_));
 sky130_fd_sc_hd__a311o_1 _12367_ (.A1(\rbzero.tex_b0[32] ),
    .A2(_04788_),
    .A3(_04829_),
    .B1(_05531_),
    .C1(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__a31o_1 _12368_ (.A1(_04783_),
    .A2(_05529_),
    .A3(_05533_),
    .B1(_04825_),
    .X(_05534_));
 sky130_fd_sc_hd__a31o_1 _12369_ (.A1(_04865_),
    .A2(_05521_),
    .A3(_05525_),
    .B1(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__o311a_1 _12370_ (.A1(_04885_),
    .A2(_05508_),
    .A3(_05517_),
    .B1(_04821_),
    .C1(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__or2_1 _12371_ (.A(\rbzero.tex_b0[10] ),
    .B(_05144_),
    .X(_05537_));
 sky130_fd_sc_hd__o211a_1 _12372_ (.A1(\rbzero.tex_b0[11] ),
    .A2(_04811_),
    .B1(_05537_),
    .C1(_04835_),
    .X(_05538_));
 sky130_fd_sc_hd__clkbuf_4 _12373_ (.A(_05144_),
    .X(_05539_));
 sky130_fd_sc_hd__a31o_1 _12374_ (.A1(\rbzero.tex_b0[9] ),
    .A2(_04874_),
    .A3(_05539_),
    .B1(_04773_),
    .X(_05540_));
 sky130_fd_sc_hd__a311o_1 _12375_ (.A1(\rbzero.tex_b0[8] ),
    .A2(_04840_),
    .A3(_04812_),
    .B1(_05538_),
    .C1(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__or2_1 _12376_ (.A(\rbzero.tex_b0[14] ),
    .B(_04798_),
    .X(_05542_));
 sky130_fd_sc_hd__o211a_1 _12377_ (.A1(\rbzero.tex_b0[15] ),
    .A2(_04811_),
    .B1(_05542_),
    .C1(_04835_),
    .X(_05543_));
 sky130_fd_sc_hd__a31o_1 _12378_ (.A1(\rbzero.tex_b0[13] ),
    .A2(_04874_),
    .A3(_05145_),
    .B1(_04786_),
    .X(_05544_));
 sky130_fd_sc_hd__a311o_1 _12379_ (.A1(\rbzero.tex_b0[12] ),
    .A2(_04840_),
    .A3(_04812_),
    .B1(_05543_),
    .C1(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__or2_1 _12380_ (.A(\rbzero.tex_b0[6] ),
    .B(_05144_),
    .X(_05546_));
 sky130_fd_sc_hd__o211a_1 _12381_ (.A1(\rbzero.tex_b0[7] ),
    .A2(_05370_),
    .B1(_05546_),
    .C1(_04777_),
    .X(_05547_));
 sky130_fd_sc_hd__a31o_1 _12382_ (.A1(\rbzero.tex_b0[5] ),
    .A2(_04838_),
    .A3(_05144_),
    .B1(_04785_),
    .X(_05548_));
 sky130_fd_sc_hd__a31o_1 _12383_ (.A1(\rbzero.tex_b0[4] ),
    .A2(_04839_),
    .A3(_05370_),
    .B1(_05548_),
    .X(_05549_));
 sky130_fd_sc_hd__or2_1 _12384_ (.A(\rbzero.tex_b0[2] ),
    .B(_05144_),
    .X(_05550_));
 sky130_fd_sc_hd__o211a_1 _12385_ (.A1(\rbzero.tex_b0[3] ),
    .A2(_05370_),
    .B1(_05550_),
    .C1(_04777_),
    .X(_05551_));
 sky130_fd_sc_hd__a31o_1 _12386_ (.A1(\rbzero.tex_b0[1] ),
    .A2(_04838_),
    .A3(_05144_),
    .B1(_04772_),
    .X(_05552_));
 sky130_fd_sc_hd__a31o_1 _12387_ (.A1(\rbzero.tex_b0[0] ),
    .A2(_04874_),
    .A3(_04833_),
    .B1(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__o221a_1 _12388_ (.A1(_05547_),
    .A2(_05549_),
    .B1(_05551_),
    .B2(_05553_),
    .C1(_04783_),
    .X(_05554_));
 sky130_fd_sc_hd__a31o_1 _12389_ (.A1(_04868_),
    .A2(_05541_),
    .A3(_05545_),
    .B1(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__or2_1 _12390_ (.A(\rbzero.tex_b0[22] ),
    .B(_04797_),
    .X(_05556_));
 sky130_fd_sc_hd__o211a_1 _12391_ (.A1(\rbzero.tex_b0[23] ),
    .A2(_05104_),
    .B1(_05556_),
    .C1(_04776_),
    .X(_05557_));
 sky130_fd_sc_hd__a31o_1 _12392_ (.A1(\rbzero.tex_b0[21] ),
    .A2(_04787_),
    .A3(_05122_),
    .B1(_04785_),
    .X(_05558_));
 sky130_fd_sc_hd__a31o_1 _12393_ (.A1(\rbzero.tex_b0[20] ),
    .A2(_04838_),
    .A3(_04810_),
    .B1(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__or2_1 _12394_ (.A(\rbzero.tex_b0[18] ),
    .B(_04797_),
    .X(_05560_));
 sky130_fd_sc_hd__o211a_1 _12395_ (.A1(\rbzero.tex_b0[19] ),
    .A2(_04810_),
    .B1(_05560_),
    .C1(_04776_),
    .X(_05561_));
 sky130_fd_sc_hd__a31o_1 _12396_ (.A1(\rbzero.tex_b0[17] ),
    .A2(_04787_),
    .A3(_05122_),
    .B1(_04772_),
    .X(_05562_));
 sky130_fd_sc_hd__a31o_1 _12397_ (.A1(\rbzero.tex_b0[16] ),
    .A2(_04838_),
    .A3(_04810_),
    .B1(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__o221a_1 _12398_ (.A1(_05557_),
    .A2(_05559_),
    .B1(_05561_),
    .B2(_05563_),
    .C1(_04783_),
    .X(_05564_));
 sky130_fd_sc_hd__or2_1 _12399_ (.A(\rbzero.tex_b0[26] ),
    .B(_04797_),
    .X(_05565_));
 sky130_fd_sc_hd__o211a_1 _12400_ (.A1(\rbzero.tex_b0[27] ),
    .A2(_05104_),
    .B1(_05565_),
    .C1(_04776_),
    .X(_05566_));
 sky130_fd_sc_hd__a31o_1 _12401_ (.A1(\rbzero.tex_b0[25] ),
    .A2(_04787_),
    .A3(_05122_),
    .B1(_04772_),
    .X(_05567_));
 sky130_fd_sc_hd__a31o_1 _12402_ (.A1(\rbzero.tex_b0[24] ),
    .A2(_04838_),
    .A3(_04810_),
    .B1(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__or2_1 _12403_ (.A(\rbzero.tex_b0[30] ),
    .B(_04797_),
    .X(_05569_));
 sky130_fd_sc_hd__o211a_1 _12404_ (.A1(\rbzero.tex_b0[31] ),
    .A2(_05104_),
    .B1(_05569_),
    .C1(_04776_),
    .X(_05570_));
 sky130_fd_sc_hd__a31o_1 _12405_ (.A1(\rbzero.tex_b0[29] ),
    .A2(_04787_),
    .A3(_05122_),
    .B1(_04785_),
    .X(_05571_));
 sky130_fd_sc_hd__a31o_1 _12406_ (.A1(\rbzero.tex_b0[28] ),
    .A2(_04838_),
    .A3(_04810_),
    .B1(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__o221a_1 _12407_ (.A1(_05566_),
    .A2(_05568_),
    .B1(_05570_),
    .B2(_05572_),
    .C1(_04770_),
    .X(_05573_));
 sky130_fd_sc_hd__or2_1 _12408_ (.A(_05564_),
    .B(_05573_),
    .X(_05574_));
 sky130_fd_sc_hd__and3_1 _12409_ (.A(_04826_),
    .B(_04908_),
    .C(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__a21oi_1 _12410_ (.A1(_04898_),
    .A2(_05555_),
    .B1(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__or2b_1 _12411_ (.A(_05536_),
    .B_N(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__a22o_1 _12412_ (.A1(_05322_),
    .A2(_05498_),
    .B1(_05577_),
    .B2(_04818_),
    .X(_05578_));
 sky130_fd_sc_hd__mux2_1 _12413_ (.A0(_05496_),
    .A1(_05578_),
    .S(_04989_),
    .X(_05579_));
 sky130_fd_sc_hd__or2_1 _12414_ (.A(_04699_),
    .B(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__o311a_1 _12415_ (.A1(_05319_),
    .A2(_05494_),
    .A3(_05495_),
    .B1(_05580_),
    .C1(_05320_),
    .X(_05581_));
 sky130_fd_sc_hd__o21a_4 _12416_ (.A1(_04685_),
    .A2(_05581_),
    .B1(_05080_),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_4 _12417_ (.A0(\reg_rgb[22] ),
    .A1(_05582_),
    .S(_05082_),
    .X(_05583_));
 sky130_fd_sc_hd__clkbuf_1 _12418_ (.A(_05583_),
    .X(net68));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_04700_),
    .X(_05584_));
 sky130_fd_sc_hd__or2_1 _12420_ (.A(\rbzero.tex_b1[22] ),
    .B(_05539_),
    .X(_05585_));
 sky130_fd_sc_hd__o211a_1 _12421_ (.A1(\rbzero.tex_b1[23] ),
    .A2(_04895_),
    .B1(_05585_),
    .C1(_04836_),
    .X(_05586_));
 sky130_fd_sc_hd__a31o_1 _12422_ (.A1(\rbzero.tex_b1[21] ),
    .A2(_04789_),
    .A3(_05403_),
    .B1(_05409_),
    .X(_05587_));
 sky130_fd_sc_hd__a31o_1 _12423_ (.A1(\rbzero.tex_b1[20] ),
    .A2(_05407_),
    .A3(_04888_),
    .B1(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__or2_1 _12424_ (.A(\rbzero.tex_b1[18] ),
    .B(_05539_),
    .X(_05589_));
 sky130_fd_sc_hd__o211a_1 _12425_ (.A1(\rbzero.tex_b1[19] ),
    .A2(_04888_),
    .B1(_05589_),
    .C1(_04836_),
    .X(_05590_));
 sky130_fd_sc_hd__a31o_1 _12426_ (.A1(\rbzero.tex_b1[17] ),
    .A2(_05406_),
    .A3(_05403_),
    .B1(_04773_),
    .X(_05591_));
 sky130_fd_sc_hd__a31o_1 _12427_ (.A1(\rbzero.tex_b1[16] ),
    .A2(_05407_),
    .A3(_04888_),
    .B1(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__o221a_1 _12428_ (.A1(_05586_),
    .A2(_05588_),
    .B1(_05590_),
    .B2(_05592_),
    .C1(_04850_),
    .X(_05593_));
 sky130_fd_sc_hd__or2_1 _12429_ (.A(\rbzero.tex_b1[26] ),
    .B(_05501_),
    .X(_05594_));
 sky130_fd_sc_hd__o211a_1 _12430_ (.A1(\rbzero.tex_b1[27] ),
    .A2(_04830_),
    .B1(_05594_),
    .C1(_04844_),
    .X(_05595_));
 sky130_fd_sc_hd__a31o_1 _12431_ (.A1(\rbzero.tex_b1[25] ),
    .A2(_04789_),
    .A3(_05403_),
    .B1(_04773_),
    .X(_05596_));
 sky130_fd_sc_hd__a311o_1 _12432_ (.A1(\rbzero.tex_b1[24] ),
    .A2(_05089_),
    .A3(_04895_),
    .B1(_05595_),
    .C1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__or2_1 _12433_ (.A(\rbzero.tex_b1[30] ),
    .B(_05501_),
    .X(_05598_));
 sky130_fd_sc_hd__o211a_1 _12434_ (.A1(\rbzero.tex_b1[31] ),
    .A2(_04830_),
    .B1(_05598_),
    .C1(_04777_),
    .X(_05599_));
 sky130_fd_sc_hd__a31o_1 _12435_ (.A1(\rbzero.tex_b1[29] ),
    .A2(_04789_),
    .A3(_05403_),
    .B1(_05409_),
    .X(_05600_));
 sky130_fd_sc_hd__a311o_1 _12436_ (.A1(\rbzero.tex_b1[28] ),
    .A2(_05089_),
    .A3(_04895_),
    .B1(_05599_),
    .C1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__a31o_1 _12437_ (.A1(_04868_),
    .A2(_05597_),
    .A3(_05601_),
    .B1(_04885_),
    .X(_05602_));
 sky130_fd_sc_hd__or2_1 _12438_ (.A(\rbzero.tex_b1[10] ),
    .B(_05539_),
    .X(_05603_));
 sky130_fd_sc_hd__o211a_1 _12439_ (.A1(\rbzero.tex_b1[11] ),
    .A2(_04888_),
    .B1(_05603_),
    .C1(_04890_),
    .X(_05604_));
 sky130_fd_sc_hd__a31o_1 _12440_ (.A1(\rbzero.tex_b1[9] ),
    .A2(_05406_),
    .A3(_05403_),
    .B1(_04773_),
    .X(_05605_));
 sky130_fd_sc_hd__a31o_1 _12441_ (.A1(\rbzero.tex_b1[8] ),
    .A2(_05407_),
    .A3(_04888_),
    .B1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__or2_1 _12442_ (.A(\rbzero.tex_b1[14] ),
    .B(_05403_),
    .X(_05607_));
 sky130_fd_sc_hd__o211a_1 _12443_ (.A1(\rbzero.tex_b1[15] ),
    .A2(_04888_),
    .B1(_05607_),
    .C1(_04890_),
    .X(_05608_));
 sky130_fd_sc_hd__a31o_1 _12444_ (.A1(\rbzero.tex_b1[13] ),
    .A2(_05406_),
    .A3(_05408_),
    .B1(_05409_),
    .X(_05609_));
 sky130_fd_sc_hd__a31o_1 _12445_ (.A1(\rbzero.tex_b1[12] ),
    .A2(_05407_),
    .A3(_05402_),
    .B1(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__o221a_1 _12446_ (.A1(_05604_),
    .A2(_05606_),
    .B1(_05608_),
    .B2(_05610_),
    .C1(_04868_),
    .X(_05611_));
 sky130_fd_sc_hd__or2_1 _12447_ (.A(\rbzero.tex_b1[6] ),
    .B(_05501_),
    .X(_05612_));
 sky130_fd_sc_hd__o211a_1 _12448_ (.A1(\rbzero.tex_b1[7] ),
    .A2(_04830_),
    .B1(_05612_),
    .C1(_04844_),
    .X(_05613_));
 sky130_fd_sc_hd__a31o_1 _12449_ (.A1(\rbzero.tex_b1[5] ),
    .A2(_05406_),
    .A3(_05403_),
    .B1(_05409_),
    .X(_05614_));
 sky130_fd_sc_hd__a311o_1 _12450_ (.A1(\rbzero.tex_b1[4] ),
    .A2(_05407_),
    .A3(_04895_),
    .B1(_05613_),
    .C1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__or2_1 _12451_ (.A(\rbzero.tex_b1[2] ),
    .B(_05501_),
    .X(_05616_));
 sky130_fd_sc_hd__o211a_1 _12452_ (.A1(\rbzero.tex_b1[3] ),
    .A2(_04830_),
    .B1(_05616_),
    .C1(_04844_),
    .X(_05617_));
 sky130_fd_sc_hd__a31o_1 _12453_ (.A1(\rbzero.tex_b1[1] ),
    .A2(_05406_),
    .A3(_05403_),
    .B1(_05332_),
    .X(_05618_));
 sky130_fd_sc_hd__a311o_1 _12454_ (.A1(\rbzero.tex_b1[0] ),
    .A2(_05407_),
    .A3(_04895_),
    .B1(_05617_),
    .C1(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__a31o_1 _12455_ (.A1(_04850_),
    .A2(_05615_),
    .A3(_05619_),
    .B1(_04826_),
    .X(_05620_));
 sky130_fd_sc_hd__o221a_1 _12456_ (.A1(_05593_),
    .A2(_05602_),
    .B1(_05611_),
    .B2(_05620_),
    .C1(_04908_),
    .X(_05621_));
 sky130_fd_sc_hd__or2_1 _12457_ (.A(\rbzero.tex_b1[54] ),
    .B(_05539_),
    .X(_05622_));
 sky130_fd_sc_hd__o211a_1 _12458_ (.A1(\rbzero.tex_b1[55] ),
    .A2(_04895_),
    .B1(_05622_),
    .C1(_04836_),
    .X(_05623_));
 sky130_fd_sc_hd__a31o_1 _12459_ (.A1(\rbzero.tex_b1[53] ),
    .A2(_04789_),
    .A3(_05539_),
    .B1(_04786_),
    .X(_05624_));
 sky130_fd_sc_hd__a31o_1 _12460_ (.A1(\rbzero.tex_b1[52] ),
    .A2(_05089_),
    .A3(_04895_),
    .B1(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__or2_1 _12461_ (.A(\rbzero.tex_b1[50] ),
    .B(_05539_),
    .X(_05626_));
 sky130_fd_sc_hd__o211a_1 _12462_ (.A1(\rbzero.tex_b1[51] ),
    .A2(_04895_),
    .B1(_05626_),
    .C1(_04836_),
    .X(_05627_));
 sky130_fd_sc_hd__a31o_1 _12463_ (.A1(\rbzero.tex_b1[49] ),
    .A2(_04789_),
    .A3(_05539_),
    .B1(_04773_),
    .X(_05628_));
 sky130_fd_sc_hd__a31o_1 _12464_ (.A1(\rbzero.tex_b1[48] ),
    .A2(_05407_),
    .A3(_04888_),
    .B1(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__o221a_1 _12465_ (.A1(_05623_),
    .A2(_05625_),
    .B1(_05627_),
    .B2(_05629_),
    .C1(_04849_),
    .X(_05630_));
 sky130_fd_sc_hd__or2_1 _12466_ (.A(\rbzero.tex_b1[58] ),
    .B(_05539_),
    .X(_05631_));
 sky130_fd_sc_hd__o211a_1 _12467_ (.A1(\rbzero.tex_b1[59] ),
    .A2(_04895_),
    .B1(_05631_),
    .C1(_04836_),
    .X(_05632_));
 sky130_fd_sc_hd__a31o_1 _12468_ (.A1(\rbzero.tex_b1[57] ),
    .A2(_04789_),
    .A3(_05403_),
    .B1(_04773_),
    .X(_05633_));
 sky130_fd_sc_hd__a31o_1 _12469_ (.A1(\rbzero.tex_b1[56] ),
    .A2(_05407_),
    .A3(_04888_),
    .B1(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__or2_1 _12470_ (.A(\rbzero.tex_b1[62] ),
    .B(_05539_),
    .X(_05635_));
 sky130_fd_sc_hd__o211a_1 _12471_ (.A1(\rbzero.tex_b1[63] ),
    .A2(_04888_),
    .B1(_05635_),
    .C1(_04890_),
    .X(_05636_));
 sky130_fd_sc_hd__a31o_1 _12472_ (.A1(\rbzero.tex_b1[61] ),
    .A2(_05406_),
    .A3(_05408_),
    .B1(_05409_),
    .X(_05637_));
 sky130_fd_sc_hd__a31o_1 _12473_ (.A1(\rbzero.tex_b1[60] ),
    .A2(_05407_),
    .A3(_05402_),
    .B1(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__o221a_1 _12474_ (.A1(_05632_),
    .A2(_05634_),
    .B1(_05636_),
    .B2(_05638_),
    .C1(_04868_),
    .X(_05639_));
 sky130_fd_sc_hd__or2_1 _12475_ (.A(\rbzero.tex_b1[42] ),
    .B(_05123_),
    .X(_05640_));
 sky130_fd_sc_hd__o211a_1 _12476_ (.A1(\rbzero.tex_b1[43] ),
    .A2(_05121_),
    .B1(_05640_),
    .C1(_05130_),
    .X(_05641_));
 sky130_fd_sc_hd__a31o_1 _12477_ (.A1(\rbzero.tex_b1[41] ),
    .A2(_05139_),
    .A3(_04927_),
    .B1(_05332_),
    .X(_05642_));
 sky130_fd_sc_hd__a311o_1 _12478_ (.A1(\rbzero.tex_b1[40] ),
    .A2(_04858_),
    .A3(_04813_),
    .B1(_05641_),
    .C1(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__or2_1 _12479_ (.A(\rbzero.tex_b1[46] ),
    .B(_05123_),
    .X(_05644_));
 sky130_fd_sc_hd__o211a_1 _12480_ (.A1(\rbzero.tex_b1[47] ),
    .A2(_05121_),
    .B1(_05644_),
    .C1(_05130_),
    .X(_05645_));
 sky130_fd_sc_hd__a31o_1 _12481_ (.A1(\rbzero.tex_b1[45] ),
    .A2(_05139_),
    .A3(_05408_),
    .B1(_05409_),
    .X(_05646_));
 sky130_fd_sc_hd__a311o_1 _12482_ (.A1(\rbzero.tex_b1[44] ),
    .A2(_04858_),
    .A3(_05402_),
    .B1(_05645_),
    .C1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__or2_1 _12483_ (.A(\rbzero.tex_b1[38] ),
    .B(_05122_),
    .X(_05648_));
 sky130_fd_sc_hd__o211a_1 _12484_ (.A1(\rbzero.tex_b1[39] ),
    .A2(_05085_),
    .B1(_05648_),
    .C1(_05129_),
    .X(_05649_));
 sky130_fd_sc_hd__a31o_1 _12485_ (.A1(\rbzero.tex_b1[37] ),
    .A2(_04856_),
    .A3(_05145_),
    .B1(_04786_),
    .X(_05650_));
 sky130_fd_sc_hd__a311o_1 _12486_ (.A1(\rbzero.tex_b1[36] ),
    .A2(_04857_),
    .A3(_05136_),
    .B1(_05649_),
    .C1(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__or2_1 _12487_ (.A(\rbzero.tex_b1[34] ),
    .B(_05122_),
    .X(_05652_));
 sky130_fd_sc_hd__o211a_1 _12488_ (.A1(\rbzero.tex_b1[35] ),
    .A2(_05085_),
    .B1(_05652_),
    .C1(_05129_),
    .X(_05653_));
 sky130_fd_sc_hd__a31o_1 _12489_ (.A1(\rbzero.tex_b1[33] ),
    .A2(_04856_),
    .A3(_04799_),
    .B1(_04862_),
    .X(_05654_));
 sky130_fd_sc_hd__a311o_1 _12490_ (.A1(\rbzero.tex_b1[32] ),
    .A2(_04857_),
    .A3(_05136_),
    .B1(_05653_),
    .C1(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__a31o_1 _12491_ (.A1(_04849_),
    .A2(_05651_),
    .A3(_05655_),
    .B1(_04825_),
    .X(_05656_));
 sky130_fd_sc_hd__a31o_1 _12492_ (.A1(_04868_),
    .A2(_05643_),
    .A3(_05647_),
    .B1(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__o311a_1 _12493_ (.A1(_04885_),
    .A2(_05630_),
    .A3(_05639_),
    .B1(_04821_),
    .C1(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__o21a_1 _12494_ (.A1(_05621_),
    .A2(_05658_),
    .B1(_04818_),
    .X(_05659_));
 sky130_fd_sc_hd__and2_1 _12495_ (.A(\rbzero.row_render.texu[0] ),
    .B(_04927_),
    .X(_05660_));
 sky130_fd_sc_hd__nor2_1 _12496_ (.A(_04800_),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__or3b_1 _12497_ (.A(_04780_),
    .B(_04702_),
    .C_N(\rbzero.row_render.wall[1] ),
    .X(_05662_));
 sky130_fd_sc_hd__o21ai_1 _12498_ (.A1(_04804_),
    .A2(_04800_),
    .B1(_04702_),
    .Y(_05663_));
 sky130_fd_sc_hd__o21ai_1 _12499_ (.A1(_04807_),
    .A2(_04804_),
    .B1(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__a22o_1 _12500_ (.A1(\rbzero.row_render.wall[0] ),
    .A2(_05662_),
    .B1(_05664_),
    .B2(_04706_),
    .X(_05665_));
 sky130_fd_sc_hd__o211a_1 _12501_ (.A1(_04703_),
    .A2(_05661_),
    .B1(_05665_),
    .C1(_04704_),
    .X(_05666_));
 sky130_fd_sc_hd__or3b_1 _12502_ (.A(_05659_),
    .B(_05666_),
    .C_N(_04989_),
    .X(_05667_));
 sky130_fd_sc_hd__o211a_1 _12503_ (.A1(_04989_),
    .A2(_05584_),
    .B1(_05667_),
    .C1(_05319_),
    .X(_05668_));
 sky130_fd_sc_hd__and3_1 _12504_ (.A(_04699_),
    .B(_05011_),
    .C(_05495_),
    .X(_05669_));
 sky130_fd_sc_hd__o21ba_1 _12505_ (.A1(_05668_),
    .A2(_05669_),
    .B1_N(_04688_),
    .X(_05670_));
 sky130_fd_sc_hd__o21a_4 _12506_ (.A1(_04685_),
    .A2(_05670_),
    .B1(_05315_),
    .X(_05671_));
 sky130_fd_sc_hd__mux2_4 _12507_ (.A0(\reg_rgb[23] ),
    .A1(_05671_),
    .S(_05082_),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _12508_ (.A(_05672_),
    .X(net69));
 sky130_fd_sc_hd__mux2_2 _12509_ (.A0(reg_vsync),
    .A1(_04466_),
    .S(_05082_),
    .X(_05673_));
 sky130_fd_sc_hd__clkbuf_1 _12510_ (.A(_05673_),
    .X(net76));
 sky130_fd_sc_hd__clkinv_2 _12511_ (.A(\rbzero.hsync ),
    .Y(_05674_));
 sky130_fd_sc_hd__mux2_2 _12512_ (.A0(reg_hsync),
    .A1(_05674_),
    .S(_05082_),
    .X(_05675_));
 sky130_fd_sc_hd__clkbuf_1 _12513_ (.A(_05675_),
    .X(net64));
 sky130_fd_sc_hd__inv_2 _12514_ (.A(net8),
    .Y(_05676_));
 sky130_fd_sc_hd__clkbuf_4 _12515_ (.A(net4),
    .X(_05677_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(_05081_),
    .A1(_05317_),
    .S(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__mux4_1 _12517_ (.A0(_05399_),
    .A1(_05492_),
    .A2(_05582_),
    .A3(_05671_),
    .S0(_05677_),
    .S1(net7),
    .X(_05679_));
 sky130_fd_sc_hd__and2_1 _12518_ (.A(net8),
    .B(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__a31o_1 _12519_ (.A1(net7),
    .A2(_05676_),
    .A3(_05678_),
    .B1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__and4b_1 _12520_ (.A_N(net9),
    .B(_05681_),
    .C(net5),
    .D(net6),
    .X(_05682_));
 sky130_fd_sc_hd__and2b_1 _12521_ (.A_N(net7),
    .B(net6),
    .X(_05683_));
 sky130_fd_sc_hd__nor2_1 _12522_ (.A(net5),
    .B(_05677_),
    .Y(_05684_));
 sky130_fd_sc_hd__and2b_1 _12523_ (.A_N(net5),
    .B(_05677_),
    .X(_05685_));
 sky130_fd_sc_hd__a22o_1 _12524_ (.A1(_05079_),
    .A2(_05684_),
    .B1(_05685_),
    .B2(net73),
    .X(_05686_));
 sky130_fd_sc_hd__and2b_1 _12525_ (.A_N(net4),
    .B(net5),
    .X(_05687_));
 sky130_fd_sc_hd__and2_1 _12526_ (.A(net5),
    .B(net4),
    .X(_05688_));
 sky130_fd_sc_hd__a22o_1 _12527_ (.A1(net44),
    .A2(_05687_),
    .B1(_05688_),
    .B2(_05077_),
    .X(_05689_));
 sky130_fd_sc_hd__nor2_1 _12528_ (.A(net7),
    .B(net6),
    .Y(_05690_));
 sky130_fd_sc_hd__a22o_1 _12529_ (.A1(_05683_),
    .A2(_05686_),
    .B1(_05689_),
    .B2(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__nor2_1 _12530_ (.A(net9),
    .B(net8),
    .Y(_05692_));
 sky130_fd_sc_hd__a22o_1 _12531_ (.A1(net54),
    .A2(_05684_),
    .B1(_05687_),
    .B2(net57),
    .X(_05693_));
 sky130_fd_sc_hd__a21o_1 _12532_ (.A1(net55),
    .A2(_05685_),
    .B1(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__a21oi_2 _12533_ (.A1(net129),
    .A2(net5),
    .B1(_05677_),
    .Y(_05695_));
 sky130_fd_sc_hd__a221o_2 _12534_ (.A1(_04094_),
    .A2(_05685_),
    .B1(_05688_),
    .B2(\gpout0.clk_div[1] ),
    .C1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__a22o_2 _12535_ (.A1(_05683_),
    .A2(_05694_),
    .B1(_05696_),
    .B2(_05690_),
    .X(_05697_));
 sky130_fd_sc_hd__clkbuf_8 _12536_ (.A(net56),
    .X(_05698_));
 sky130_fd_sc_hd__a21o_1 _12537_ (.A1(_05698_),
    .A2(_05692_),
    .B1(net52),
    .X(_05699_));
 sky130_fd_sc_hd__a22o_1 _12538_ (.A1(net51),
    .A2(_05687_),
    .B1(_05688_),
    .B2(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__nand2_1 _12539_ (.A(_05700_),
    .B(_05683_),
    .Y(_05701_));
 sky130_fd_sc_hd__a22o_1 _12540_ (.A1(net41),
    .A2(_05687_),
    .B1(_05688_),
    .B2(_04704_),
    .X(_05702_));
 sky130_fd_sc_hd__a221o_1 _12541_ (.A1(net53),
    .A2(_05684_),
    .B1(_05685_),
    .B2(net40),
    .C1(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__inv_2 _12542_ (.A(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__a221oi_1 _12543_ (.A1(net43),
    .A2(_05684_),
    .B1(_05685_),
    .B2(net46),
    .C1(net7),
    .Y(_05705_));
 sky130_fd_sc_hd__a211o_1 _12544_ (.A1(net7),
    .A2(_05704_),
    .B1(_05705_),
    .C1(net6),
    .X(_05706_));
 sky130_fd_sc_hd__and4_1 _12545_ (.A(_05698_),
    .B(_05688_),
    .C(_05692_),
    .D(_05683_),
    .X(_05707_));
 sky130_fd_sc_hd__a21oi_1 _12546_ (.A1(net9),
    .A2(_05676_),
    .B1(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__a21oi_1 _12547_ (.A1(_05701_),
    .A2(_05706_),
    .B1(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__a21o_1 _12548_ (.A1(net5),
    .A2(net6),
    .B1(net7),
    .X(_05710_));
 sky130_fd_sc_hd__buf_2 _12549_ (.A(_04678_),
    .X(_05711_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(_04675_),
    .A1(_05711_),
    .S(_05677_),
    .X(_05712_));
 sky130_fd_sc_hd__mux2_1 _12551_ (.A0(_04683_),
    .A1(_04671_),
    .S(_05677_),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(_05186_),
    .A1(_05016_),
    .S(_05677_),
    .X(_05714_));
 sky130_fd_sc_hd__buf_2 _12553_ (.A(\gpout0.vpos[8] ),
    .X(_05715_));
 sky130_fd_sc_hd__buf_2 _12554_ (.A(\gpout0.vpos[9] ),
    .X(_05716_));
 sky130_fd_sc_hd__mux4_1 _12555_ (.A0(\gpout0.vpos[0] ),
    .A1(\gpout0.vpos[1] ),
    .A2(_05715_),
    .A3(_05716_),
    .S0(_05677_),
    .S1(net7),
    .X(_05717_));
 sky130_fd_sc_hd__mux4_1 _12556_ (.A0(_05712_),
    .A1(_05713_),
    .A2(_05714_),
    .A3(_05717_),
    .S0(net6),
    .S1(net5),
    .X(_05718_));
 sky130_fd_sc_hd__mux4_1 _12557_ (.A0(_04484_),
    .A1(_04452_),
    .A2(_04458_),
    .A3(_04014_),
    .S0(_05677_),
    .S1(net5),
    .X(_05719_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(_04017_),
    .A1(_04018_),
    .S(net4),
    .X(_05720_));
 sky130_fd_sc_hd__mux4_1 _12559_ (.A0(_04010_),
    .A1(_04584_),
    .A2(\gpout0.hpos[2] ),
    .A3(_04482_),
    .S0(net4),
    .S1(net5),
    .X(_05721_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(_05720_),
    .A1(_05721_),
    .S(net7),
    .X(_05722_));
 sky130_fd_sc_hd__or2b_1 _12561_ (.A(_05722_),
    .B_N(net6),
    .X(_05723_));
 sky130_fd_sc_hd__nor2_1 _12562_ (.A(_05676_),
    .B(_05710_),
    .Y(_05724_));
 sky130_fd_sc_hd__a31o_1 _12563_ (.A1(net7),
    .A2(net6),
    .A3(_05676_),
    .B1(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__o2111a_1 _12564_ (.A1(net6),
    .A2(_05719_),
    .B1(_05723_),
    .C1(net9),
    .D1(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__a41o_1 _12565_ (.A1(net9),
    .A2(net8),
    .A3(_05710_),
    .A4(_05718_),
    .B1(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__a211o_2 _12566_ (.A1(_05692_),
    .A2(_05697_),
    .B1(_05709_),
    .C1(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__a31o_2 _12567_ (.A1(net9),
    .A2(_05676_),
    .A3(_05691_),
    .B1(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__nand3_1 _12568_ (.A(_05684_),
    .B(_05692_),
    .C(_05690_),
    .Y(_05730_));
 sky130_fd_sc_hd__o22a_2 _12569_ (.A1(_05682_),
    .A2(_05729_),
    .B1(_05730_),
    .B2(_05399_),
    .X(_05731_));
 sky130_fd_sc_hd__mux2_2 _12570_ (.A0(\reg_gpout[0] ),
    .A1(clknet_1_0__leaf__05731_),
    .S(_05082_),
    .X(_05732_));
 sky130_fd_sc_hd__buf_1 _12571_ (.A(_05732_),
    .X(net58));
 sky130_fd_sc_hd__and2b_1 _12572_ (.A_N(net14),
    .B(net13),
    .X(_05733_));
 sky130_fd_sc_hd__clkbuf_4 _12573_ (.A(net10),
    .X(_05734_));
 sky130_fd_sc_hd__mux2_1 _12574_ (.A0(_05081_),
    .A1(_05317_),
    .S(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__mux4_1 _12575_ (.A0(_05399_),
    .A1(_05492_),
    .A2(_05582_),
    .A3(_05671_),
    .S0(_05734_),
    .S1(net13),
    .X(_05736_));
 sky130_fd_sc_hd__a22o_1 _12576_ (.A1(_05733_),
    .A2(_05735_),
    .B1(_05736_),
    .B2(net14),
    .X(_05737_));
 sky130_fd_sc_hd__and4b_1 _12577_ (.A_N(net15),
    .B(_05737_),
    .C(net11),
    .D(net12),
    .X(_05738_));
 sky130_fd_sc_hd__and2b_1 _12578_ (.A_N(net14),
    .B(net15),
    .X(_05739_));
 sky130_fd_sc_hd__inv_2 _12579_ (.A(net12),
    .Y(_05740_));
 sky130_fd_sc_hd__nor2_1 _12580_ (.A(net13),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__nor2_2 _12581_ (.A(net11),
    .B(net10),
    .Y(_05742_));
 sky130_fd_sc_hd__inv_2 _12582_ (.A(net11),
    .Y(_05743_));
 sky130_fd_sc_hd__and2_1 _12583_ (.A(_05743_),
    .B(net10),
    .X(_05744_));
 sky130_fd_sc_hd__a22o_1 _12584_ (.A1(_05079_),
    .A2(_05742_),
    .B1(_05744_),
    .B2(net73),
    .X(_05745_));
 sky130_fd_sc_hd__nor2_2 _12585_ (.A(_05743_),
    .B(_05734_),
    .Y(_05746_));
 sky130_fd_sc_hd__and2_1 _12586_ (.A(net11),
    .B(net10),
    .X(_05747_));
 sky130_fd_sc_hd__a22o_1 _12587_ (.A1(net44),
    .A2(_05746_),
    .B1(_05747_),
    .B2(_05077_),
    .X(_05748_));
 sky130_fd_sc_hd__nor2_1 _12588_ (.A(net13),
    .B(net12),
    .Y(_05749_));
 sky130_fd_sc_hd__a22o_1 _12589_ (.A1(_05741_),
    .A2(_05745_),
    .B1(_05748_),
    .B2(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__nor2_1 _12590_ (.A(net15),
    .B(net14),
    .Y(_05751_));
 sky130_fd_sc_hd__a41o_1 _12591_ (.A1(_05698_),
    .A2(_05751_),
    .A3(_05747_),
    .A4(_05741_),
    .B1(_05739_),
    .X(_05752_));
 sky130_fd_sc_hd__a21o_1 _12592_ (.A1(net56),
    .A2(_05751_),
    .B1(net52),
    .X(_05753_));
 sky130_fd_sc_hd__a22o_1 _12593_ (.A1(net51),
    .A2(_05746_),
    .B1(_05747_),
    .B2(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__a22o_1 _12594_ (.A1(net43),
    .A2(_05742_),
    .B1(_05744_),
    .B2(net46),
    .X(_05755_));
 sky130_fd_sc_hd__a22o_1 _12595_ (.A1(net53),
    .A2(_05742_),
    .B1(_05744_),
    .B2(net40),
    .X(_05756_));
 sky130_fd_sc_hd__a221o_1 _12596_ (.A1(net41),
    .A2(_05746_),
    .B1(_05747_),
    .B2(_04704_),
    .C1(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__mux2_1 _12597_ (.A0(_05755_),
    .A1(_05757_),
    .S(net13),
    .X(_05758_));
 sky130_fd_sc_hd__a22o_1 _12598_ (.A1(_05754_),
    .A2(_05741_),
    .B1(_05758_),
    .B2(_05740_),
    .X(_05759_));
 sky130_fd_sc_hd__a22o_1 _12599_ (.A1(net57),
    .A2(_05746_),
    .B1(_05744_),
    .B2(net55),
    .X(_05760_));
 sky130_fd_sc_hd__a21o_1 _12600_ (.A1(net54),
    .A2(_05742_),
    .B1(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__buf_1 _12601_ (.A(clknet_opt_8_0_i_clk),
    .X(_05762_));
 sky130_fd_sc_hd__a221o_2 _12602_ (.A1(_05743_),
    .A2(net50),
    .B1(_05746_),
    .B2(clknet_1_0__leaf__05762_),
    .C1(_05742_),
    .X(_05763_));
 sky130_fd_sc_hd__a21o_2 _12603_ (.A1(\gpout1.clk_div[1] ),
    .A2(_05747_),
    .B1(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__a22o_2 _12604_ (.A1(_05741_),
    .A2(_05761_),
    .B1(_05764_),
    .B2(_05749_),
    .X(_05765_));
 sky130_fd_sc_hd__a22o_2 _12605_ (.A1(_05752_),
    .A2(_05759_),
    .B1(_05765_),
    .B2(_05751_),
    .X(_05766_));
 sky130_fd_sc_hd__a21o_1 _12606_ (.A1(net11),
    .A2(net12),
    .B1(net13),
    .X(_05767_));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(_05186_),
    .A1(_05016_),
    .S(_05734_),
    .X(_05768_));
 sky130_fd_sc_hd__buf_2 _12608_ (.A(\gpout0.vpos[0] ),
    .X(_05769_));
 sky130_fd_sc_hd__buf_2 _12609_ (.A(\gpout0.vpos[1] ),
    .X(_05770_));
 sky130_fd_sc_hd__mux4_1 _12610_ (.A0(_05769_),
    .A1(_05770_),
    .A2(_05715_),
    .A3(_05716_),
    .S0(_05734_),
    .S1(net13),
    .X(_05771_));
 sky130_fd_sc_hd__mux2_1 _12611_ (.A0(_04675_),
    .A1(_05711_),
    .S(_05734_),
    .X(_05772_));
 sky130_fd_sc_hd__mux2_1 _12612_ (.A0(_04683_),
    .A1(_04671_),
    .S(_05734_),
    .X(_05773_));
 sky130_fd_sc_hd__mux4_1 _12613_ (.A0(_05768_),
    .A1(_05771_),
    .A2(_05772_),
    .A3(_05773_),
    .S0(net12),
    .S1(_05743_),
    .X(_05774_));
 sky130_fd_sc_hd__mux2_1 _12614_ (.A0(_04017_),
    .A1(_04018_),
    .S(_05734_),
    .X(_05775_));
 sky130_fd_sc_hd__mux4_1 _12615_ (.A0(_04010_),
    .A1(_04584_),
    .A2(_04587_),
    .A3(_04482_),
    .S0(_05734_),
    .S1(net11),
    .X(_05776_));
 sky130_fd_sc_hd__mux2_1 _12616_ (.A0(_05775_),
    .A1(_05776_),
    .S(net13),
    .X(_05777_));
 sky130_fd_sc_hd__mux4_1 _12617_ (.A0(_04484_),
    .A1(_04452_),
    .A2(_04458_),
    .A3(_04014_),
    .S0(_05734_),
    .S1(net11),
    .X(_05778_));
 sky130_fd_sc_hd__or2_1 _12618_ (.A(net12),
    .B(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__a21oi_1 _12619_ (.A1(net13),
    .A2(net12),
    .B1(net14),
    .Y(_05780_));
 sky130_fd_sc_hd__a21oi_1 _12620_ (.A1(net14),
    .A2(_05767_),
    .B1(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__o2111a_1 _12621_ (.A1(_05740_),
    .A2(_05777_),
    .B1(_05779_),
    .C1(net15),
    .D1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__a41o_1 _12622_ (.A1(net15),
    .A2(net14),
    .A3(_05767_),
    .A4(_05774_),
    .B1(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__a211o_2 _12623_ (.A1(_05739_),
    .A2(_05750_),
    .B1(_05766_),
    .C1(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__and4b_1 _12624_ (.A_N(_05492_),
    .B(_05751_),
    .C(_05742_),
    .D(_05749_),
    .X(_05785_));
 sky130_fd_sc_hd__o21ba_2 _12625_ (.A1(_05738_),
    .A2(_05784_),
    .B1_N(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__mux2_2 _12626_ (.A0(\reg_gpout[1] ),
    .A1(clknet_1_0__leaf__05786_),
    .S(_05082_),
    .X(_05787_));
 sky130_fd_sc_hd__buf_1 _12627_ (.A(_05787_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 _12628_ (.A(net16),
    .X(_05788_));
 sky130_fd_sc_hd__mux4_1 _12629_ (.A0(_05399_),
    .A1(_05492_),
    .A2(_05582_),
    .A3(_05671_),
    .S0(_05788_),
    .S1(net19),
    .X(_05789_));
 sky130_fd_sc_hd__inv_2 _12630_ (.A(net19),
    .Y(_05790_));
 sky130_fd_sc_hd__nor2_1 _12631_ (.A(_05790_),
    .B(net20),
    .Y(_05791_));
 sky130_fd_sc_hd__mux2_1 _12632_ (.A0(_05081_),
    .A1(_05317_),
    .S(_05788_),
    .X(_05792_));
 sky130_fd_sc_hd__a22o_1 _12633_ (.A1(net20),
    .A2(_05789_),
    .B1(_05791_),
    .B2(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__and4b_1 _12634_ (.A_N(net21),
    .B(_05793_),
    .C(net17),
    .D(net18),
    .X(_05794_));
 sky130_fd_sc_hd__and2b_1 _12635_ (.A_N(net20),
    .B(net21),
    .X(_05795_));
 sky130_fd_sc_hd__inv_2 _12636_ (.A(net18),
    .Y(_05796_));
 sky130_fd_sc_hd__nor2_1 _12637_ (.A(net19),
    .B(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__nor2_2 _12638_ (.A(net17),
    .B(net16),
    .Y(_05798_));
 sky130_fd_sc_hd__inv_2 _12639_ (.A(net17),
    .Y(_05799_));
 sky130_fd_sc_hd__and2_1 _12640_ (.A(_05799_),
    .B(net16),
    .X(_05800_));
 sky130_fd_sc_hd__a22o_1 _12641_ (.A1(_05079_),
    .A2(_05798_),
    .B1(_05800_),
    .B2(net73),
    .X(_05801_));
 sky130_fd_sc_hd__and2_1 _12642_ (.A(net17),
    .B(net16),
    .X(_05802_));
 sky130_fd_sc_hd__nor2_1 _12643_ (.A(_05799_),
    .B(_05788_),
    .Y(_05803_));
 sky130_fd_sc_hd__a22o_1 _12644_ (.A1(_05077_),
    .A2(_05802_),
    .B1(_05803_),
    .B2(net44),
    .X(_05804_));
 sky130_fd_sc_hd__nor2_1 _12645_ (.A(net19),
    .B(net18),
    .Y(_05805_));
 sky130_fd_sc_hd__a22o_1 _12646_ (.A1(_05797_),
    .A2(_05801_),
    .B1(_05804_),
    .B2(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__nor2_1 _12647_ (.A(net21),
    .B(net20),
    .Y(_05807_));
 sky130_fd_sc_hd__a41o_1 _12648_ (.A1(_05698_),
    .A2(_05802_),
    .A3(_05807_),
    .A4(_05797_),
    .B1(_05795_),
    .X(_05808_));
 sky130_fd_sc_hd__a22o_1 _12649_ (.A1(net53),
    .A2(_05798_),
    .B1(_05800_),
    .B2(net40),
    .X(_05809_));
 sky130_fd_sc_hd__a22o_1 _12650_ (.A1(_04704_),
    .A2(_05802_),
    .B1(_05803_),
    .B2(net41),
    .X(_05810_));
 sky130_fd_sc_hd__or3_1 _12651_ (.A(_05790_),
    .B(_05809_),
    .C(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__a221o_1 _12652_ (.A1(net43),
    .A2(_05798_),
    .B1(_05800_),
    .B2(net46),
    .C1(net19),
    .X(_05812_));
 sky130_fd_sc_hd__a21o_1 _12653_ (.A1(_05698_),
    .A2(_05807_),
    .B1(net52),
    .X(_05813_));
 sky130_fd_sc_hd__a22o_1 _12654_ (.A1(net51),
    .A2(_05803_),
    .B1(_05813_),
    .B2(_05802_),
    .X(_05814_));
 sky130_fd_sc_hd__a32o_1 _12655_ (.A1(_05796_),
    .A2(_05811_),
    .A3(_05812_),
    .B1(_05797_),
    .B2(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__a22o_1 _12656_ (.A1(net55),
    .A2(_05800_),
    .B1(_05803_),
    .B2(net57),
    .X(_05816_));
 sky130_fd_sc_hd__a21o_1 _12657_ (.A1(net54),
    .A2(_05798_),
    .B1(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__a221o_2 _12658_ (.A1(_05799_),
    .A2(net49),
    .B1(_05803_),
    .B2(clknet_1_0__leaf__05762_),
    .C1(_05798_),
    .X(_05818_));
 sky130_fd_sc_hd__a21o_2 _12659_ (.A1(\gpout2.clk_div[1] ),
    .A2(_05802_),
    .B1(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__a22o_2 _12660_ (.A1(_05797_),
    .A2(_05817_),
    .B1(_05819_),
    .B2(_05805_),
    .X(_05820_));
 sky130_fd_sc_hd__a22o_2 _12661_ (.A1(_05808_),
    .A2(_05815_),
    .B1(_05820_),
    .B2(_05807_),
    .X(_05821_));
 sky130_fd_sc_hd__a21oi_1 _12662_ (.A1(net17),
    .A2(net18),
    .B1(net19),
    .Y(_05822_));
 sky130_fd_sc_hd__and3b_1 _12663_ (.A_N(_05822_),
    .B(net20),
    .C(net21),
    .X(_05823_));
 sky130_fd_sc_hd__mux2_1 _12664_ (.A0(_05186_),
    .A1(_05016_),
    .S(_05788_),
    .X(_05824_));
 sky130_fd_sc_hd__mux4_1 _12665_ (.A0(_05769_),
    .A1(_05770_),
    .A2(_05715_),
    .A3(_05716_),
    .S0(_05788_),
    .S1(net19),
    .X(_05825_));
 sky130_fd_sc_hd__mux2_1 _12666_ (.A0(_04675_),
    .A1(_05711_),
    .S(_05788_),
    .X(_05826_));
 sky130_fd_sc_hd__mux2_1 _12667_ (.A0(_04683_),
    .A1(_04671_),
    .S(_05788_),
    .X(_05827_));
 sky130_fd_sc_hd__mux4_1 _12668_ (.A0(_05824_),
    .A1(_05825_),
    .A2(_05826_),
    .A3(_05827_),
    .S0(net18),
    .S1(_05799_),
    .X(_05828_));
 sky130_fd_sc_hd__mux4_1 _12669_ (.A0(_04484_),
    .A1(_04452_),
    .A2(_04458_),
    .A3(_04014_),
    .S0(_05788_),
    .S1(net17),
    .X(_05829_));
 sky130_fd_sc_hd__or2_1 _12670_ (.A(net18),
    .B(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__mux2_1 _12671_ (.A0(_04017_),
    .A1(_04018_),
    .S(_05788_),
    .X(_05831_));
 sky130_fd_sc_hd__mux4_1 _12672_ (.A0(_04010_),
    .A1(_04584_),
    .A2(_04587_),
    .A3(_04482_),
    .S0(_05788_),
    .S1(net17),
    .X(_05832_));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(_05831_),
    .A1(_05832_),
    .S(net19),
    .X(_05833_));
 sky130_fd_sc_hd__a22o_1 _12674_ (.A1(net18),
    .A2(_05791_),
    .B1(_05822_),
    .B2(net20),
    .X(_05834_));
 sky130_fd_sc_hd__o211a_1 _12675_ (.A1(_05796_),
    .A2(_05833_),
    .B1(_05834_),
    .C1(net21),
    .X(_05835_));
 sky130_fd_sc_hd__a22o_1 _12676_ (.A1(_05823_),
    .A2(_05828_),
    .B1(_05830_),
    .B2(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__a211o_2 _12677_ (.A1(_05795_),
    .A2(_05806_),
    .B1(_05821_),
    .C1(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__and4b_1 _12678_ (.A_N(_05081_),
    .B(_05798_),
    .C(_05807_),
    .D(_05805_),
    .X(_05838_));
 sky130_fd_sc_hd__o21ba_2 _12679_ (.A1(_05794_),
    .A2(_05837_),
    .B1_N(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__mux2_2 _12680_ (.A0(\reg_gpout[2] ),
    .A1(clknet_1_1__leaf__05839_),
    .S(net45),
    .X(_05840_));
 sky130_fd_sc_hd__buf_1 _12681_ (.A(_05840_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 _12682_ (.A(net22),
    .X(_05841_));
 sky130_fd_sc_hd__mux4_1 _12683_ (.A0(_05399_),
    .A1(_05492_),
    .A2(_05582_),
    .A3(_05671_),
    .S0(_05841_),
    .S1(net25),
    .X(_05842_));
 sky130_fd_sc_hd__inv_2 _12684_ (.A(net26),
    .Y(_05843_));
 sky130_fd_sc_hd__and2_1 _12685_ (.A(net25),
    .B(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__mux2_1 _12686_ (.A0(_05081_),
    .A1(_05317_),
    .S(_05841_),
    .X(_05845_));
 sky130_fd_sc_hd__a22o_1 _12687_ (.A1(net26),
    .A2(_05842_),
    .B1(_05844_),
    .B2(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__and4b_1 _12688_ (.A_N(net27),
    .B(_05846_),
    .C(net23),
    .D(net24),
    .X(_05847_));
 sky130_fd_sc_hd__nor2_1 _12689_ (.A(net26),
    .B(net27),
    .Y(_05848_));
 sky130_fd_sc_hd__and2b_1 _12690_ (.A_N(net25),
    .B(net24),
    .X(_05849_));
 sky130_fd_sc_hd__inv_2 _12691_ (.A(net23),
    .Y(_05850_));
 sky130_fd_sc_hd__and2_1 _12692_ (.A(_05850_),
    .B(_05841_),
    .X(_05851_));
 sky130_fd_sc_hd__nor2_2 _12693_ (.A(_05850_),
    .B(net22),
    .Y(_05852_));
 sky130_fd_sc_hd__nor2_2 _12694_ (.A(net23),
    .B(_05841_),
    .Y(_05853_));
 sky130_fd_sc_hd__and2_1 _12695_ (.A(net54),
    .B(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__a221o_1 _12696_ (.A1(net55),
    .A2(_05851_),
    .B1(_05852_),
    .B2(net57),
    .C1(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__and2_1 _12697_ (.A(net23),
    .B(net22),
    .X(_05856_));
 sky130_fd_sc_hd__a221o_2 _12698_ (.A1(net48),
    .A2(_05850_),
    .B1(_05852_),
    .B2(clknet_1_0__leaf__05762_),
    .C1(_05853_),
    .X(_05857_));
 sky130_fd_sc_hd__a21o_2 _12699_ (.A1(\gpout3.clk_div[1] ),
    .A2(_05856_),
    .B1(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__nor2_1 _12700_ (.A(net25),
    .B(net24),
    .Y(_05859_));
 sky130_fd_sc_hd__a22o_2 _12701_ (.A1(_05849_),
    .A2(_05855_),
    .B1(_05858_),
    .B2(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__a21o_1 _12702_ (.A1(_05698_),
    .A2(_05848_),
    .B1(net52),
    .X(_05861_));
 sky130_fd_sc_hd__a22o_1 _12703_ (.A1(net51),
    .A2(_05852_),
    .B1(_05861_),
    .B2(_05856_),
    .X(_05862_));
 sky130_fd_sc_hd__nand2_1 _12704_ (.A(_05862_),
    .B(_05849_),
    .Y(_05863_));
 sky130_fd_sc_hd__a22o_1 _12705_ (.A1(_04704_),
    .A2(_05856_),
    .B1(_05852_),
    .B2(net41),
    .X(_05864_));
 sky130_fd_sc_hd__a221o_1 _12706_ (.A1(net40),
    .A2(_05851_),
    .B1(_05853_),
    .B2(net53),
    .C1(_05864_),
    .X(_05865_));
 sky130_fd_sc_hd__inv_2 _12707_ (.A(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__a221oi_1 _12708_ (.A1(net46),
    .A2(_05851_),
    .B1(_05853_),
    .B2(net43),
    .C1(net25),
    .Y(_05867_));
 sky130_fd_sc_hd__a211o_1 _12709_ (.A1(net25),
    .A2(_05866_),
    .B1(_05867_),
    .C1(net24),
    .X(_05868_));
 sky130_fd_sc_hd__and4_1 _12710_ (.A(_05698_),
    .B(_05856_),
    .C(_05848_),
    .D(_05849_),
    .X(_05869_));
 sky130_fd_sc_hd__a21oi_1 _12711_ (.A1(_05843_),
    .A2(net27),
    .B1(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__a21oi_1 _12712_ (.A1(_05863_),
    .A2(_05868_),
    .B1(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__a21oi_1 _12713_ (.A1(net23),
    .A2(net24),
    .B1(net25),
    .Y(_05872_));
 sky130_fd_sc_hd__nor2_1 _12714_ (.A(_05843_),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(_05186_),
    .A1(_05016_),
    .S(_05841_),
    .X(_05874_));
 sky130_fd_sc_hd__mux4_1 _12716_ (.A0(\gpout0.vpos[0] ),
    .A1(_05770_),
    .A2(_05715_),
    .A3(_05716_),
    .S0(_05841_),
    .S1(net25),
    .X(_05875_));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(_04675_),
    .A1(_05711_),
    .S(_05841_),
    .X(_05876_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(_04683_),
    .A1(_04671_),
    .S(_05841_),
    .X(_05877_));
 sky130_fd_sc_hd__mux4_1 _12719_ (.A0(_05874_),
    .A1(_05875_),
    .A2(_05876_),
    .A3(_05877_),
    .S0(net24),
    .S1(_05850_),
    .X(_05878_));
 sky130_fd_sc_hd__mux4_1 _12720_ (.A0(_04484_),
    .A1(_04452_),
    .A2(_04458_),
    .A3(_04014_),
    .S0(_05841_),
    .S1(net23),
    .X(_05879_));
 sky130_fd_sc_hd__mux2_1 _12721_ (.A0(_04017_),
    .A1(_04018_),
    .S(_05841_),
    .X(_05880_));
 sky130_fd_sc_hd__mux4_1 _12722_ (.A0(_04010_),
    .A1(_04584_),
    .A2(\gpout0.hpos[2] ),
    .A3(_04482_),
    .S0(net22),
    .S1(net23),
    .X(_05881_));
 sky130_fd_sc_hd__mux2_1 _12723_ (.A0(_05880_),
    .A1(_05881_),
    .S(net25),
    .X(_05882_));
 sky130_fd_sc_hd__or2b_1 _12724_ (.A(_05882_),
    .B_N(net24),
    .X(_05883_));
 sky130_fd_sc_hd__a22o_1 _12725_ (.A1(net24),
    .A2(_05844_),
    .B1(_05872_),
    .B2(net26),
    .X(_05884_));
 sky130_fd_sc_hd__o2111a_1 _12726_ (.A1(net24),
    .A2(_05879_),
    .B1(_05883_),
    .C1(net27),
    .D1(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__a31o_1 _12727_ (.A1(net27),
    .A2(_05873_),
    .A3(_05878_),
    .B1(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__a211o_2 _12728_ (.A1(_05848_),
    .A2(_05860_),
    .B1(_05871_),
    .C1(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__a22o_1 _12729_ (.A1(net73),
    .A2(_05851_),
    .B1(_05853_),
    .B2(_05079_),
    .X(_05888_));
 sky130_fd_sc_hd__a22o_1 _12730_ (.A1(_05077_),
    .A2(_05856_),
    .B1(_05852_),
    .B2(net44),
    .X(_05889_));
 sky130_fd_sc_hd__a22o_1 _12731_ (.A1(_05849_),
    .A2(_05888_),
    .B1(_05889_),
    .B2(_05859_),
    .X(_05890_));
 sky130_fd_sc_hd__and3_1 _12732_ (.A(_05843_),
    .B(net27),
    .C(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__nand3_1 _12733_ (.A(_05853_),
    .B(_05848_),
    .C(_05859_),
    .Y(_05892_));
 sky130_fd_sc_hd__o32a_2 _12734_ (.A1(_05847_),
    .A2(_05887_),
    .A3(_05891_),
    .B1(_05892_),
    .B2(_05317_),
    .X(_05893_));
 sky130_fd_sc_hd__mux2_2 _12735_ (.A0(\reg_gpout[3] ),
    .A1(clknet_1_0__leaf__05893_),
    .S(net45),
    .X(_05894_));
 sky130_fd_sc_hd__buf_1 _12736_ (.A(_05894_),
    .X(net61));
 sky130_fd_sc_hd__a21oi_1 _12737_ (.A1(net29),
    .A2(net30),
    .B1(net31),
    .Y(_05895_));
 sky130_fd_sc_hd__and3b_1 _12738_ (.A_N(_05895_),
    .B(net33),
    .C(net32),
    .X(_05896_));
 sky130_fd_sc_hd__clkbuf_4 _12739_ (.A(net28),
    .X(_05897_));
 sky130_fd_sc_hd__mux2_1 _12740_ (.A0(_04675_),
    .A1(_05711_),
    .S(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(_04683_),
    .A1(_04671_),
    .S(_05897_),
    .X(_05899_));
 sky130_fd_sc_hd__mux2_1 _12742_ (.A0(_05186_),
    .A1(_05016_),
    .S(_05897_),
    .X(_05900_));
 sky130_fd_sc_hd__mux4_1 _12743_ (.A0(_05769_),
    .A1(_05770_),
    .A2(_05715_),
    .A3(_05716_),
    .S0(_05897_),
    .S1(net31),
    .X(_05901_));
 sky130_fd_sc_hd__mux4_1 _12744_ (.A0(_05898_),
    .A1(_05899_),
    .A2(_05900_),
    .A3(_05901_),
    .S0(net30),
    .S1(net29),
    .X(_05902_));
 sky130_fd_sc_hd__mux4_1 _12745_ (.A0(_04484_),
    .A1(_04452_),
    .A2(_04458_),
    .A3(_04014_),
    .S0(_05897_),
    .S1(net29),
    .X(_05903_));
 sky130_fd_sc_hd__or2_1 _12746_ (.A(net30),
    .B(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__inv_2 _12747_ (.A(net30),
    .Y(_05905_));
 sky130_fd_sc_hd__mux2_1 _12748_ (.A0(_04017_),
    .A1(_04018_),
    .S(_05897_),
    .X(_05906_));
 sky130_fd_sc_hd__mux4_1 _12749_ (.A0(_04010_),
    .A1(_04584_),
    .A2(_04587_),
    .A3(_04482_),
    .S0(_05897_),
    .S1(net29),
    .X(_05907_));
 sky130_fd_sc_hd__mux2_1 _12750_ (.A0(_05906_),
    .A1(_05907_),
    .S(net31),
    .X(_05908_));
 sky130_fd_sc_hd__and2b_1 _12751_ (.A_N(net32),
    .B(net31),
    .X(_05909_));
 sky130_fd_sc_hd__a22o_1 _12752_ (.A1(net30),
    .A2(_05909_),
    .B1(_05895_),
    .B2(net32),
    .X(_05910_));
 sky130_fd_sc_hd__o211a_1 _12753_ (.A1(_05905_),
    .A2(_05908_),
    .B1(_05910_),
    .C1(net33),
    .X(_05911_));
 sky130_fd_sc_hd__a22o_1 _12754_ (.A1(_05896_),
    .A2(_05902_),
    .B1(_05904_),
    .B2(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__and2_1 _12755_ (.A(net29),
    .B(net28),
    .X(_05913_));
 sky130_fd_sc_hd__nor2_1 _12756_ (.A(net32),
    .B(net33),
    .Y(_05914_));
 sky130_fd_sc_hd__nor2_1 _12757_ (.A(net31),
    .B(_05905_),
    .Y(_05915_));
 sky130_fd_sc_hd__and2b_1 _12758_ (.A_N(net32),
    .B(net33),
    .X(_05916_));
 sky130_fd_sc_hd__a41o_1 _12759_ (.A1(_05698_),
    .A2(_05913_),
    .A3(_05914_),
    .A4(_05915_),
    .B1(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__and2b_1 _12760_ (.A_N(net28),
    .B(net29),
    .X(_05918_));
 sky130_fd_sc_hd__a21o_1 _12761_ (.A1(_05698_),
    .A2(_05914_),
    .B1(net52),
    .X(_05919_));
 sky130_fd_sc_hd__a22o_1 _12762_ (.A1(net51),
    .A2(_05918_),
    .B1(_05913_),
    .B2(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__nor2_1 _12763_ (.A(net29),
    .B(net28),
    .Y(_05921_));
 sky130_fd_sc_hd__and2b_1 _12764_ (.A_N(net29),
    .B(net28),
    .X(_05922_));
 sky130_fd_sc_hd__a22o_1 _12765_ (.A1(net43),
    .A2(_05921_),
    .B1(_05922_),
    .B2(net46),
    .X(_05923_));
 sky130_fd_sc_hd__a22o_1 _12766_ (.A1(net41),
    .A2(_05918_),
    .B1(_05913_),
    .B2(_04704_),
    .X(_05924_));
 sky130_fd_sc_hd__a221o_1 _12767_ (.A1(net53),
    .A2(_05921_),
    .B1(_05922_),
    .B2(net40),
    .C1(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__mux2_1 _12768_ (.A0(_05923_),
    .A1(_05925_),
    .S(net31),
    .X(_05926_));
 sky130_fd_sc_hd__a22o_1 _12769_ (.A1(_05920_),
    .A2(_05915_),
    .B1(_05926_),
    .B2(_05905_),
    .X(_05927_));
 sky130_fd_sc_hd__a22o_1 _12770_ (.A1(net54),
    .A2(_05921_),
    .B1(_05922_),
    .B2(net55),
    .X(_05928_));
 sky130_fd_sc_hd__a21o_1 _12771_ (.A1(net57),
    .A2(_05918_),
    .B1(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__a21oi_1 _12772_ (.A1(_04672_),
    .A2(_05897_),
    .B1(net29),
    .Y(_05930_));
 sky130_fd_sc_hd__a221o_2 _12773_ (.A1(clknet_1_0__leaf__05762_),
    .A2(_05918_),
    .B1(_05913_),
    .B2(\gpout4.clk_div[1] ),
    .C1(_05930_),
    .X(_05931_));
 sky130_fd_sc_hd__nor2_1 _12774_ (.A(net31),
    .B(net30),
    .Y(_05932_));
 sky130_fd_sc_hd__a22o_2 _12775_ (.A1(_05915_),
    .A2(_05929_),
    .B1(_05931_),
    .B2(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__a22o_2 _12776_ (.A1(_05917_),
    .A2(_05927_),
    .B1(_05933_),
    .B2(_05914_),
    .X(_05934_));
 sky130_fd_sc_hd__mux4_1 _12777_ (.A0(_05399_),
    .A1(_05492_),
    .A2(_05582_),
    .A3(_05671_),
    .S0(_05897_),
    .S1(net31),
    .X(_05935_));
 sky130_fd_sc_hd__mux2_1 _12778_ (.A0(_05081_),
    .A1(_05317_),
    .S(_05897_),
    .X(_05936_));
 sky130_fd_sc_hd__a22o_1 _12779_ (.A1(net32),
    .A2(_05935_),
    .B1(_05909_),
    .B2(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__and3b_1 _12780_ (.A_N(net33),
    .B(net30),
    .C(net29),
    .X(_05938_));
 sky130_fd_sc_hd__a22o_1 _12781_ (.A1(_05079_),
    .A2(_05921_),
    .B1(_05922_),
    .B2(net73),
    .X(_05939_));
 sky130_fd_sc_hd__a22o_1 _12782_ (.A1(net44),
    .A2(_05918_),
    .B1(_05913_),
    .B2(_05077_),
    .X(_05940_));
 sky130_fd_sc_hd__a22o_1 _12783_ (.A1(_05915_),
    .A2(_05939_),
    .B1(_05940_),
    .B2(_05932_),
    .X(_05941_));
 sky130_fd_sc_hd__a22o_1 _12784_ (.A1(_05937_),
    .A2(_05938_),
    .B1(_05916_),
    .B2(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__nand4b_1 _12785_ (.A_N(_05582_),
    .B(_05921_),
    .C(_05914_),
    .D(_05932_),
    .Y(_05943_));
 sky130_fd_sc_hd__o31a_2 _12786_ (.A1(_05912_),
    .A2(_05934_),
    .A3(_05942_),
    .B1(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__mux2_2 _12787_ (.A0(\reg_gpout[4] ),
    .A1(clknet_1_1__leaf__05944_),
    .S(net45),
    .X(_05945_));
 sky130_fd_sc_hd__buf_1 _12788_ (.A(_05945_),
    .X(net62));
 sky130_fd_sc_hd__buf_2 _12789_ (.A(net35),
    .X(_05946_));
 sky130_fd_sc_hd__clkbuf_4 _12790_ (.A(net34),
    .X(_05947_));
 sky130_fd_sc_hd__or4_1 _12791_ (.A(_05946_),
    .B(_05947_),
    .C(net38),
    .D(net39),
    .X(_05948_));
 sky130_fd_sc_hd__inv_2 _12792_ (.A(net39),
    .Y(_05949_));
 sky130_fd_sc_hd__mux4_1 _12793_ (.A0(_05399_),
    .A1(_05492_),
    .A2(_05582_),
    .A3(_05671_),
    .S0(_05947_),
    .S1(net37),
    .X(_05950_));
 sky130_fd_sc_hd__inv_2 _12794_ (.A(net37),
    .Y(_05951_));
 sky130_fd_sc_hd__nor2_1 _12795_ (.A(_05951_),
    .B(net38),
    .Y(_05952_));
 sky130_fd_sc_hd__mux2_1 _12796_ (.A0(_05081_),
    .A1(_05317_),
    .S(_05947_),
    .X(_05953_));
 sky130_fd_sc_hd__a22o_1 _12797_ (.A1(net38),
    .A2(_05950_),
    .B1(_05952_),
    .B2(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__nor2_1 _12798_ (.A(_05946_),
    .B(_05947_),
    .Y(_05955_));
 sky130_fd_sc_hd__and2b_1 _12799_ (.A_N(net34),
    .B(net35),
    .X(_05956_));
 sky130_fd_sc_hd__and2b_1 _12800_ (.A_N(net35),
    .B(net34),
    .X(_05957_));
 sky130_fd_sc_hd__and3_1 _12801_ (.A(net56),
    .B(_05946_),
    .C(_05947_),
    .X(_05958_));
 sky130_fd_sc_hd__a221o_1 _12802_ (.A1(net57),
    .A2(_05956_),
    .B1(_05957_),
    .B2(net55),
    .C1(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__inv_2 _12803_ (.A(net36),
    .Y(_05960_));
 sky130_fd_sc_hd__a211o_1 _12804_ (.A1(net54),
    .A2(_05955_),
    .B1(_05959_),
    .C1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__and2_1 _12805_ (.A(net35),
    .B(net34),
    .X(_05962_));
 sky130_fd_sc_hd__a21oi_2 _12806_ (.A1(net128),
    .A2(_05946_),
    .B1(_05947_),
    .Y(_05963_));
 sky130_fd_sc_hd__a211o_2 _12807_ (.A1(\gpout5.clk_div[1] ),
    .A2(_05962_),
    .B1(_05963_),
    .C1(net36),
    .X(_05964_));
 sky130_fd_sc_hd__nor2_1 _12808_ (.A(net38),
    .B(net39),
    .Y(_05965_));
 sky130_fd_sc_hd__a221o_1 _12809_ (.A1(net53),
    .A2(_05955_),
    .B1(_05957_),
    .B2(net40),
    .C1(_05951_),
    .X(_05966_));
 sky130_fd_sc_hd__a22o_1 _12810_ (.A1(net52),
    .A2(_05962_),
    .B1(_05956_),
    .B2(net51),
    .X(_05967_));
 sky130_fd_sc_hd__a221o_1 _12811_ (.A1(_05079_),
    .A2(_05955_),
    .B1(_05957_),
    .B2(net73),
    .C1(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__a22o_1 _12812_ (.A1(_05960_),
    .A2(_05966_),
    .B1(_05968_),
    .B2(_05951_),
    .X(_05969_));
 sky130_fd_sc_hd__mux4_1 _12813_ (.A0(net43),
    .A1(net46),
    .A2(net44),
    .A3(_05077_),
    .S0(_05947_),
    .S1(_05946_),
    .X(_05970_));
 sky130_fd_sc_hd__or3_1 _12814_ (.A(net37),
    .B(net36),
    .C(_05970_),
    .X(_05971_));
 sky130_fd_sc_hd__and3b_1 _12815_ (.A_N(net38),
    .B(_05969_),
    .C(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__and3_1 _12816_ (.A(_04482_),
    .B(net35),
    .C(net34),
    .X(_05973_));
 sky130_fd_sc_hd__a221o_1 _12817_ (.A1(_04010_),
    .A2(_05955_),
    .B1(_05957_),
    .B2(_04584_),
    .C1(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__a211o_1 _12818_ (.A1(_04587_),
    .A2(_05956_),
    .B1(_05974_),
    .C1(_05960_),
    .X(_05975_));
 sky130_fd_sc_hd__a221o_1 _12819_ (.A1(_04704_),
    .A2(_05962_),
    .B1(_05956_),
    .B2(net41),
    .C1(net36),
    .X(_05976_));
 sky130_fd_sc_hd__and3_1 _12820_ (.A(_05952_),
    .B(_05975_),
    .C(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__mux4_1 _12821_ (.A0(_04675_),
    .A1(_04678_),
    .A2(_04683_),
    .A3(_04671_),
    .S0(_05947_),
    .S1(net36),
    .X(_05978_));
 sky130_fd_sc_hd__mux4_1 _12822_ (.A0(_05186_),
    .A1(_05016_),
    .A2(\gpout0.vpos[8] ),
    .A3(\gpout0.vpos[9] ),
    .S0(_05947_),
    .S1(net36),
    .X(_05979_));
 sky130_fd_sc_hd__mux2_1 _12823_ (.A0(_05978_),
    .A1(_05979_),
    .S(_05946_),
    .X(_05980_));
 sky130_fd_sc_hd__mux2_1 _12824_ (.A0(_04458_),
    .A1(_04014_),
    .S(_05947_),
    .X(_05981_));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(\gpout0.vpos[0] ),
    .A1(\gpout0.vpos[1] ),
    .S(net34),
    .X(_05982_));
 sky130_fd_sc_hd__a31o_1 _12826_ (.A1(_05946_),
    .A2(net36),
    .A3(_05982_),
    .B1(net37),
    .X(_05983_));
 sky130_fd_sc_hd__mux4_1 _12827_ (.A0(_04484_),
    .A1(_04017_),
    .A2(_04452_),
    .A3(_04018_),
    .S0(net36),
    .S1(net34),
    .X(_05984_));
 sky130_fd_sc_hd__and2b_1 _12828_ (.A_N(_05946_),
    .B(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__a311o_1 _12829_ (.A1(_05946_),
    .A2(_05960_),
    .A3(_05981_),
    .B1(_05983_),
    .C1(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__o211a_1 _12830_ (.A1(_05951_),
    .A2(_05980_),
    .B1(_05986_),
    .C1(net38),
    .X(_05987_));
 sky130_fd_sc_hd__o31a_1 _12831_ (.A1(_05972_),
    .A2(_05977_),
    .A3(_05987_),
    .B1(net39),
    .X(_05988_));
 sky130_fd_sc_hd__a41o_2 _12832_ (.A1(_05951_),
    .A2(_05961_),
    .A3(_05964_),
    .A4(_05965_),
    .B1(_05988_),
    .X(_05989_));
 sky130_fd_sc_hd__a41o_2 _12833_ (.A1(_05946_),
    .A2(net36),
    .A3(_05949_),
    .A4(_05954_),
    .B1(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__o41a_2 _12834_ (.A1(net37),
    .A2(net36),
    .A3(_05671_),
    .A4(_05948_),
    .B1(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__mux2_2 _12835_ (.A0(\reg_gpout[5] ),
    .A1(clknet_1_1__leaf__05991_),
    .S(net45),
    .X(_05992_));
 sky130_fd_sc_hd__buf_1 _12836_ (.A(_05992_),
    .X(net63));
 sky130_fd_sc_hd__clkinv_2 _12837_ (.A(\rbzero.map_rom.i_row[4] ),
    .Y(_05993_));
 sky130_fd_sc_hd__inv_2 _12838_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .Y(_05994_));
 sky130_fd_sc_hd__nand2_1 _12839_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_05995_));
 sky130_fd_sc_hd__or2_1 _12840_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_05996_));
 sky130_fd_sc_hd__nand3_1 _12841_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .C(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__and2_1 _12842_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_05998_));
 sky130_fd_sc_hd__or2_1 _12843_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_05999_));
 sky130_fd_sc_hd__or2b_1 _12844_ (.A(_05998_),
    .B_N(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__nand2_1 _12845_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06001_));
 sky130_fd_sc_hd__or2_1 _12846_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_06002_));
 sky130_fd_sc_hd__nand2_1 _12847_ (.A(_06001_),
    .B(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__or2_1 _12848_ (.A(_06000_),
    .B(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__nand2_1 _12849_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_06005_));
 sky130_fd_sc_hd__or2_1 _12850_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_06006_));
 sky130_fd_sc_hd__and2_1 _12851_ (.A(_06005_),
    .B(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__nor2_1 _12852_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06008_));
 sky130_fd_sc_hd__and2_1 _12853_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_06009_));
 sky130_fd_sc_hd__nor2_1 _12854_ (.A(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2_1 _12855_ (.A(_06007_),
    .B(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__or2_1 _12856_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_06012_));
 sky130_fd_sc_hd__or2_1 _12857_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06013_));
 sky130_fd_sc_hd__xor2_1 _12858_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06014_));
 sky130_fd_sc_hd__and2_1 _12859_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06015_));
 sky130_fd_sc_hd__a31o_1 _12860_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_06014_),
    .B1(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__and2_1 _12861_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06017_));
 sky130_fd_sc_hd__a221o_1 _12862_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_06013_),
    .B2(_06016_),
    .C1(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__or4bb_1 _12863_ (.A(_06004_),
    .B(_06011_),
    .C_N(_06012_),
    .D_N(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06020_));
 sky130_fd_sc_hd__a21o_1 _12865_ (.A1(_06005_),
    .A2(_06020_),
    .B1(_06008_),
    .X(_06021_));
 sky130_fd_sc_hd__a31o_1 _12866_ (.A1(\rbzero.debug_overlay.facingY[-3] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .A3(_05999_),
    .B1(_05998_),
    .X(_06022_));
 sky130_fd_sc_hd__o21ba_1 _12867_ (.A1(_06004_),
    .A2(_06021_),
    .B1_N(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__nand2_1 _12868_ (.A(_05996_),
    .B(_05995_),
    .Y(_06024_));
 sky130_fd_sc_hd__nand2_1 _12869_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_06025_));
 sky130_fd_sc_hd__or2_1 _12870_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_06026_));
 sky130_fd_sc_hd__nand2_1 _12871_ (.A(_06025_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__a211o_1 _12872_ (.A1(_06019_),
    .A2(_06023_),
    .B1(_06024_),
    .C1(_06027_),
    .X(_06028_));
 sky130_fd_sc_hd__nand2_1 _12873_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06029_));
 sky130_fd_sc_hd__nor2_1 _12874_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06030_));
 sky130_fd_sc_hd__a41o_1 _12875_ (.A1(_05995_),
    .A2(_05997_),
    .A3(_06028_),
    .A4(_06029_),
    .B1(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__or2_1 _12876_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_06032_));
 sky130_fd_sc_hd__nand2_1 _12877_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_06033_));
 sky130_fd_sc_hd__nand2_1 _12878_ (.A(_06032_),
    .B(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__xor2_2 _12879_ (.A(_06031_),
    .B(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__and2b_1 _12880_ (.A_N(_06030_),
    .B(_06029_),
    .X(_06036_));
 sky130_fd_sc_hd__a31oi_1 _12881_ (.A1(_05995_),
    .A2(_05997_),
    .A3(_06028_),
    .B1(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__and4_1 _12882_ (.A(_05995_),
    .B(_05997_),
    .C(_06028_),
    .D(_06036_),
    .X(_06038_));
 sky130_fd_sc_hd__or2_1 _12883_ (.A(_06037_),
    .B(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__nand3_1 _12884_ (.A(_06012_),
    .B(_06018_),
    .C(_06007_),
    .Y(_06040_));
 sky130_fd_sc_hd__a311o_1 _12885_ (.A1(_06005_),
    .A2(_06040_),
    .A3(_06020_),
    .B1(_06008_),
    .C1(_06003_),
    .X(_06041_));
 sky130_fd_sc_hd__a21oi_1 _12886_ (.A1(_06001_),
    .A2(_06041_),
    .B1(_06000_),
    .Y(_06042_));
 sky130_fd_sc_hd__and3_1 _12887_ (.A(_06000_),
    .B(_06001_),
    .C(_06041_),
    .X(_06043_));
 sky130_fd_sc_hd__nor2_1 _12888_ (.A(_06042_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__inv_2 _12889_ (.A(_06008_),
    .Y(_06045_));
 sky130_fd_sc_hd__a32o_1 _12890_ (.A1(_06012_),
    .A2(_06018_),
    .A3(_06007_),
    .B1(\rbzero.wall_tracer.rayAddendY[3] ),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .X(_06046_));
 sky130_fd_sc_hd__a221o_1 _12891_ (.A1(_06001_),
    .A2(_06002_),
    .B1(_06045_),
    .B2(_06046_),
    .C1(_06009_),
    .X(_06047_));
 sky130_fd_sc_hd__and2_1 _12892_ (.A(_06041_),
    .B(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__a21oi_1 _12893_ (.A1(_06019_),
    .A2(_06023_),
    .B1(_06027_),
    .Y(_06049_));
 sky130_fd_sc_hd__and3_1 _12894_ (.A(_06027_),
    .B(_06019_),
    .C(_06023_),
    .X(_06050_));
 sky130_fd_sc_hd__nor2_1 _12895_ (.A(_06049_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__xor2_2 _12896_ (.A(_06010_),
    .B(_06046_),
    .X(_06052_));
 sky130_fd_sc_hd__a21o_1 _12897_ (.A1(_06012_),
    .A2(_06018_),
    .B1(_06007_),
    .X(_06053_));
 sky130_fd_sc_hd__and2_1 _12898_ (.A(_06040_),
    .B(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__nand2_1 _12899_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_06055_));
 sky130_fd_sc_hd__nand2_1 _12900_ (.A(_06012_),
    .B(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__a21o_1 _12901_ (.A1(_06013_),
    .A2(_06016_),
    .B1(_06017_),
    .X(_06057_));
 sky130_fd_sc_hd__xnor2_1 _12902_ (.A(_06056_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__and2b_1 _12903_ (.A_N(_06017_),
    .B(_06013_),
    .X(_06059_));
 sky130_fd_sc_hd__xor2_2 _12904_ (.A(_06059_),
    .B(_06016_),
    .X(_06060_));
 sky130_fd_sc_hd__nand2_1 _12905_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_06061_));
 sky130_fd_sc_hd__xnor2_1 _12906_ (.A(_06061_),
    .B(_06014_),
    .Y(_06062_));
 sky130_fd_sc_hd__xor2_1 _12907_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_06063_));
 sky130_fd_sc_hd__or4_1 _12908_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C(_06062_),
    .D(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__or4_1 _12909_ (.A(_06054_),
    .B(_06058_),
    .C(_06060_),
    .D(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__or3_1 _12910_ (.A(_06051_),
    .B(_06052_),
    .C(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__a21o_1 _12911_ (.A1(_06019_),
    .A2(_06023_),
    .B1(_06027_),
    .X(_06067_));
 sky130_fd_sc_hd__a21o_1 _12912_ (.A1(_06025_),
    .A2(_06067_),
    .B1(_06024_),
    .X(_06068_));
 sky130_fd_sc_hd__nand3_1 _12913_ (.A(_06025_),
    .B(_06067_),
    .C(_06024_),
    .Y(_06069_));
 sky130_fd_sc_hd__nand2_1 _12914_ (.A(_06068_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__or3b_1 _12915_ (.A(_06048_),
    .B(_06066_),
    .C_N(_06070_),
    .X(_06071_));
 sky130_fd_sc_hd__inv_2 _12916_ (.A(_06033_),
    .Y(_06072_));
 sky130_fd_sc_hd__o21ai_1 _12917_ (.A1(_06072_),
    .A2(_06031_),
    .B1(_06032_),
    .Y(_06073_));
 sky130_fd_sc_hd__o41a_4 _12918_ (.A1(_06035_),
    .A2(_06039_),
    .A3(_06044_),
    .A4(_06071_),
    .B1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__buf_4 _12919_ (.A(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__buf_4 _12920_ (.A(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__a21oi_1 _12921_ (.A1(_05993_),
    .A2(_05994_),
    .B1(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__xnor2_1 _12922_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .B(_06076_),
    .Y(_06078_));
 sky130_fd_sc_hd__clkinv_2 _12923_ (.A(\rbzero.map_rom.a6 ),
    .Y(_06079_));
 sky130_fd_sc_hd__nor2_1 _12924_ (.A(_06079_),
    .B(_06076_),
    .Y(_06080_));
 sky130_fd_sc_hd__clkinv_4 _12925_ (.A(_06075_),
    .Y(_06081_));
 sky130_fd_sc_hd__nor2_1 _12926_ (.A(\rbzero.map_rom.a6 ),
    .B(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__clkinv_2 _12927_ (.A(\rbzero.map_rom.b6 ),
    .Y(_06083_));
 sky130_fd_sc_hd__inv_2 _12928_ (.A(\rbzero.map_rom.c6 ),
    .Y(_06084_));
 sky130_fd_sc_hd__nor2_1 _12929_ (.A(_06084_),
    .B(_06075_),
    .Y(_06085_));
 sky130_fd_sc_hd__buf_2 _12930_ (.A(\rbzero.map_rom.d6 ),
    .X(_06086_));
 sky130_fd_sc_hd__nor2_1 _12931_ (.A(\rbzero.map_rom.c6 ),
    .B(_06081_),
    .Y(_06087_));
 sky130_fd_sc_hd__nor2_1 _12932_ (.A(_06085_),
    .B(_06087_),
    .Y(_06088_));
 sky130_fd_sc_hd__and2_1 _12933_ (.A(_06086_),
    .B(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__xnor2_1 _12934_ (.A(\rbzero.map_rom.b6 ),
    .B(_06075_),
    .Y(_06090_));
 sky130_fd_sc_hd__o21ai_1 _12935_ (.A1(_06085_),
    .A2(_06089_),
    .B1(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__o21ai_1 _12936_ (.A1(_06083_),
    .A2(_06076_),
    .B1(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__and2b_1 _12937_ (.A_N(_06082_),
    .B(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__xnor2_1 _12938_ (.A(\rbzero.map_rom.i_row[4] ),
    .B(_06076_),
    .Y(_06094_));
 sky130_fd_sc_hd__o21a_1 _12939_ (.A1(_06080_),
    .A2(_06093_),
    .B1(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__and2_1 _12940_ (.A(_06078_),
    .B(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__xnor2_1 _12941_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_06076_),
    .Y(_06097_));
 sky130_fd_sc_hd__o21ai_1 _12942_ (.A1(_06077_),
    .A2(_06096_),
    .B1(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__or3_1 _12943_ (.A(_06097_),
    .B(_06077_),
    .C(_06096_),
    .X(_06099_));
 sky130_fd_sc_hd__or2_1 _12944_ (.A(_04465_),
    .B(_04473_),
    .X(_06100_));
 sky130_fd_sc_hd__buf_4 _12945_ (.A(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__buf_6 _12946_ (.A(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__nand2_1 _12947_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(\rbzero.wall_tracer.mapX[5] ),
    .Y(_06103_));
 sky130_fd_sc_hd__or2_1 _12948_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .B(\rbzero.wall_tracer.mapX[5] ),
    .X(_06104_));
 sky130_fd_sc_hd__buf_2 _12949_ (.A(\rbzero.map_rom.f1 ),
    .X(_06105_));
 sky130_fd_sc_hd__nand2_1 _12950_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__or2_1 _12951_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_06105_),
    .X(_06107_));
 sky130_fd_sc_hd__buf_2 _12952_ (.A(\rbzero.map_rom.f4 ),
    .X(_06108_));
 sky130_fd_sc_hd__xor2_1 _12953_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__a221o_1 _12954_ (.A1(_06103_),
    .A2(_06104_),
    .B1(_06106_),
    .B2(_06107_),
    .C1(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__or4_1 _12955_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(\rbzero.wall_tracer.mapY[9] ),
    .C(\rbzero.wall_tracer.mapY[8] ),
    .D(\rbzero.wall_tracer.mapY[10] ),
    .X(_06111_));
 sky130_fd_sc_hd__or4_1 _12956_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(\rbzero.wall_tracer.mapX[8] ),
    .C(\rbzero.wall_tracer.mapX[10] ),
    .D(\rbzero.wall_tracer.mapY[7] ),
    .X(_06112_));
 sky130_fd_sc_hd__inv_2 _12957_ (.A(\rbzero.map_rom.d6 ),
    .Y(_06113_));
 sky130_fd_sc_hd__a211o_1 _12958_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_06084_),
    .B1(\rbzero.wall_tracer.mapX[6] ),
    .C1(\rbzero.wall_tracer.mapX[7] ),
    .X(_06114_));
 sky130_fd_sc_hd__a221o_1 _12959_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_06113_),
    .B1(_06079_),
    .B2(\rbzero.debug_overlay.playerY[3] ),
    .C1(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__clkinv_2 _12960_ (.A(\rbzero.map_rom.i_col[4] ),
    .Y(_06116_));
 sky130_fd_sc_hd__buf_2 _12961_ (.A(\rbzero.map_rom.f2 ),
    .X(_06117_));
 sky130_fd_sc_hd__o22a_1 _12962_ (.A1(_05000_),
    .A2(_06117_),
    .B1(_06113_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .X(_06118_));
 sky130_fd_sc_hd__o21ai_1 _12963_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_06116_),
    .B1(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__a22o_1 _12964_ (.A1(_05000_),
    .A2(\rbzero.map_rom.f2 ),
    .B1(_05994_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .X(_06120_));
 sky130_fd_sc_hd__a221o_1 _12965_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_06116_),
    .B1(_06083_),
    .B2(\rbzero.debug_overlay.playerY[2] ),
    .C1(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__clkinv_2 _12966_ (.A(\rbzero.map_rom.f3 ),
    .Y(_06122_));
 sky130_fd_sc_hd__inv_2 _12967_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .Y(_06123_));
 sky130_fd_sc_hd__a2bb2o_1 _12968_ (.A1_N(\rbzero.debug_overlay.playerY[1] ),
    .A2_N(_06084_),
    .B1(_05993_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .X(_06124_));
 sky130_fd_sc_hd__a221o_1 _12969_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_06122_),
    .B1(\rbzero.wall_tracer.mapY[5] ),
    .B2(_06123_),
    .C1(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__clkbuf_4 _12970_ (.A(\rbzero.map_rom.f3 ),
    .X(_06126_));
 sky130_fd_sc_hd__inv_2 _12971_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .Y(_06127_));
 sky130_fd_sc_hd__a22o_1 _12972_ (.A1(_06127_),
    .A2(\rbzero.map_rom.b6 ),
    .B1(\rbzero.map_rom.a6 ),
    .B2(_04993_),
    .X(_06128_));
 sky130_fd_sc_hd__a221o_1 _12973_ (.A1(_04998_),
    .A2(_06126_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_04997_),
    .C1(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__or4_1 _12974_ (.A(_06119_),
    .B(_06121_),
    .C(_06125_),
    .D(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__or4_1 _12975_ (.A(_06111_),
    .B(_06112_),
    .C(_06115_),
    .D(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__or4_1 _12976_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(\rbzero.wall_tracer.visualWallDist[2] ),
    .C(\rbzero.wall_tracer.visualWallDist[1] ),
    .D(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_06132_));
 sky130_fd_sc_hd__or4_1 _12977_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(\rbzero.wall_tracer.visualWallDist[-2] ),
    .C(\rbzero.wall_tracer.visualWallDist[-3] ),
    .D(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__or4_1 _12978_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(\rbzero.wall_tracer.visualWallDist[6] ),
    .C(\rbzero.wall_tracer.visualWallDist[5] ),
    .D(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_06134_));
 sky130_fd_sc_hd__inv_2 _12979_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .Y(_06135_));
 sky130_fd_sc_hd__o41a_2 _12980_ (.A1(\rbzero.wall_tracer.visualWallDist[9] ),
    .A2(\rbzero.wall_tracer.visualWallDist[8] ),
    .A3(_06133_),
    .A4(_06134_),
    .B1(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__o21ai_4 _12981_ (.A1(_06110_),
    .A2(_06131_),
    .B1(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__or2_1 _12982_ (.A(\rbzero.map_rom.d6 ),
    .B(\rbzero.map_rom.c6 ),
    .X(_06138_));
 sky130_fd_sc_hd__and4b_1 _12983_ (.A_N(_06138_),
    .B(_05993_),
    .C(_06079_),
    .D(_06083_),
    .X(_06139_));
 sky130_fd_sc_hd__xor2_1 _12984_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(\rbzero.map_rom.b6 ),
    .X(_06140_));
 sky130_fd_sc_hd__a221o_1 _12985_ (.A1(\rbzero.map_overlay.i_mapdy[1] ),
    .A2(_06084_),
    .B1(_05993_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__xnor2_1 _12986_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_rom.a6 ),
    .Y(_06142_));
 sky130_fd_sc_hd__o221a_1 _12987_ (.A1(_05022_),
    .A2(_06086_),
    .B1(_05993_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__o221a_1 _12988_ (.A1(\rbzero.map_overlay.i_mapdy[0] ),
    .A2(_06113_),
    .B1(_06084_),
    .B2(\rbzero.map_overlay.i_mapdy[1] ),
    .C1(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__nor4b_4 _12989_ (.A(_06137_),
    .B(_06139_),
    .C(_06141_),
    .D_N(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__clkinv_2 _12990_ (.A(_06117_),
    .Y(_06146_));
 sky130_fd_sc_hd__a22o_1 _12991_ (.A1(\rbzero.map_overlay.i_mapdx[2] ),
    .A2(_06146_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .B2(_05026_),
    .X(_06147_));
 sky130_fd_sc_hd__nor2_1 _12992_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06108_),
    .Y(_06148_));
 sky130_fd_sc_hd__and2_1 _12993_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06108_),
    .X(_06149_));
 sky130_fd_sc_hd__xnor2_1 _12994_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_06105_),
    .Y(_06150_));
 sky130_fd_sc_hd__o221a_1 _12995_ (.A1(\rbzero.map_overlay.i_mapdx[1] ),
    .A2(_06122_),
    .B1(_06146_),
    .B2(\rbzero.map_overlay.i_mapdx[2] ),
    .C1(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__o221a_1 _12996_ (.A1(_05027_),
    .A2(_06126_),
    .B1(_06148_),
    .B2(_06149_),
    .C1(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__a21o_1 _12997_ (.A1(_05026_),
    .A2(_05031_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .X(_06153_));
 sky130_fd_sc_hd__and4bb_1 _12998_ (.A_N(_06137_),
    .B_N(_06147_),
    .C(_06152_),
    .D(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__or2_2 _12999_ (.A(_06145_),
    .B(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__nor2_2 _13000_ (.A(_06101_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__and2b_1 _13001_ (.A_N(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .X(_06157_));
 sky130_fd_sc_hd__nand2_4 _13002_ (.A(\rbzero.trace_state[1] ),
    .B(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__nor2_1 _13003_ (.A(\rbzero.trace_state[0] ),
    .B(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__buf_4 _13004_ (.A(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__buf_4 _13005_ (.A(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__buf_4 _13006_ (.A(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__buf_6 _13007_ (.A(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__inv_2 _13008_ (.A(\rbzero.map_rom.f4 ),
    .Y(_06164_));
 sky130_fd_sc_hd__nand2_1 _13009_ (.A(_06086_),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06165_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(_06138_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__a22o_1 _13011_ (.A1(_06164_),
    .A2(_06113_),
    .B1(_06166_),
    .B2(_06126_),
    .X(_06167_));
 sky130_fd_sc_hd__and3_1 _13012_ (.A(\rbzero.map_rom.b6 ),
    .B(\rbzero.map_rom.a6 ),
    .C(\rbzero.map_rom.i_row[4] ),
    .X(_06168_));
 sky130_fd_sc_hd__and3_1 _13013_ (.A(_06117_),
    .B(\rbzero.map_rom.f1 ),
    .C(\rbzero.map_rom.i_col[4] ),
    .X(_06169_));
 sky130_fd_sc_hd__a31o_1 _13014_ (.A1(\rbzero.map_rom.f4 ),
    .A2(_06126_),
    .A3(_06169_),
    .B1(_06139_),
    .X(_06170_));
 sky130_fd_sc_hd__a31o_1 _13015_ (.A1(_06086_),
    .A2(\rbzero.map_rom.c6 ),
    .A3(_06168_),
    .B1(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__a31o_1 _13016_ (.A1(_06117_),
    .A2(\rbzero.map_rom.b6 ),
    .A3(_06167_),
    .B1(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__or2_1 _13017_ (.A(_06126_),
    .B(\rbzero.map_rom.i_col[4] ),
    .X(_06173_));
 sky130_fd_sc_hd__or4_1 _13018_ (.A(_06108_),
    .B(_06117_),
    .C(_06105_),
    .D(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__a22o_1 _13019_ (.A1(_06164_),
    .A2(_06113_),
    .B1(\rbzero.map_rom.b6 ),
    .B2(_06117_),
    .X(_06175_));
 sky130_fd_sc_hd__a2111o_1 _13020_ (.A1(_06146_),
    .A2(_06083_),
    .B1(\rbzero.map_rom.a6 ),
    .C1(_06175_),
    .D1(_06105_),
    .X(_06176_));
 sky130_fd_sc_hd__a22o_1 _13021_ (.A1(_06108_),
    .A2(_06086_),
    .B1(\rbzero.map_rom.c6 ),
    .B2(_06126_),
    .X(_06177_));
 sky130_fd_sc_hd__a211o_1 _13022_ (.A1(_06122_),
    .A2(_06084_),
    .B1(_06176_),
    .C1(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__or4_1 _13023_ (.A(_06108_),
    .B(_06117_),
    .C(_06086_),
    .D(\rbzero.map_rom.b6 ),
    .X(_06179_));
 sky130_fd_sc_hd__and4b_1 _13024_ (.A_N(_06172_),
    .B(_06174_),
    .C(_06178_),
    .D(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__or4b_1 _13025_ (.A(_06084_),
    .B(\rbzero.map_rom.i_row[4] ),
    .C(_06079_),
    .D_N(_06105_),
    .X(_06181_));
 sky130_fd_sc_hd__xnor2_1 _13026_ (.A(_06117_),
    .B(\rbzero.map_rom.a6 ),
    .Y(_06182_));
 sky130_fd_sc_hd__o22ai_1 _13027_ (.A1(_06126_),
    .A2(_06086_),
    .B1(\rbzero.map_rom.c6 ),
    .B2(\rbzero.map_rom.f1 ),
    .Y(_06183_));
 sky130_fd_sc_hd__a221o_1 _13028_ (.A1(_06105_),
    .A2(\rbzero.map_rom.c6 ),
    .B1(\rbzero.map_rom.b6 ),
    .B2(\rbzero.map_rom.f4 ),
    .C1(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__a22o_1 _13029_ (.A1(_06126_),
    .A2(_06086_),
    .B1(_06083_),
    .B2(_06164_),
    .X(_06185_));
 sky130_fd_sc_hd__or3_1 _13030_ (.A(_06182_),
    .B(_06184_),
    .C(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__o31a_1 _13031_ (.A1(_06173_),
    .A2(_06179_),
    .A3(_06181_),
    .B1(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__inv_2 _13032_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .Y(_06188_));
 sky130_fd_sc_hd__a22o_1 _13033_ (.A1(\rbzero.map_overlay.i_otherx[2] ),
    .A2(_06146_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_05039_),
    .X(_06189_));
 sky130_fd_sc_hd__a221o_1 _13034_ (.A1(_06188_),
    .A2(_06108_),
    .B1(_06113_),
    .B2(\rbzero.map_overlay.i_othery[0] ),
    .C1(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__o22a_1 _13035_ (.A1(\rbzero.map_overlay.i_othery[2] ),
    .A2(_06083_),
    .B1(_06079_),
    .B2(\rbzero.map_overlay.i_othery[3] ),
    .X(_06191_));
 sky130_fd_sc_hd__o221ai_1 _13036_ (.A1(_06188_),
    .A2(\rbzero.map_rom.f4 ),
    .B1(_06084_),
    .B2(\rbzero.map_overlay.i_othery[1] ),
    .C1(_06191_),
    .Y(_06192_));
 sky130_fd_sc_hd__a2bb2o_1 _13037_ (.A1_N(\rbzero.map_overlay.i_otherx[4] ),
    .A2_N(_06116_),
    .B1(_06083_),
    .B2(\rbzero.map_overlay.i_othery[2] ),
    .X(_06193_));
 sky130_fd_sc_hd__a22o_1 _13038_ (.A1(_05050_),
    .A2(\rbzero.map_rom.f1 ),
    .B1(_06079_),
    .B2(\rbzero.map_overlay.i_othery[3] ),
    .X(_06194_));
 sky130_fd_sc_hd__a221o_1 _13039_ (.A1(_05047_),
    .A2(_06126_),
    .B1(_05993_),
    .B2(\rbzero.map_overlay.i_othery[4] ),
    .C1(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__o22a_1 _13040_ (.A1(\rbzero.map_overlay.i_otherx[2] ),
    .A2(_06146_),
    .B1(_06113_),
    .B2(\rbzero.map_overlay.i_othery[0] ),
    .X(_06196_));
 sky130_fd_sc_hd__or4b_1 _13041_ (.A(_06192_),
    .B(_06193_),
    .C(_06195_),
    .D_N(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__a2bb2o_1 _13042_ (.A1_N(_05050_),
    .A2_N(\rbzero.map_rom.f1 ),
    .B1(\rbzero.map_overlay.i_otherx[1] ),
    .B2(_06122_),
    .X(_06198_));
 sky130_fd_sc_hd__a221o_1 _13043_ (.A1(\rbzero.map_overlay.i_otherx[4] ),
    .A2(_06116_),
    .B1(_06084_),
    .B2(\rbzero.map_overlay.i_othery[1] ),
    .C1(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__or3_1 _13044_ (.A(_06190_),
    .B(_06197_),
    .C(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__a31o_2 _13045_ (.A1(_06180_),
    .A2(_06187_),
    .A3(_06200_),
    .B1(_06137_),
    .X(_06201_));
 sky130_fd_sc_hd__or3b_4 _13046_ (.A(_06145_),
    .B(_06154_),
    .C_N(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__nor2_2 _13047_ (.A(_06101_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__inv_2 _13048_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .Y(_06204_));
 sky130_fd_sc_hd__inv_2 _13049_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .Y(_06205_));
 sky130_fd_sc_hd__nand2_1 _13050_ (.A(_06205_),
    .B(\rbzero.wall_tracer.trackDistX[9] ),
    .Y(_06206_));
 sky130_fd_sc_hd__inv_2 _13051_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .Y(_06207_));
 sky130_fd_sc_hd__inv_2 _13052_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .Y(_06208_));
 sky130_fd_sc_hd__inv_2 _13053_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .Y(_06209_));
 sky130_fd_sc_hd__inv_2 _13054_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .Y(_06210_));
 sky130_fd_sc_hd__inv_2 _13055_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .Y(_06211_));
 sky130_fd_sc_hd__inv_2 _13056_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .Y(_06212_));
 sky130_fd_sc_hd__inv_2 _13057_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .Y(_06213_));
 sky130_fd_sc_hd__inv_2 _13058_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .Y(_06214_));
 sky130_fd_sc_hd__inv_2 _13059_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .Y(_06215_));
 sky130_fd_sc_hd__inv_2 _13060_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .Y(_06216_));
 sky130_fd_sc_hd__a2bb2o_1 _13061_ (.A1_N(_06216_),
    .A2_N(\rbzero.wall_tracer.trackDistY[-1] ),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_06215_),
    .X(_06217_));
 sky130_fd_sc_hd__o21ai_1 _13062_ (.A1(_06215_),
    .A2(\rbzero.wall_tracer.trackDistX[0] ),
    .B1(_06217_),
    .Y(_06218_));
 sky130_fd_sc_hd__inv_2 _13063_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .Y(_06219_));
 sky130_fd_sc_hd__inv_2 _13064_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .Y(_06220_));
 sky130_fd_sc_hd__a22o_1 _13065_ (.A1(\rbzero.wall_tracer.trackDistY[0] ),
    .A2(_06219_),
    .B1(\rbzero.wall_tracer.trackDistY[-2] ),
    .B2(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__inv_2 _13066_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .Y(_06222_));
 sky130_fd_sc_hd__inv_2 _13067_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .Y(_06223_));
 sky130_fd_sc_hd__inv_2 _13068_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .Y(_06224_));
 sky130_fd_sc_hd__inv_2 _13069_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .Y(_06225_));
 sky130_fd_sc_hd__inv_2 _13070_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .Y(_06226_));
 sky130_fd_sc_hd__inv_2 _13071_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .Y(_06227_));
 sky130_fd_sc_hd__inv_2 _13072_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .Y(_06228_));
 sky130_fd_sc_hd__inv_2 _13073_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .Y(_06229_));
 sky130_fd_sc_hd__inv_2 _13074_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .Y(_06230_));
 sky130_fd_sc_hd__o211a_1 _13075_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(_06229_),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .C1(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__a221o_1 _13076_ (.A1(\rbzero.wall_tracer.trackDistY[-9] ),
    .A2(_06228_),
    .B1(\rbzero.wall_tracer.trackDistY[-10] ),
    .B2(_06229_),
    .C1(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__o221a_1 _13077_ (.A1(\rbzero.wall_tracer.trackDistY[-8] ),
    .A2(_06227_),
    .B1(\rbzero.wall_tracer.trackDistY[-9] ),
    .B2(_06228_),
    .C1(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__a221o_1 _13078_ (.A1(_06226_),
    .A2(\rbzero.wall_tracer.trackDistY[-7] ),
    .B1(\rbzero.wall_tracer.trackDistY[-8] ),
    .B2(_06227_),
    .C1(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__o221a_1 _13079_ (.A1(\rbzero.wall_tracer.trackDistY[-6] ),
    .A2(_06225_),
    .B1(_06226_),
    .B2(\rbzero.wall_tracer.trackDistY[-7] ),
    .C1(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__a221o_1 _13080_ (.A1(\rbzero.wall_tracer.trackDistY[-5] ),
    .A2(_06224_),
    .B1(\rbzero.wall_tracer.trackDistY[-6] ),
    .B2(_06225_),
    .C1(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__o221a_1 _13081_ (.A1(\rbzero.wall_tracer.trackDistY[-4] ),
    .A2(_06223_),
    .B1(\rbzero.wall_tracer.trackDistY[-5] ),
    .B2(_06224_),
    .C1(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__a221o_1 _13082_ (.A1(_06222_),
    .A2(\rbzero.wall_tracer.trackDistY[-3] ),
    .B1(\rbzero.wall_tracer.trackDistY[-4] ),
    .B2(_06223_),
    .C1(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__o221a_1 _13083_ (.A1(\rbzero.wall_tracer.trackDistY[-2] ),
    .A2(_06220_),
    .B1(_06222_),
    .B2(\rbzero.wall_tracer.trackDistY[-3] ),
    .C1(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__a2111o_1 _13084_ (.A1(\rbzero.wall_tracer.trackDistY[-1] ),
    .A2(_06216_),
    .B1(_06217_),
    .C1(_06221_),
    .D1(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__o2bb2a_1 _13085_ (.A1_N(_06218_),
    .A2_N(_06240_),
    .B1(\rbzero.wall_tracer.trackDistX[1] ),
    .B2(_06214_),
    .X(_06241_));
 sky130_fd_sc_hd__a221o_1 _13086_ (.A1(_06213_),
    .A2(\rbzero.wall_tracer.trackDistX[2] ),
    .B1(\rbzero.wall_tracer.trackDistX[1] ),
    .B2(_06214_),
    .C1(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__o221a_1 _13087_ (.A1(_06212_),
    .A2(\rbzero.wall_tracer.trackDistX[3] ),
    .B1(_06213_),
    .B2(\rbzero.wall_tracer.trackDistX[2] ),
    .C1(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__a221o_1 _13088_ (.A1(_06211_),
    .A2(\rbzero.wall_tracer.trackDistX[4] ),
    .B1(_06212_),
    .B2(\rbzero.wall_tracer.trackDistX[3] ),
    .C1(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__o221a_1 _13089_ (.A1(\rbzero.wall_tracer.trackDistX[5] ),
    .A2(_06210_),
    .B1(_06211_),
    .B2(\rbzero.wall_tracer.trackDistX[4] ),
    .C1(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__a221o_1 _13090_ (.A1(_06209_),
    .A2(\rbzero.wall_tracer.trackDistX[6] ),
    .B1(\rbzero.wall_tracer.trackDistX[5] ),
    .B2(_06210_),
    .C1(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__o221a_1 _13091_ (.A1(_06208_),
    .A2(\rbzero.wall_tracer.trackDistX[7] ),
    .B1(_06209_),
    .B2(\rbzero.wall_tracer.trackDistX[6] ),
    .C1(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__a221o_1 _13092_ (.A1(_06207_),
    .A2(\rbzero.wall_tracer.trackDistX[8] ),
    .B1(_06208_),
    .B2(\rbzero.wall_tracer.trackDistX[7] ),
    .C1(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__o221a_1 _13093_ (.A1(_06205_),
    .A2(\rbzero.wall_tracer.trackDistX[9] ),
    .B1(_06207_),
    .B2(\rbzero.wall_tracer.trackDistX[8] ),
    .C1(_06248_),
    .X(_06249_));
 sky130_fd_sc_hd__o2bb2a_1 _13094_ (.A1_N(_06206_),
    .A2_N(_06249_),
    .B1(_06204_),
    .B2(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_06250_));
 sky130_fd_sc_hd__a22o_2 _13095_ (.A1(_06204_),
    .A2(\rbzero.wall_tracer.trackDistY[10] ),
    .B1(_06206_),
    .B2(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__nand2_2 _13096_ (.A(_06203_),
    .B(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__or3_1 _13097_ (.A(_06101_),
    .B(_06155_),
    .C(_06201_),
    .X(_06253_));
 sky130_fd_sc_hd__and3_1 _13098_ (.A(_04468_),
    .B(_06252_),
    .C(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__o21ai_4 _13099_ (.A1(_06156_),
    .A2(_06163_),
    .B1(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__nor2_2 _13100_ (.A(_06102_),
    .B(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__a32o_1 _13101_ (.A1(_06098_),
    .A2(_06099_),
    .A3(_06256_),
    .B1(_06255_),
    .B2(\rbzero.wall_tracer.mapY[6] ),
    .X(_00386_));
 sky130_fd_sc_hd__xnor2_1 _13102_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .B(_06076_),
    .Y(_06257_));
 sky130_fd_sc_hd__a21bo_1 _13103_ (.A1(\rbzero.wall_tracer.mapY[6] ),
    .A2(_06081_),
    .B1_N(_06098_),
    .X(_06258_));
 sky130_fd_sc_hd__o21ai_1 _13104_ (.A1(_06257_),
    .A2(_06258_),
    .B1(_06256_),
    .Y(_06259_));
 sky130_fd_sc_hd__a21o_1 _13105_ (.A1(_06257_),
    .A2(_06258_),
    .B1(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__a21bo_1 _13106_ (.A1(\rbzero.wall_tracer.mapY[7] ),
    .A2(_06255_),
    .B1_N(_06260_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _13107_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06081_),
    .X(_06261_));
 sky130_fd_sc_hd__nor2_1 _13108_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06081_),
    .Y(_06262_));
 sky130_fd_sc_hd__nor2_1 _13109_ (.A(_06261_),
    .B(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__o41a_1 _13110_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(\rbzero.wall_tracer.mapY[5] ),
    .A3(\rbzero.wall_tracer.mapY[7] ),
    .A4(\rbzero.wall_tracer.mapY[6] ),
    .B1(_06081_),
    .X(_06264_));
 sky130_fd_sc_hd__a31o_1 _13111_ (.A1(_06097_),
    .A2(_06096_),
    .A3(_06257_),
    .B1(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__xor2_1 _13112_ (.A(_06263_),
    .B(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__a22o_1 _13113_ (.A1(\rbzero.wall_tracer.mapY[8] ),
    .A2(_06255_),
    .B1(_06256_),
    .B2(_06266_),
    .X(_00388_));
 sky130_fd_sc_hd__a21o_1 _13114_ (.A1(_06263_),
    .A2(_06265_),
    .B1(_06261_),
    .X(_06267_));
 sky130_fd_sc_hd__xnor2_1 _13115_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(_06076_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_1 _13116_ (.A(_06267_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__or2_1 _13117_ (.A(_06267_),
    .B(_06268_),
    .X(_06270_));
 sky130_fd_sc_hd__a32o_1 _13118_ (.A1(_06256_),
    .A2(_06269_),
    .A3(_06270_),
    .B1(_06255_),
    .B2(\rbzero.wall_tracer.mapY[9] ),
    .X(_00389_));
 sky130_fd_sc_hd__o21a_1 _13119_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06081_),
    .B1(_06267_),
    .X(_06271_));
 sky130_fd_sc_hd__a21o_1 _13120_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06081_),
    .B1(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__xor2_1 _13121_ (.A(\rbzero.wall_tracer.mapY[10] ),
    .B(_06076_),
    .X(_06273_));
 sky130_fd_sc_hd__xnor2_1 _13122_ (.A(_06272_),
    .B(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__a22o_1 _13123_ (.A1(\rbzero.wall_tracer.mapY[10] ),
    .A2(_06255_),
    .B1(_06256_),
    .B2(_06274_),
    .X(_00390_));
 sky130_fd_sc_hd__inv_2 _13124_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06275_));
 sky130_fd_sc_hd__buf_4 _13125_ (.A(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__a31o_1 _13126_ (.A1(_05995_),
    .A2(_05997_),
    .A3(_06028_),
    .B1(_06030_),
    .X(_06277_));
 sky130_fd_sc_hd__inv_2 _13127_ (.A(_04463_),
    .Y(_06278_));
 sky130_fd_sc_hd__buf_2 _13128_ (.A(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__a311o_4 _13129_ (.A1(_06032_),
    .A2(_06029_),
    .A3(_06277_),
    .B1(_06072_),
    .C1(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__and2_1 _13130_ (.A(_06276_),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__or2_1 _13131_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_04464_),
    .X(_06282_));
 sky130_fd_sc_hd__and2_1 _13132_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .X(_06283_));
 sky130_fd_sc_hd__nand2_1 _13133_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_06284_));
 sky130_fd_sc_hd__or2_1 _13134_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_06285_));
 sky130_fd_sc_hd__nand3_1 _13135_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .C(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__xor2_2 _13136_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06287_));
 sky130_fd_sc_hd__nand2_1 _13137_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_06288_));
 sky130_fd_sc_hd__or2_1 _13138_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06289_));
 sky130_fd_sc_hd__nand3_1 _13139_ (.A(_06287_),
    .B(_06288_),
    .C(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__and2_1 _13140_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_06291_));
 sky130_fd_sc_hd__a21o_1 _13141_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[4] ),
    .B1(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__o21ai_1 _13142_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[4] ),
    .B1(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__nor2_1 _13143_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06294_));
 sky130_fd_sc_hd__nor2_1 _13144_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06295_));
 sky130_fd_sc_hd__nand2_2 _13145_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_06296_));
 sky130_fd_sc_hd__nor2_1 _13146_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06297_));
 sky130_fd_sc_hd__nand2_1 _13147_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06298_));
 sky130_fd_sc_hd__nand2_1 _13148_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06299_));
 sky130_fd_sc_hd__o211a_1 _13149_ (.A1(_06296_),
    .A2(_06297_),
    .B1(_06298_),
    .C1(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__nand2_1 _13150_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06301_));
 sky130_fd_sc_hd__o31ai_4 _13151_ (.A1(_06294_),
    .A2(_06295_),
    .A3(_06300_),
    .B1(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__xor2_2 _13152_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_06303_));
 sky130_fd_sc_hd__xor2_2 _13153_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_06304_));
 sky130_fd_sc_hd__and2_1 _13154_ (.A(_06303_),
    .B(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__and2b_1 _13155_ (.A_N(_06290_),
    .B(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__a2bb2o_1 _13156_ (.A1_N(_06290_),
    .A2_N(_06293_),
    .B1(_06302_),
    .B2(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__and2_1 _13157_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06308_));
 sky130_fd_sc_hd__a21bo_1 _13158_ (.A1(_06308_),
    .A2(_06289_),
    .B1_N(_06288_),
    .X(_06309_));
 sky130_fd_sc_hd__nand2_1 _13159_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_06310_));
 sky130_fd_sc_hd__or2_1 _13160_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_06311_));
 sky130_fd_sc_hd__nand2_1 _13161_ (.A(_06310_),
    .B(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__inv_2 _13162_ (.A(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__o2111ai_1 _13163_ (.A1(_06307_),
    .A2(_06309_),
    .B1(_06313_),
    .C1(_06284_),
    .D1(_06285_),
    .Y(_06314_));
 sky130_fd_sc_hd__nand2_1 _13164_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_06315_));
 sky130_fd_sc_hd__nor2_1 _13165_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_06316_));
 sky130_fd_sc_hd__a41o_2 _13166_ (.A1(_06284_),
    .A2(_06286_),
    .A3(_06314_),
    .A4(_06315_),
    .B1(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__or2_1 _13167_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .X(_06318_));
 sky130_fd_sc_hd__o211a_4 _13168_ (.A1(_06283_),
    .A2(_06317_),
    .B1(_04479_),
    .C1(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__a21oi_2 _13169_ (.A1(_06281_),
    .A2(_06282_),
    .B1(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__or2_1 _13170_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_04464_),
    .X(_06321_));
 sky130_fd_sc_hd__a31o_1 _13171_ (.A1(_06276_),
    .A2(_06280_),
    .A3(_06321_),
    .B1(_06319_),
    .X(_06322_));
 sky130_fd_sc_hd__a21o_1 _13172_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_06279_),
    .B1(_04480_),
    .X(_06323_));
 sky130_fd_sc_hd__a21o_1 _13173_ (.A1(_04464_),
    .A2(_06035_),
    .B1(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__nand2_1 _13174_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_06325_));
 sky130_fd_sc_hd__nand2_1 _13175_ (.A(_06318_),
    .B(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__xnor2_2 _13176_ (.A(_06317_),
    .B(_06326_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand2_1 _13177_ (.A(_04480_),
    .B(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__and3_1 _13178_ (.A(_06284_),
    .B(_06286_),
    .C(_06314_),
    .X(_06329_));
 sky130_fd_sc_hd__and2b_1 _13179_ (.A_N(_06316_),
    .B(_06315_),
    .X(_06330_));
 sky130_fd_sc_hd__xnor2_2 _13180_ (.A(_06329_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__or3_1 _13181_ (.A(_06279_),
    .B(_06037_),
    .C(_06038_),
    .X(_06332_));
 sky130_fd_sc_hd__o21a_1 _13182_ (.A1(\rbzero.wall_tracer.visualWallDist[1] ),
    .A2(_04463_),
    .B1(_06276_),
    .X(_06333_));
 sky130_fd_sc_hd__a22o_1 _13183_ (.A1(_04480_),
    .A2(_06331_),
    .B1(_06332_),
    .B2(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__a21o_1 _13184_ (.A1(_06324_),
    .A2(_06328_),
    .B1(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__or2_1 _13185_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_04464_),
    .X(_06336_));
 sky130_fd_sc_hd__a31oi_4 _13186_ (.A1(_06276_),
    .A2(_06280_),
    .A3(_06336_),
    .B1(_06319_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _13187_ (.A(_06288_),
    .B(_06289_),
    .Y(_06338_));
 sky130_fd_sc_hd__a21bo_1 _13188_ (.A1(_06302_),
    .A2(_06305_),
    .B1_N(_06293_),
    .X(_06339_));
 sky130_fd_sc_hd__a21oi_1 _13189_ (.A1(_06287_),
    .A2(_06339_),
    .B1(_06308_),
    .Y(_06340_));
 sky130_fd_sc_hd__xnor2_2 _13190_ (.A(_06338_),
    .B(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__and2_1 _13191_ (.A(_04479_),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__a21oi_1 _13192_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_06279_),
    .B1(_04479_),
    .Y(_06343_));
 sky130_fd_sc_hd__o31a_1 _13193_ (.A1(_06279_),
    .A2(_06042_),
    .A3(_06043_),
    .B1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__xnor2_2 _13194_ (.A(_06287_),
    .B(_06339_),
    .Y(_06345_));
 sky130_fd_sc_hd__a21o_1 _13195_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_06278_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06346_));
 sky130_fd_sc_hd__a31o_1 _13196_ (.A1(_04463_),
    .A2(_06041_),
    .A3(_06047_),
    .B1(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__a21bo_2 _13197_ (.A1(_04479_),
    .A2(_06345_),
    .B1_N(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__a21o_1 _13198_ (.A1(_06302_),
    .A2(_06303_),
    .B1(_06291_),
    .X(_06349_));
 sky130_fd_sc_hd__xnor2_2 _13199_ (.A(_06304_),
    .B(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__nand2_1 _13200_ (.A(_04463_),
    .B(_06052_),
    .Y(_06351_));
 sky130_fd_sc_hd__a21oi_1 _13201_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_06279_),
    .B1(_04479_),
    .Y(_06352_));
 sky130_fd_sc_hd__a22o_4 _13202_ (.A1(_04479_),
    .A2(_06350_),
    .B1(_06351_),
    .B2(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__xnor2_2 _13203_ (.A(_06302_),
    .B(_06303_),
    .Y(_06354_));
 sky130_fd_sc_hd__a21o_1 _13204_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_06279_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06355_));
 sky130_fd_sc_hd__and3_1 _13205_ (.A(_04463_),
    .B(_06040_),
    .C(_06053_),
    .X(_06356_));
 sky130_fd_sc_hd__o2bb2a_2 _13206_ (.A1_N(_04479_),
    .A2_N(_06354_),
    .B1(_06355_),
    .B2(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__or2_1 _13207_ (.A(_06294_),
    .B(_06300_),
    .X(_06358_));
 sky130_fd_sc_hd__and2b_1 _13208_ (.A_N(_06295_),
    .B(_06301_),
    .X(_06359_));
 sky130_fd_sc_hd__xnor2_2 _13209_ (.A(_06358_),
    .B(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__or2_1 _13210_ (.A(_06278_),
    .B(_06058_),
    .X(_06361_));
 sky130_fd_sc_hd__o21a_1 _13211_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_04463_),
    .B1(_06276_),
    .X(_06362_));
 sky130_fd_sc_hd__o21ai_1 _13212_ (.A1(_06296_),
    .A2(_06297_),
    .B1(_06298_),
    .Y(_06363_));
 sky130_fd_sc_hd__and2_1 _13213_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_06364_));
 sky130_fd_sc_hd__nor2_1 _13214_ (.A(_06364_),
    .B(_06294_),
    .Y(_06365_));
 sky130_fd_sc_hd__xnor2_1 _13215_ (.A(_06363_),
    .B(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__nand2_1 _13216_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__a21o_1 _13217_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_06278_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06368_));
 sky130_fd_sc_hd__a21o_1 _13218_ (.A1(_04463_),
    .A2(_06060_),
    .B1(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06370_));
 sky130_fd_sc_hd__mux2_2 _13220_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_06370_),
    .S(_06275_),
    .X(_06371_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06372_));
 sky130_fd_sc_hd__mux2_2 _13222_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_06372_),
    .S(_06275_),
    .X(_06373_));
 sky130_fd_sc_hd__or2_1 _13223_ (.A(_06371_),
    .B(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__or2_1 _13224_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_06375_));
 sky130_fd_sc_hd__and2_1 _13225_ (.A(_06296_),
    .B(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__mux2_1 _13226_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_06063_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06377_));
 sky130_fd_sc_hd__mux2_2 _13227_ (.A0(_06376_),
    .A1(_06377_),
    .S(_06275_),
    .X(_06378_));
 sky130_fd_sc_hd__or2_1 _13228_ (.A(_06374_),
    .B(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__or2b_1 _13229_ (.A(_06297_),
    .B_N(_06298_),
    .X(_06380_));
 sky130_fd_sc_hd__xor2_2 _13230_ (.A(_06296_),
    .B(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__mux2_1 _13231_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_06062_),
    .S(_04463_),
    .X(_06382_));
 sky130_fd_sc_hd__mux2_4 _13232_ (.A0(_06381_),
    .A1(_06382_),
    .S(_06276_),
    .X(_06383_));
 sky130_fd_sc_hd__a211o_1 _13233_ (.A1(_06367_),
    .A2(_06369_),
    .B1(_06379_),
    .C1(_06383_),
    .X(_06384_));
 sky130_fd_sc_hd__a221o_1 _13234_ (.A1(\rbzero.wall_tracer.rcp_sel[0] ),
    .A2(_06360_),
    .B1(_06361_),
    .B2(_06362_),
    .C1(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__nor2_2 _13235_ (.A(_06357_),
    .B(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__o2111a_1 _13236_ (.A1(_06342_),
    .A2(_06344_),
    .B1(_06348_),
    .C1(_06353_),
    .D1(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__o21ai_1 _13237_ (.A1(_06307_),
    .A2(_06309_),
    .B1(_06313_),
    .Y(_06388_));
 sky130_fd_sc_hd__nand2_1 _13238_ (.A(_06285_),
    .B(_06284_),
    .Y(_06389_));
 sky130_fd_sc_hd__a21oi_1 _13239_ (.A1(_06310_),
    .A2(_06388_),
    .B1(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__and3_1 _13240_ (.A(_06310_),
    .B(_06388_),
    .C(_06389_),
    .X(_06391_));
 sky130_fd_sc_hd__o21ai_1 _13241_ (.A1(_06390_),
    .A2(_06391_),
    .B1(_04480_),
    .Y(_06392_));
 sky130_fd_sc_hd__a21o_1 _13242_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_06279_),
    .B1(_04479_),
    .X(_06393_));
 sky130_fd_sc_hd__a31o_1 _13243_ (.A1(_04464_),
    .A2(_06068_),
    .A3(_06069_),
    .B1(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__or3_1 _13244_ (.A(_06307_),
    .B(_06309_),
    .C(_06313_),
    .X(_06395_));
 sky130_fd_sc_hd__nand2_2 _13245_ (.A(_06388_),
    .B(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__a21oi_1 _13246_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_06279_),
    .B1(_04479_),
    .Y(_06397_));
 sky130_fd_sc_hd__o31a_1 _13247_ (.A1(_06279_),
    .A2(_06049_),
    .A3(_06050_),
    .B1(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__a21oi_1 _13248_ (.A1(_04480_),
    .A2(_06396_),
    .B1(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__a21oi_1 _13249_ (.A1(_06392_),
    .A2(_06394_),
    .B1(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__nand3_1 _13250_ (.A(_06337_),
    .B(_06387_),
    .C(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__or2_1 _13251_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_04464_),
    .X(_06402_));
 sky130_fd_sc_hd__a31o_1 _13252_ (.A1(_06276_),
    .A2(_06280_),
    .A3(_06402_),
    .B1(_06319_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_4 _13253_ (.A(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__o31a_1 _13254_ (.A1(_06322_),
    .A2(_06335_),
    .A3(_06401_),
    .B1(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__xnor2_2 _13255_ (.A(_06320_),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__o21ai_1 _13256_ (.A1(_06335_),
    .A2(_06401_),
    .B1(_06404_),
    .Y(_06407_));
 sky130_fd_sc_hd__xnor2_2 _13257_ (.A(_06322_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__or2_2 _13258_ (.A(_06406_),
    .B(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__or2_1 _13259_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_04464_),
    .X(_06410_));
 sky130_fd_sc_hd__a21oi_1 _13260_ (.A1(_06280_),
    .A2(_06410_),
    .B1(_04480_),
    .Y(_06411_));
 sky130_fd_sc_hd__clkinv_2 _13261_ (.A(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__o21ai_2 _13262_ (.A1(_06283_),
    .A2(_06317_),
    .B1(_06318_),
    .Y(_06413_));
 sky130_fd_sc_hd__a21o_1 _13263_ (.A1(_04480_),
    .A2(_06413_),
    .B1(_06411_),
    .X(_06414_));
 sky130_fd_sc_hd__nor3_1 _13264_ (.A(_06322_),
    .B(_06335_),
    .C(_06401_),
    .Y(_06415_));
 sky130_fd_sc_hd__o21a_1 _13265_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_04464_),
    .B1(_06281_),
    .X(_06416_));
 sky130_fd_sc_hd__or2_1 _13266_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_04463_),
    .X(_06417_));
 sky130_fd_sc_hd__a31oi_4 _13267_ (.A1(_06276_),
    .A2(_06280_),
    .A3(_06417_),
    .B1(_06319_),
    .Y(_06418_));
 sky130_fd_sc_hd__a21bo_1 _13268_ (.A1(_06281_),
    .A2(_06282_),
    .B1_N(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__or2_1 _13269_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_04464_),
    .X(_06420_));
 sky130_fd_sc_hd__a31o_1 _13270_ (.A1(_06276_),
    .A2(_06280_),
    .A3(_06420_),
    .B1(_06319_),
    .X(_06421_));
 sky130_fd_sc_hd__nor3_1 _13271_ (.A(_06416_),
    .B(_06419_),
    .C(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__a31oi_1 _13272_ (.A1(_06276_),
    .A2(_06280_),
    .A3(_06402_),
    .B1(_06319_),
    .Y(_06423_));
 sky130_fd_sc_hd__clkbuf_4 _13273_ (.A(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__a21o_1 _13274_ (.A1(_06415_),
    .A2(_06422_),
    .B1(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__mux2_2 _13275_ (.A0(_06412_),
    .A1(_06414_),
    .S(_06425_),
    .X(_06426_));
 sky130_fd_sc_hd__nand2_1 _13276_ (.A(_06281_),
    .B(_06402_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand2_1 _13277_ (.A(_06415_),
    .B(_06422_),
    .Y(_06428_));
 sky130_fd_sc_hd__or3_2 _13278_ (.A(_06427_),
    .B(_06428_),
    .C(_06410_),
    .X(_06429_));
 sky130_fd_sc_hd__or4_1 _13279_ (.A(_06322_),
    .B(_06335_),
    .C(_06401_),
    .D(_06419_),
    .X(_06430_));
 sky130_fd_sc_hd__or2_1 _13280_ (.A(_06319_),
    .B(_06416_),
    .X(_06431_));
 sky130_fd_sc_hd__o211a_1 _13281_ (.A1(_06421_),
    .A2(_06430_),
    .B1(_06431_),
    .C1(_06404_),
    .X(_06432_));
 sky130_fd_sc_hd__a21oi_1 _13282_ (.A1(_06281_),
    .A2(_06420_),
    .B1(_06319_),
    .Y(_06433_));
 sky130_fd_sc_hd__nor2_1 _13283_ (.A(_06424_),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__a211oi_1 _13284_ (.A1(_06404_),
    .A2(_06430_),
    .B1(_06431_),
    .C1(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__or3b_1 _13285_ (.A(_06424_),
    .B(_06421_),
    .C_N(_06430_),
    .X(_06436_));
 sky130_fd_sc_hd__a21o_1 _13286_ (.A1(_06404_),
    .A2(_06430_),
    .B1(_06433_),
    .X(_06437_));
 sky130_fd_sc_hd__o211a_1 _13287_ (.A1(_06432_),
    .A2(_06435_),
    .B1(_06436_),
    .C1(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__a21oi_2 _13288_ (.A1(_06415_),
    .A2(_06320_),
    .B1(_06424_),
    .Y(_06439_));
 sky130_fd_sc_hd__xor2_2 _13289_ (.A(_06418_),
    .B(_06439_),
    .X(_06440_));
 sky130_fd_sc_hd__nand4_4 _13290_ (.A(_06426_),
    .B(_06429_),
    .C(_06438_),
    .D(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__a21o_1 _13291_ (.A1(_06387_),
    .A2(_06400_),
    .B1(_06423_),
    .X(_06442_));
 sky130_fd_sc_hd__a21bo_1 _13292_ (.A1(_06403_),
    .A2(_06335_),
    .B1_N(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__xnor2_2 _13293_ (.A(_06337_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__xnor2_2 _13294_ (.A(_06334_),
    .B(_06442_),
    .Y(_06445_));
 sky130_fd_sc_hd__and2_1 _13295_ (.A(_06392_),
    .B(_06394_),
    .X(_06446_));
 sky130_fd_sc_hd__a21o_1 _13296_ (.A1(_04480_),
    .A2(_06396_),
    .B1(_06398_),
    .X(_06447_));
 sky130_fd_sc_hd__a21o_1 _13297_ (.A1(_06447_),
    .A2(_06387_),
    .B1(_06424_),
    .X(_06448_));
 sky130_fd_sc_hd__xnor2_2 _13298_ (.A(_06446_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__nand2_1 _13299_ (.A(_06324_),
    .B(_06328_),
    .Y(_06450_));
 sky130_fd_sc_hd__o2111ai_1 _13300_ (.A1(_06342_),
    .A2(_06344_),
    .B1(_06348_),
    .C1(_06353_),
    .D1(_06386_),
    .Y(_06451_));
 sky130_fd_sc_hd__a21o_1 _13301_ (.A1(_06392_),
    .A2(_06394_),
    .B1(_06399_),
    .X(_06452_));
 sky130_fd_sc_hd__o31a_1 _13302_ (.A1(_06334_),
    .A2(_06451_),
    .A3(_06452_),
    .B1(_06403_),
    .X(_06453_));
 sky130_fd_sc_hd__xnor2_2 _13303_ (.A(_06450_),
    .B(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__or3_1 _13304_ (.A(_06445_),
    .B(_06449_),
    .C(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__or2_1 _13305_ (.A(_06444_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__nor2_1 _13306_ (.A(_06424_),
    .B(_06387_),
    .Y(_06457_));
 sky130_fd_sc_hd__xnor2_2 _13307_ (.A(_06447_),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__nor2_1 _13308_ (.A(_06456_),
    .B(_06458_),
    .Y(_06459_));
 sky130_fd_sc_hd__or3b_4 _13309_ (.A(_06409_),
    .B(_06441_),
    .C_N(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_4 _13310_ (.A(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__nor2_2 _13311_ (.A(_06342_),
    .B(_06344_),
    .Y(_06462_));
 sky130_fd_sc_hd__a31oi_4 _13312_ (.A1(_06348_),
    .A2(_06353_),
    .A3(_06386_),
    .B1(_06424_),
    .Y(_06463_));
 sky130_fd_sc_hd__xor2_4 _13313_ (.A(_06462_),
    .B(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__nor2_1 _13314_ (.A(_06406_),
    .B(_06408_),
    .Y(_06465_));
 sky130_fd_sc_hd__and4_1 _13315_ (.A(_06426_),
    .B(_06429_),
    .C(_06438_),
    .D(_06440_),
    .X(_06466_));
 sky130_fd_sc_hd__and3_2 _13316_ (.A(_06465_),
    .B(_06466_),
    .C(_06459_),
    .X(_06467_));
 sky130_fd_sc_hd__nand2_2 _13317_ (.A(_06367_),
    .B(_06369_),
    .Y(_06468_));
 sky130_fd_sc_hd__nor2_1 _13318_ (.A(_06379_),
    .B(_06383_),
    .Y(_06469_));
 sky130_fd_sc_hd__or2_2 _13319_ (.A(_06469_),
    .B(_06424_),
    .X(_06470_));
 sky130_fd_sc_hd__xor2_4 _13320_ (.A(_06468_),
    .B(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__a21o_1 _13321_ (.A1(_06353_),
    .A2(_06386_),
    .B1(_06424_),
    .X(_06472_));
 sky130_fd_sc_hd__xor2_4 _13322_ (.A(_06348_),
    .B(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__nand2_2 _13323_ (.A(_06404_),
    .B(_06385_),
    .Y(_06474_));
 sky130_fd_sc_hd__xnor2_4 _13324_ (.A(_06357_),
    .B(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__nor2_2 _13325_ (.A(_06424_),
    .B(_06386_),
    .Y(_06476_));
 sky130_fd_sc_hd__xnor2_4 _13326_ (.A(_06353_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__a22o_2 _13327_ (.A1(_04480_),
    .A2(_06360_),
    .B1(_06361_),
    .B2(_06362_),
    .X(_06478_));
 sky130_fd_sc_hd__nand2_2 _13328_ (.A(_06404_),
    .B(_06384_),
    .Y(_06479_));
 sky130_fd_sc_hd__xnor2_2 _13329_ (.A(_06478_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__or3_1 _13330_ (.A(_06475_),
    .B(_06477_),
    .C(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__nor3_1 _13331_ (.A(_06471_),
    .B(_06473_),
    .C(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__and4b_1 _13332_ (.A_N(_06464_),
    .B(_06467_),
    .C(_06482_),
    .D(_06469_),
    .X(_06483_));
 sky130_fd_sc_hd__clkbuf_4 _13333_ (.A(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__or4b_2 _13334_ (.A(_06409_),
    .B(_06441_),
    .C(_06464_),
    .D_N(_06459_),
    .X(_06485_));
 sky130_fd_sc_hd__and2_2 _13335_ (.A(_06379_),
    .B(_06404_),
    .X(_06486_));
 sky130_fd_sc_hd__xor2_4 _13336_ (.A(_06383_),
    .B(_06486_),
    .X(_06487_));
 sky130_fd_sc_hd__nand2_1 _13337_ (.A(_06374_),
    .B(_06404_),
    .Y(_06488_));
 sky130_fd_sc_hd__xnor2_4 _13338_ (.A(_06378_),
    .B(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__nor2_1 _13339_ (.A(_06487_),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_06371_),
    .B(_06404_),
    .Y(_06491_));
 sky130_fd_sc_hd__xor2_2 _13341_ (.A(_06373_),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__and3_1 _13342_ (.A(_06371_),
    .B(_06490_),
    .C(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__and3b_1 _13343_ (.A_N(_06485_),
    .B(_06482_),
    .C(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__and2b_1 _13344_ (.A_N(_06464_),
    .B(_06473_),
    .X(_06495_));
 sky130_fd_sc_hd__and4_1 _13345_ (.A(_06465_),
    .B(_06466_),
    .C(_06459_),
    .D(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__or4b_1 _13346_ (.A(_06445_),
    .B(_06449_),
    .C(_06458_),
    .D_N(_06464_),
    .X(_06497_));
 sky130_fd_sc_hd__or2_1 _13347_ (.A(_06454_),
    .B(_06444_),
    .X(_06498_));
 sky130_fd_sc_hd__nor2_1 _13348_ (.A(_06409_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__nor3b_1 _13349_ (.A(_06441_),
    .B(_06497_),
    .C_N(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__or2_1 _13350_ (.A(_06458_),
    .B(_06464_),
    .X(_06501_));
 sky130_fd_sc_hd__or3_1 _13351_ (.A(_06473_),
    .B(_06456_),
    .C(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__xor2_1 _13352_ (.A(_06357_),
    .B(_06474_),
    .X(_06503_));
 sky130_fd_sc_hd__nor2_1 _13353_ (.A(_06503_),
    .B(_06477_),
    .Y(_06504_));
 sky130_fd_sc_hd__or4b_1 _13354_ (.A(_06409_),
    .B(_06441_),
    .C(_06502_),
    .D_N(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__or3b_4 _13355_ (.A(_06496_),
    .B(_06500_),
    .C_N(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__nand2_1 _13356_ (.A(_06426_),
    .B(_06429_),
    .Y(_06507_));
 sky130_fd_sc_hd__or2b_1 _13357_ (.A(_06507_),
    .B_N(_06438_),
    .X(_06508_));
 sky130_fd_sc_hd__nor4b_1 _13358_ (.A(_06473_),
    .B(_06456_),
    .C(_06501_),
    .D_N(_06477_),
    .Y(_06509_));
 sky130_fd_sc_hd__nor2_1 _13359_ (.A(_06501_),
    .B(_06492_),
    .Y(_06510_));
 sky130_fd_sc_hd__and4b_1 _13360_ (.A_N(_06456_),
    .B(_06482_),
    .C(_06490_),
    .D(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__and4bb_1 _13361_ (.A_N(_06509_),
    .B_N(_06511_),
    .C(_06440_),
    .D(_06465_),
    .X(_06512_));
 sky130_fd_sc_hd__or3b_1 _13362_ (.A(_06409_),
    .B(_06441_),
    .C_N(_06444_),
    .X(_06513_));
 sky130_fd_sc_hd__o21ai_2 _13363_ (.A1(_06508_),
    .A2(_06512_),
    .B1(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__or4_1 _13364_ (.A(_06484_),
    .B(_06494_),
    .C(_06506_),
    .D(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__clkbuf_8 _13365_ (.A(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__or2_1 _13366_ (.A(_06455_),
    .B(_06458_),
    .X(_06517_));
 sky130_fd_sc_hd__nor2_1 _13367_ (.A(_06409_),
    .B(_06444_),
    .Y(_06518_));
 sky130_fd_sc_hd__and2_1 _13368_ (.A(_06466_),
    .B(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__and3_1 _13369_ (.A(_06465_),
    .B(_06466_),
    .C(_06509_),
    .X(_06520_));
 sky130_fd_sc_hd__a21o_1 _13370_ (.A1(_06517_),
    .A2(_06519_),
    .B1(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__or2_2 _13371_ (.A(_06506_),
    .B(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__xnor2_4 _13372_ (.A(_06516_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__or3_1 _13373_ (.A(_06471_),
    .B(_06473_),
    .C(_06481_),
    .X(_06524_));
 sky130_fd_sc_hd__inv_2 _13374_ (.A(_06489_),
    .Y(_06525_));
 sky130_fd_sc_hd__o41a_4 _13375_ (.A1(_06485_),
    .A2(_06524_),
    .A3(_06487_),
    .A4(_06525_),
    .B1(_06505_),
    .X(_06526_));
 sky130_fd_sc_hd__and4bb_2 _13376_ (.A_N(_06441_),
    .B_N(_06455_),
    .C(_06458_),
    .D(_06518_),
    .X(_06527_));
 sky130_fd_sc_hd__a311o_1 _13377_ (.A1(_06466_),
    .A2(_06445_),
    .A3(_06499_),
    .B1(_06527_),
    .C1(_06496_),
    .X(_06528_));
 sky130_fd_sc_hd__xnor2_1 _13378_ (.A(_06468_),
    .B(_06470_),
    .Y(_06529_));
 sky130_fd_sc_hd__or4_1 _13379_ (.A(_06529_),
    .B(_06473_),
    .C(_06485_),
    .D(_06481_),
    .X(_06530_));
 sky130_fd_sc_hd__inv_2 _13380_ (.A(_06406_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_1 _13381_ (.A(_06436_),
    .B(_06437_),
    .Y(_06532_));
 sky130_fd_sc_hd__or2_1 _13382_ (.A(_06432_),
    .B(_06435_),
    .X(_06533_));
 sky130_fd_sc_hd__nand2_1 _13383_ (.A(_06532_),
    .B(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__o2111a_1 _13384_ (.A1(_06531_),
    .A2(_06441_),
    .B1(_06513_),
    .C1(_06534_),
    .D1(_06426_),
    .X(_06535_));
 sky130_fd_sc_hd__and4bb_4 _13385_ (.A_N(_06494_),
    .B_N(_06528_),
    .C(_06530_),
    .D(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__nor2_1 _13386_ (.A(_06520_),
    .B(_06527_),
    .Y(_06537_));
 sky130_fd_sc_hd__nor3b_1 _13387_ (.A(_06498_),
    .B(_06445_),
    .C_N(_06449_),
    .Y(_06538_));
 sky130_fd_sc_hd__and4bb_1 _13388_ (.A_N(_06456_),
    .B_N(_06501_),
    .C(_06482_),
    .D(_06487_),
    .X(_06539_));
 sky130_fd_sc_hd__o311ai_1 _13389_ (.A1(_06408_),
    .A2(_06538_),
    .A3(_06539_),
    .B1(_06466_),
    .C1(_06531_),
    .Y(_06540_));
 sky130_fd_sc_hd__o211a_1 _13390_ (.A1(_06507_),
    .A2(_06438_),
    .B1(_06513_),
    .C1(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__and4b_1 _13391_ (.A_N(_06484_),
    .B(_06537_),
    .C(_06526_),
    .D(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__a211o_2 _13392_ (.A1(_06526_),
    .A2(_06536_),
    .B1(_06542_),
    .C1(_06516_),
    .X(_06543_));
 sky130_fd_sc_hd__a21oi_4 _13393_ (.A1(_06523_),
    .A2(_06543_),
    .B1(_06527_),
    .Y(_06544_));
 sky130_fd_sc_hd__buf_4 _13394_ (.A(_06484_),
    .X(_06545_));
 sky130_fd_sc_hd__buf_4 _13395_ (.A(_06542_),
    .X(_06546_));
 sky130_fd_sc_hd__a21oi_4 _13396_ (.A1(_06526_),
    .A2(_06536_),
    .B1(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__xnor2_4 _13397_ (.A(_06516_),
    .B(_06547_),
    .Y(_06548_));
 sky130_fd_sc_hd__buf_2 _13398_ (.A(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__nor2_1 _13399_ (.A(_06545_),
    .B(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__nand2_2 _13400_ (.A(_06526_),
    .B(_06536_),
    .Y(_06551_));
 sky130_fd_sc_hd__buf_2 _13401_ (.A(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__clkbuf_4 _13402_ (.A(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__buf_2 _13403_ (.A(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__clkbuf_4 _13404_ (.A(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__or2_4 _13405_ (.A(_06460_),
    .B(_06544_),
    .X(_06556_));
 sky130_fd_sc_hd__nor2_2 _13406_ (.A(_06485_),
    .B(_06524_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_4 _13407_ (.A(_06469_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__nand4_4 _13408_ (.A(_06558_),
    .B(_06537_),
    .C(_06526_),
    .D(_06541_),
    .Y(_06559_));
 sky130_fd_sc_hd__clkbuf_4 _13409_ (.A(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__and3_1 _13410_ (.A(_06477_),
    .B(_06526_),
    .C(_06536_),
    .X(_06561_));
 sky130_fd_sc_hd__a21o_1 _13411_ (.A1(_06473_),
    .A2(_06560_),
    .B1(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__and3_1 _13412_ (.A(_06480_),
    .B(_06526_),
    .C(_06536_),
    .X(_06563_));
 sky130_fd_sc_hd__a21o_1 _13413_ (.A1(_06475_),
    .A2(_06553_),
    .B1(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__and3_1 _13414_ (.A(_06526_),
    .B(_06546_),
    .C(_06536_),
    .X(_06565_));
 sky130_fd_sc_hd__nor2_4 _13415_ (.A(_06547_),
    .B(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__mux2_1 _13416_ (.A0(_06562_),
    .A1(_06564_),
    .S(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__xnor2_1 _13417_ (.A(_06373_),
    .B(_06491_),
    .Y(_06568_));
 sky130_fd_sc_hd__and2_1 _13418_ (.A(_06526_),
    .B(_06536_),
    .X(_06569_));
 sky130_fd_sc_hd__buf_2 _13419_ (.A(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__mux4_1 _13420_ (.A0(_06471_),
    .A1(_06489_),
    .A2(_06568_),
    .A3(_06487_),
    .S0(_06546_),
    .S1(_06570_),
    .X(_06571_));
 sky130_fd_sc_hd__mux2_1 _13421_ (.A0(_06567_),
    .A1(_06571_),
    .S(_06548_),
    .X(_06572_));
 sky130_fd_sc_hd__nor2_4 _13422_ (.A(_06516_),
    .B(_06546_),
    .Y(_06573_));
 sky130_fd_sc_hd__xnor2_2 _13423_ (.A(_06383_),
    .B(_06486_),
    .Y(_06574_));
 sky130_fd_sc_hd__nand2_4 _13424_ (.A(_06557_),
    .B(_06574_),
    .Y(_06575_));
 sky130_fd_sc_hd__a31o_1 _13425_ (.A1(_06371_),
    .A2(_06554_),
    .A3(_06573_),
    .B1(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__or2_2 _13426_ (.A(_06516_),
    .B(_06521_),
    .X(_06577_));
 sky130_fd_sc_hd__nor3b_4 _13427_ (.A(_06506_),
    .B(_06520_),
    .C_N(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__mux2_1 _13428_ (.A0(_06449_),
    .A1(_06458_),
    .S(_06552_),
    .X(_06579_));
 sky130_fd_sc_hd__mux2_1 _13429_ (.A0(_06473_),
    .A1(_06464_),
    .S(_06570_),
    .X(_06580_));
 sky130_fd_sc_hd__mux2_1 _13430_ (.A0(_06579_),
    .A1(_06580_),
    .S(_06559_),
    .X(_06581_));
 sky130_fd_sc_hd__mux2_1 _13431_ (.A0(_06408_),
    .A1(_06444_),
    .S(_06552_),
    .X(_06582_));
 sky130_fd_sc_hd__mux2_1 _13432_ (.A0(_06445_),
    .A1(_06454_),
    .S(_06570_),
    .X(_06583_));
 sky130_fd_sc_hd__mux2_1 _13433_ (.A0(_06582_),
    .A1(_06583_),
    .S(_06559_),
    .X(_06584_));
 sky130_fd_sc_hd__clkbuf_4 _13434_ (.A(_06516_),
    .X(_06585_));
 sky130_fd_sc_hd__mux2_2 _13435_ (.A0(_06581_),
    .A1(_06584_),
    .S(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__clkbuf_4 _13436_ (.A(_06546_),
    .X(_06587_));
 sky130_fd_sc_hd__xnor2_1 _13437_ (.A(_06418_),
    .B(_06439_),
    .Y(_06588_));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(_06588_),
    .A1(_06406_),
    .S(_06553_),
    .X(_06589_));
 sky130_fd_sc_hd__a21o_1 _13439_ (.A1(_06532_),
    .A2(_06553_),
    .B1(_06560_),
    .X(_06590_));
 sky130_fd_sc_hd__o21a_1 _13440_ (.A1(_06587_),
    .A2(_06589_),
    .B1(_06590_),
    .X(_06591_));
 sky130_fd_sc_hd__a211o_1 _13441_ (.A1(_06578_),
    .A2(_06586_),
    .B1(_06591_),
    .C1(_06467_),
    .X(_06592_));
 sky130_fd_sc_hd__o211a_2 _13442_ (.A1(_06556_),
    .A2(_06572_),
    .B1(_06576_),
    .C1(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__inv_2 _13443_ (.A(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__buf_4 _13444_ (.A(_06578_),
    .X(_06595_));
 sky130_fd_sc_hd__mux2_1 _13445_ (.A0(_06454_),
    .A1(_06444_),
    .S(_06570_),
    .X(_06596_));
 sky130_fd_sc_hd__mux2_1 _13446_ (.A0(_06445_),
    .A1(_06449_),
    .S(_06551_),
    .X(_06597_));
 sky130_fd_sc_hd__mux2_1 _13447_ (.A0(_06596_),
    .A1(_06597_),
    .S(_06559_),
    .X(_06598_));
 sky130_fd_sc_hd__mux2_1 _13448_ (.A0(_06458_),
    .A1(_06464_),
    .S(_06551_),
    .X(_06599_));
 sky130_fd_sc_hd__mux2_1 _13449_ (.A0(_06473_),
    .A1(_06477_),
    .S(_06551_),
    .X(_06600_));
 sky130_fd_sc_hd__mux2_1 _13450_ (.A0(_06599_),
    .A1(_06600_),
    .S(_06559_),
    .X(_06601_));
 sky130_fd_sc_hd__or2_2 _13451_ (.A(_06484_),
    .B(_06494_),
    .X(_06602_));
 sky130_fd_sc_hd__nor3_4 _13452_ (.A(_06602_),
    .B(_06506_),
    .C(_06514_),
    .Y(_06603_));
 sky130_fd_sc_hd__mux2_1 _13453_ (.A0(_06598_),
    .A1(_06601_),
    .S(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(_06406_),
    .A1(_06408_),
    .S(_06553_),
    .X(_06605_));
 sky130_fd_sc_hd__mux2_1 _13455_ (.A0(_06532_),
    .A1(_06588_),
    .S(_06553_),
    .X(_06606_));
 sky130_fd_sc_hd__mux2_2 _13456_ (.A0(_06605_),
    .A1(_06606_),
    .S(_06587_),
    .X(_06607_));
 sky130_fd_sc_hd__mux4_1 _13457_ (.A0(_06471_),
    .A1(_06475_),
    .A2(_06477_),
    .A3(_06480_),
    .S0(_06587_),
    .S1(_06554_),
    .X(_06608_));
 sky130_fd_sc_hd__inv_2 _13458_ (.A(_06371_),
    .Y(_06609_));
 sky130_fd_sc_hd__mux4_1 _13459_ (.A0(_06609_),
    .A1(_06574_),
    .A2(_06525_),
    .A3(_06492_),
    .S0(_06553_),
    .S1(_06587_),
    .X(_06610_));
 sky130_fd_sc_hd__nand2_1 _13460_ (.A(_06548_),
    .B(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__nor2_8 _13461_ (.A(_06460_),
    .B(_06544_),
    .Y(_06612_));
 sky130_fd_sc_hd__o211a_1 _13462_ (.A1(_06548_),
    .A2(_06608_),
    .B1(_06611_),
    .C1(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__a211oi_4 _13463_ (.A1(_06595_),
    .A2(_06604_),
    .B1(_06607_),
    .C1(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__xor2_2 _13464_ (.A(_06478_),
    .B(_06479_),
    .X(_06615_));
 sky130_fd_sc_hd__and3_1 _13465_ (.A(_06503_),
    .B(_06526_),
    .C(_06536_),
    .X(_06616_));
 sky130_fd_sc_hd__a211o_1 _13466_ (.A1(_06615_),
    .A2(_06552_),
    .B1(_06616_),
    .C1(_06546_),
    .X(_06617_));
 sky130_fd_sc_hd__a21boi_1 _13467_ (.A1(_06587_),
    .A2(_06600_),
    .B1_N(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__or2_1 _13468_ (.A(_06516_),
    .B(_06546_),
    .X(_06619_));
 sky130_fd_sc_hd__nor2_1 _13469_ (.A(_06489_),
    .B(_06553_),
    .Y(_06620_));
 sky130_fd_sc_hd__a211o_1 _13470_ (.A1(_06492_),
    .A2(_06553_),
    .B1(_06619_),
    .C1(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__nor2_1 _13471_ (.A(_06516_),
    .B(_06559_),
    .Y(_06622_));
 sky130_fd_sc_hd__mux2_1 _13472_ (.A0(_06471_),
    .A1(_06487_),
    .S(_06551_),
    .X(_06623_));
 sky130_fd_sc_hd__a21oi_1 _13473_ (.A1(_06622_),
    .A2(_06623_),
    .B1(_06523_),
    .Y(_06624_));
 sky130_fd_sc_hd__o211a_1 _13474_ (.A1(_06603_),
    .A2(_06618_),
    .B1(_06621_),
    .C1(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__mux2_2 _13475_ (.A0(_06597_),
    .A1(_06599_),
    .S(_06560_),
    .X(_06626_));
 sky130_fd_sc_hd__o21ai_1 _13476_ (.A1(_06577_),
    .A2(_06626_),
    .B1(_06461_),
    .Y(_06627_));
 sky130_fd_sc_hd__clkbuf_4 _13477_ (.A(_06570_),
    .X(_06628_));
 sky130_fd_sc_hd__nor2_1 _13478_ (.A(_06568_),
    .B(_06570_),
    .Y(_06629_));
 sky130_fd_sc_hd__a211o_1 _13479_ (.A1(_06609_),
    .A2(_06628_),
    .B1(_06566_),
    .C1(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__nor2_1 _13480_ (.A(_06548_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__a2bb2o_4 _13481_ (.A1_N(_06625_),
    .A2_N(_06627_),
    .B1(_06612_),
    .B2(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__a211o_1 _13482_ (.A1(_06475_),
    .A2(_06552_),
    .B1(_06561_),
    .C1(_06559_),
    .X(_06633_));
 sky130_fd_sc_hd__a211o_1 _13483_ (.A1(_06471_),
    .A2(_06552_),
    .B1(_06563_),
    .C1(_06546_),
    .X(_06634_));
 sky130_fd_sc_hd__a21o_1 _13484_ (.A1(_06633_),
    .A2(_06634_),
    .B1(_06603_),
    .X(_06635_));
 sky130_fd_sc_hd__nor2_1 _13485_ (.A(_06609_),
    .B(_06570_),
    .Y(_06636_));
 sky130_fd_sc_hd__a211o_1 _13486_ (.A1(_06568_),
    .A2(_06570_),
    .B1(_06619_),
    .C1(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__nand2_1 _13487_ (.A(_06603_),
    .B(_06546_),
    .Y(_06638_));
 sky130_fd_sc_hd__mux2_1 _13488_ (.A0(_06487_),
    .A1(_06489_),
    .S(_06552_),
    .X(_06639_));
 sky130_fd_sc_hd__or2_1 _13489_ (.A(_06638_),
    .B(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__a31o_1 _13490_ (.A1(_06635_),
    .A2(_06637_),
    .A3(_06640_),
    .B1(_06523_),
    .X(_06641_));
 sky130_fd_sc_hd__o21a_1 _13491_ (.A1(_06578_),
    .A2(_06586_),
    .B1(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__or2_1 _13492_ (.A(_06603_),
    .B(_06547_),
    .X(_06643_));
 sky130_fd_sc_hd__nand2_4 _13493_ (.A(_06643_),
    .B(_06543_),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_2 _13494_ (.A(_06612_),
    .B(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__mux2_1 _13495_ (.A0(_06525_),
    .A1(_06492_),
    .S(_06570_),
    .X(_06646_));
 sky130_fd_sc_hd__o2bb2a_1 _13496_ (.A1_N(_06587_),
    .A2_N(_06636_),
    .B1(_06646_),
    .B2(_06566_),
    .X(_06647_));
 sky130_fd_sc_hd__a21o_1 _13497_ (.A1(_06475_),
    .A2(_06552_),
    .B1(_06561_),
    .X(_06648_));
 sky130_fd_sc_hd__mux2_1 _13498_ (.A0(_06580_),
    .A1(_06648_),
    .S(_06560_),
    .X(_06649_));
 sky130_fd_sc_hd__a21o_1 _13499_ (.A1(_06471_),
    .A2(_06552_),
    .B1(_06563_),
    .X(_06650_));
 sky130_fd_sc_hd__a221o_1 _13500_ (.A1(_06622_),
    .A2(_06650_),
    .B1(_06639_),
    .B2(_06573_),
    .C1(_06523_),
    .X(_06651_));
 sky130_fd_sc_hd__a21o_1 _13501_ (.A1(_06585_),
    .A2(_06649_),
    .B1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__mux2_1 _13502_ (.A0(_06579_),
    .A1(_06583_),
    .S(_06546_),
    .X(_06653_));
 sky130_fd_sc_hd__o21a_1 _13503_ (.A1(_06585_),
    .A2(_06653_),
    .B1(_06460_),
    .X(_06654_));
 sky130_fd_sc_hd__a2bb2o_2 _13504_ (.A1_N(_06645_),
    .A2_N(_06647_),
    .B1(_06652_),
    .B2(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__a21o_4 _13505_ (.A1(_06632_),
    .A2(_06642_),
    .B1(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__a32o_1 _13506_ (.A1(_06585_),
    .A2(_06560_),
    .A3(_06636_),
    .B1(_06571_),
    .B2(_06644_),
    .X(_06657_));
 sky130_fd_sc_hd__o21ai_1 _13507_ (.A1(_06577_),
    .A2(_06584_),
    .B1(_06461_),
    .Y(_06658_));
 sky130_fd_sc_hd__a31o_1 _13508_ (.A1(_06603_),
    .A2(_06633_),
    .A3(_06634_),
    .B1(_06523_),
    .X(_06659_));
 sky130_fd_sc_hd__a21oi_1 _13509_ (.A1(_06585_),
    .A2(_06581_),
    .B1(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__o2bb2a_4 _13510_ (.A1_N(_06467_),
    .A2_N(_06657_),
    .B1(_06658_),
    .B2(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__a21oi_1 _13511_ (.A1(_06615_),
    .A2(_06552_),
    .B1(_06616_),
    .Y(_06662_));
 sky130_fd_sc_hd__a221o_1 _13512_ (.A1(_06622_),
    .A2(_06662_),
    .B1(_06623_),
    .B2(_06573_),
    .C1(_06523_),
    .X(_06663_));
 sky130_fd_sc_hd__a21oi_1 _13513_ (.A1(_06516_),
    .A2(_06601_),
    .B1(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nor2_1 _13514_ (.A(_06577_),
    .B(_06598_),
    .Y(_06665_));
 sky130_fd_sc_hd__o32a_1 _13515_ (.A1(_06467_),
    .A2(_06664_),
    .A3(_06665_),
    .B1(_06645_),
    .B2(_06610_),
    .X(_06666_));
 sky130_fd_sc_hd__buf_4 _13516_ (.A(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__nor2_4 _13517_ (.A(_06661_),
    .B(_06667_),
    .Y(_06668_));
 sky130_fd_sc_hd__buf_4 _13518_ (.A(_06467_),
    .X(_06669_));
 sky130_fd_sc_hd__nand2_1 _13519_ (.A(_06585_),
    .B(_06626_),
    .Y(_06670_));
 sky130_fd_sc_hd__o211a_1 _13520_ (.A1(_06585_),
    .A2(_06618_),
    .B1(_06670_),
    .C1(_06578_),
    .X(_06671_));
 sky130_fd_sc_hd__mux2_1 _13521_ (.A0(_06605_),
    .A1(_06596_),
    .S(_06560_),
    .X(_06672_));
 sky130_fd_sc_hd__nor2_1 _13522_ (.A(_06577_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__mux4_2 _13523_ (.A0(_06529_),
    .A1(_06574_),
    .A2(_06525_),
    .A3(_06615_),
    .S0(_06553_),
    .S1(_06560_),
    .X(_06674_));
 sky130_fd_sc_hd__o32a_1 _13524_ (.A1(_06461_),
    .A2(_06644_),
    .A3(_06630_),
    .B1(_06674_),
    .B2(_06645_),
    .X(_06675_));
 sky130_fd_sc_hd__o31ai_4 _13525_ (.A1(_06669_),
    .A2(_06671_),
    .A3(_06673_),
    .B1(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__mux2_1 _13526_ (.A0(_06649_),
    .A1(_06653_),
    .S(_06585_),
    .X(_06677_));
 sky130_fd_sc_hd__a22o_2 _13527_ (.A1(_06582_),
    .A2(_06573_),
    .B1(_06622_),
    .B2(_06589_),
    .X(_06678_));
 sky130_fd_sc_hd__mux4_1 _13528_ (.A0(_06471_),
    .A1(_06475_),
    .A2(_06480_),
    .A3(_06487_),
    .S0(_06560_),
    .S1(_06628_),
    .X(_06679_));
 sky130_fd_sc_hd__nor2_1 _13529_ (.A(_06548_),
    .B(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__a211oi_4 _13530_ (.A1(_06548_),
    .A2(_06647_),
    .B1(_06680_),
    .C1(_06556_),
    .Y(_06681_));
 sky130_fd_sc_hd__a211o_4 _13531_ (.A1(_06595_),
    .A2(_06677_),
    .B1(_06678_),
    .C1(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__a31o_1 _13532_ (.A1(_06656_),
    .A2(_06668_),
    .A3(_06676_),
    .B1(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__or3b_1 _13533_ (.A(_06594_),
    .B(_06614_),
    .C_N(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__buf_2 _13534_ (.A(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__nor2_2 _13535_ (.A(_06461_),
    .B(_06644_),
    .Y(_06686_));
 sky130_fd_sc_hd__buf_2 _13536_ (.A(_06560_),
    .X(_06687_));
 sky130_fd_sc_hd__o21ai_1 _13537_ (.A1(_06533_),
    .A2(_06628_),
    .B1(_06461_),
    .Y(_06688_));
 sky130_fd_sc_hd__a221o_1 _13538_ (.A1(_06687_),
    .A2(_06606_),
    .B1(_06672_),
    .B2(_06585_),
    .C1(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__a31oi_4 _13539_ (.A1(_06517_),
    .A2(_06519_),
    .A3(_06626_),
    .B1(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__mux4_1 _13540_ (.A0(_06473_),
    .A1(_06475_),
    .A2(_06477_),
    .A3(_06464_),
    .S0(_06560_),
    .S1(_06554_),
    .X(_06691_));
 sky130_fd_sc_hd__o22ai_2 _13541_ (.A1(_06575_),
    .A2(_06631_),
    .B1(_06691_),
    .B2(_06645_),
    .Y(_06692_));
 sky130_fd_sc_hd__a211oi_4 _13542_ (.A1(_06686_),
    .A2(_06674_),
    .B1(_06690_),
    .C1(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__clkbuf_4 _13543_ (.A(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__xnor2_1 _13544_ (.A(_06685_),
    .B(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__buf_2 _13545_ (.A(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__clkbuf_4 _13546_ (.A(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__buf_2 _13547_ (.A(_06593_),
    .X(_06698_));
 sky130_fd_sc_hd__a211o_2 _13548_ (.A1(_06595_),
    .A2(_06604_),
    .B1(_06607_),
    .C1(_06613_),
    .X(_06699_));
 sky130_fd_sc_hd__clkbuf_4 _13549_ (.A(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__buf_4 _13550_ (.A(_06683_),
    .X(_06701_));
 sky130_fd_sc_hd__a41o_2 _13551_ (.A1(_06698_),
    .A2(_06700_),
    .A3(_06701_),
    .A4(_06694_),
    .B1(_06484_),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_4 _13552_ (.A(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__nand2_8 _13553_ (.A(_06656_),
    .B(_06668_),
    .Y(_06704_));
 sky130_fd_sc_hd__a2bb2o_2 _13554_ (.A1_N(_06660_),
    .A2_N(_06658_),
    .B1(_06657_),
    .B2(_06669_),
    .X(_06705_));
 sky130_fd_sc_hd__o22a_1 _13555_ (.A1(_06645_),
    .A2(_06630_),
    .B1(_06625_),
    .B2(_06627_),
    .X(_06706_));
 sky130_fd_sc_hd__o21ai_4 _13556_ (.A1(_06578_),
    .A2(_06586_),
    .B1(_06641_),
    .Y(_06707_));
 sky130_fd_sc_hd__nor3_1 _13557_ (.A(_06706_),
    .B(_06707_),
    .C(_06667_),
    .Y(_06708_));
 sky130_fd_sc_hd__o2bb2a_2 _13558_ (.A1_N(_06652_),
    .A2_N(_06654_),
    .B1(_06645_),
    .B2(_06647_),
    .X(_06709_));
 sky130_fd_sc_hd__nor2_1 _13559_ (.A(_06709_),
    .B(_06667_),
    .Y(_06710_));
 sky130_fd_sc_hd__or3_2 _13560_ (.A(_06705_),
    .B(_06708_),
    .C(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__a21oi_2 _13561_ (.A1(_06704_),
    .A2(_06711_),
    .B1(_06614_),
    .Y(_06712_));
 sky130_fd_sc_hd__a211oi_4 _13562_ (.A1(_06595_),
    .A2(_06677_),
    .B1(_06678_),
    .C1(_06681_),
    .Y(_06713_));
 sky130_fd_sc_hd__xnor2_1 _13563_ (.A(_06656_),
    .B(_06667_),
    .Y(_06714_));
 sky130_fd_sc_hd__nor2_1 _13564_ (.A(_06713_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__xor2_4 _13565_ (.A(_06656_),
    .B(_06667_),
    .X(_06716_));
 sky130_fd_sc_hd__nand2_1 _13566_ (.A(_06700_),
    .B(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__a21o_1 _13567_ (.A1(_06704_),
    .A2(_06711_),
    .B1(_06713_),
    .X(_06718_));
 sky130_fd_sc_hd__nand2_1 _13568_ (.A(_06717_),
    .B(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__o31a_4 _13569_ (.A1(_06669_),
    .A2(_06671_),
    .A3(_06673_),
    .B1(_06675_),
    .X(_06720_));
 sky130_fd_sc_hd__nor2_4 _13570_ (.A(_06704_),
    .B(_06720_),
    .Y(_06721_));
 sky130_fd_sc_hd__a22o_1 _13571_ (.A1(_06712_),
    .A2(_06715_),
    .B1(_06719_),
    .B2(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__buf_2 _13572_ (.A(_06667_),
    .X(_06723_));
 sky130_fd_sc_hd__a21o_1 _13573_ (.A1(_06700_),
    .A2(_06701_),
    .B1(_06593_),
    .X(_06724_));
 sky130_fd_sc_hd__and2_1 _13574_ (.A(_06685_),
    .B(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__xnor2_2 _13575_ (.A(_06614_),
    .B(_06701_),
    .Y(_06726_));
 sky130_fd_sc_hd__nand4_4 _13576_ (.A(_06682_),
    .B(_06656_),
    .C(_06668_),
    .D(_06676_),
    .Y(_06727_));
 sky130_fd_sc_hd__and3_1 _13577_ (.A(_06705_),
    .B(_06701_),
    .C(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__or3b_1 _13578_ (.A(_06720_),
    .B(_06726_),
    .C_N(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__clkbuf_4 _13579_ (.A(_06676_),
    .X(_06730_));
 sky130_fd_sc_hd__xnor2_4 _13580_ (.A(_06699_),
    .B(_06701_),
    .Y(_06731_));
 sky130_fd_sc_hd__a32o_1 _13581_ (.A1(_06730_),
    .A2(_06701_),
    .A3(_06727_),
    .B1(_06731_),
    .B2(_06705_),
    .X(_06732_));
 sky130_fd_sc_hd__or4bb_1 _13582_ (.A(_06723_),
    .B(_06725_),
    .C_N(_06729_),
    .D_N(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__a2bb2o_1 _13583_ (.A1_N(_06723_),
    .A2_N(_06725_),
    .B1(_06729_),
    .B2(_06732_),
    .X(_06734_));
 sky130_fd_sc_hd__and3_1 _13584_ (.A(_06722_),
    .B(_06733_),
    .C(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__or3b_2 _13585_ (.A(_06667_),
    .B(_06726_),
    .C_N(_06728_),
    .X(_06736_));
 sky130_fd_sc_hd__nand2_1 _13586_ (.A(_06685_),
    .B(_06724_),
    .Y(_06737_));
 sky130_fd_sc_hd__clkbuf_4 _13587_ (.A(_06737_),
    .X(_06738_));
 sky130_fd_sc_hd__o21bai_1 _13588_ (.A1(_06667_),
    .A2(_06726_),
    .B1_N(_06728_),
    .Y(_06739_));
 sky130_fd_sc_hd__nand4_2 _13589_ (.A(_06655_),
    .B(_06738_),
    .C(_06736_),
    .D(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__a21oi_1 _13590_ (.A1(_06733_),
    .A2(_06734_),
    .B1(_06722_),
    .Y(_06741_));
 sky130_fd_sc_hd__a211o_1 _13591_ (.A1(_06736_),
    .A2(_06740_),
    .B1(_06741_),
    .C1(_06735_),
    .X(_06742_));
 sky130_fd_sc_hd__and2b_1 _13592_ (.A_N(_06735_),
    .B(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__or2_1 _13593_ (.A(_06709_),
    .B(_06702_),
    .X(_06744_));
 sky130_fd_sc_hd__clkbuf_4 _13594_ (.A(_06706_),
    .X(_06745_));
 sky130_fd_sc_hd__or2_1 _13595_ (.A(_06745_),
    .B(_06695_),
    .X(_06746_));
 sky130_fd_sc_hd__nor2_1 _13596_ (.A(_06723_),
    .B(_06696_),
    .Y(_06747_));
 sky130_fd_sc_hd__or3_1 _13597_ (.A(_06744_),
    .B(_06746_),
    .C(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__or2_1 _13598_ (.A(_06709_),
    .B(_06695_),
    .X(_06749_));
 sky130_fd_sc_hd__or2_1 _13599_ (.A(_06745_),
    .B(_06702_),
    .X(_06750_));
 sky130_fd_sc_hd__xor2_1 _13600_ (.A(_06744_),
    .B(_06747_),
    .X(_06751_));
 sky130_fd_sc_hd__o21ai_1 _13601_ (.A1(_06749_),
    .A2(_06750_),
    .B1(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__and2_1 _13602_ (.A(_06748_),
    .B(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__or2b_1 _13603_ (.A(_06743_),
    .B_N(_06753_),
    .X(_06754_));
 sky130_fd_sc_hd__clkbuf_4 _13604_ (.A(_06707_),
    .X(_06755_));
 sky130_fd_sc_hd__or4_1 _13605_ (.A(_06755_),
    .B(_06655_),
    .C(_06696_),
    .D(_06750_),
    .X(_06756_));
 sky130_fd_sc_hd__xnor2_1 _13606_ (.A(_06753_),
    .B(_06743_),
    .Y(_06757_));
 sky130_fd_sc_hd__or2b_1 _13607_ (.A(_06756_),
    .B_N(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__nand2_1 _13608_ (.A(_06754_),
    .B(_06758_),
    .Y(_06759_));
 sky130_fd_sc_hd__xnor2_1 _13609_ (.A(_06706_),
    .B(_06707_),
    .Y(_06760_));
 sky130_fd_sc_hd__buf_2 _13610_ (.A(_06760_),
    .X(_06761_));
 sky130_fd_sc_hd__or3_1 _13611_ (.A(_06706_),
    .B(_06707_),
    .C(_06709_),
    .X(_06762_));
 sky130_fd_sc_hd__and2_1 _13612_ (.A(_06656_),
    .B(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__and4_1 _13613_ (.A(_06558_),
    .B(_06694_),
    .C(_06761_),
    .D(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__xnor2_1 _13614_ (.A(_06632_),
    .B(_06707_),
    .Y(_06765_));
 sky130_fd_sc_hd__o2bb2a_1 _13615_ (.A1_N(_06694_),
    .A2_N(_06763_),
    .B1(_06765_),
    .B2(_06484_),
    .X(_06766_));
 sky130_fd_sc_hd__or2_1 _13616_ (.A(_06764_),
    .B(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__clkbuf_4 _13617_ (.A(_06763_),
    .X(_06768_));
 sky130_fd_sc_hd__clkbuf_4 _13618_ (.A(_06642_),
    .X(_06769_));
 sky130_fd_sc_hd__mux2_1 _13619_ (.A0(_06769_),
    .A1(_06706_),
    .S(_06693_),
    .X(_06770_));
 sky130_fd_sc_hd__nand2_1 _13620_ (.A(_06769_),
    .B(_06693_),
    .Y(_06771_));
 sky130_fd_sc_hd__nor2_1 _13621_ (.A(_06745_),
    .B(_06771_),
    .Y(_06772_));
 sky130_fd_sc_hd__a31o_1 _13622_ (.A1(_06698_),
    .A2(_06768_),
    .A3(_06770_),
    .B1(_06772_),
    .X(_06773_));
 sky130_fd_sc_hd__xor2_2 _13623_ (.A(_06767_),
    .B(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__xnor2_4 _13624_ (.A(_06704_),
    .B(_06720_),
    .Y(_06775_));
 sky130_fd_sc_hd__nand2_1 _13625_ (.A(_06682_),
    .B(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__nand2_1 _13626_ (.A(_06698_),
    .B(_06716_),
    .Y(_06777_));
 sky130_fd_sc_hd__xnor2_2 _13627_ (.A(_06712_),
    .B(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__xor2_2 _13628_ (.A(_06776_),
    .B(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__xnor2_2 _13629_ (.A(_06774_),
    .B(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__nand2_1 _13630_ (.A(_06698_),
    .B(_06763_),
    .Y(_06781_));
 sky130_fd_sc_hd__xor2_1 _13631_ (.A(_06781_),
    .B(_06770_),
    .X(_06782_));
 sky130_fd_sc_hd__nand2_1 _13632_ (.A(_06700_),
    .B(_06768_),
    .Y(_06783_));
 sky130_fd_sc_hd__nand2_1 _13633_ (.A(_06593_),
    .B(_06760_),
    .Y(_06784_));
 sky130_fd_sc_hd__xnor2_1 _13634_ (.A(_06771_),
    .B(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__nor2_1 _13635_ (.A(_06771_),
    .B(_06784_),
    .Y(_06786_));
 sky130_fd_sc_hd__o21ba_1 _13636_ (.A1(_06783_),
    .A2(_06785_),
    .B1_N(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__xor2_1 _13637_ (.A(_06782_),
    .B(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__xnor2_1 _13638_ (.A(_06717_),
    .B(_06718_),
    .Y(_06789_));
 sky130_fd_sc_hd__xnor2_1 _13639_ (.A(_06721_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__nor2_1 _13640_ (.A(_06782_),
    .B(_06787_),
    .Y(_06791_));
 sky130_fd_sc_hd__a21oi_1 _13641_ (.A1(_06788_),
    .A2(_06790_),
    .B1(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__xor2_1 _13642_ (.A(_06780_),
    .B(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__nand2_1 _13643_ (.A(_06736_),
    .B(_06740_),
    .Y(_06794_));
 sky130_fd_sc_hd__o21bai_1 _13644_ (.A1(_06735_),
    .A2(_06741_),
    .B1_N(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand3_1 _13645_ (.A(_06742_),
    .B(_06793_),
    .C(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__o21ai_2 _13646_ (.A1(_06780_),
    .A2(_06792_),
    .B1(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__nand2_1 _13647_ (.A(_06656_),
    .B(_06762_),
    .Y(_06798_));
 sky130_fd_sc_hd__clkbuf_4 _13648_ (.A(_06798_),
    .X(_06799_));
 sky130_fd_sc_hd__nor2_1 _13649_ (.A(_06799_),
    .B(_06764_),
    .Y(_06800_));
 sky130_fd_sc_hd__nand2_1 _13650_ (.A(_06700_),
    .B(_06775_),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_2 _13651_ (.A(_06704_),
    .B(_06711_),
    .Y(_06802_));
 sky130_fd_sc_hd__nand2_1 _13652_ (.A(_06698_),
    .B(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(_06694_),
    .B(_06716_),
    .Y(_06804_));
 sky130_fd_sc_hd__xor2_1 _13654_ (.A(_06803_),
    .B(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__xnor2_2 _13655_ (.A(_06801_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__xnor2_2 _13656_ (.A(_06800_),
    .B(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__or2b_1 _13657_ (.A(_06767_),
    .B_N(_06773_),
    .X(_06808_));
 sky130_fd_sc_hd__o21ai_2 _13658_ (.A1(_06774_),
    .A2(_06779_),
    .B1(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__xor2_1 _13659_ (.A(_06807_),
    .B(_06809_),
    .X(_06810_));
 sky130_fd_sc_hd__nand2_1 _13660_ (.A(_06729_),
    .B(_06733_),
    .Y(_06811_));
 sky130_fd_sc_hd__nor2_1 _13661_ (.A(_06717_),
    .B(_06803_),
    .Y(_06812_));
 sky130_fd_sc_hd__a31o_1 _13662_ (.A1(_06682_),
    .A2(_06775_),
    .A3(_06778_),
    .B1(_06812_),
    .X(_06813_));
 sky130_fd_sc_hd__nor2_1 _13663_ (.A(_06661_),
    .B(_06725_),
    .Y(_06814_));
 sky130_fd_sc_hd__nand2_1 _13664_ (.A(_06730_),
    .B(_06731_),
    .Y(_06815_));
 sky130_fd_sc_hd__or2_1 _13665_ (.A(_06713_),
    .B(_06721_),
    .X(_06816_));
 sky130_fd_sc_hd__xor2_1 _13666_ (.A(_06815_),
    .B(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__xnor2_1 _13667_ (.A(_06814_),
    .B(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__xnor2_1 _13668_ (.A(_06813_),
    .B(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__xnor2_1 _13669_ (.A(_06811_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__xor2_1 _13670_ (.A(_06810_),
    .B(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__xnor2_1 _13671_ (.A(_06797_),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__xor2_1 _13672_ (.A(_06756_),
    .B(_06757_),
    .X(_06823_));
 sky130_fd_sc_hd__nor2_1 _13673_ (.A(_06822_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__a21oi_1 _13674_ (.A1(_06797_),
    .A2(_06821_),
    .B1(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__or2b_1 _13675_ (.A(_06807_),
    .B_N(_06809_),
    .X(_06826_));
 sky130_fd_sc_hd__o21ai_1 _13676_ (.A1(_06810_),
    .A2(_06820_),
    .B1(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__and2_1 _13677_ (.A(_06694_),
    .B(_06802_),
    .X(_06828_));
 sky130_fd_sc_hd__nand2_1 _13678_ (.A(_06558_),
    .B(_06716_),
    .Y(_06829_));
 sky130_fd_sc_hd__xnor2_1 _13679_ (.A(_06828_),
    .B(_06829_),
    .Y(_06830_));
 sky130_fd_sc_hd__and2_1 _13680_ (.A(_06704_),
    .B(_06720_),
    .X(_06831_));
 sky130_fd_sc_hd__nor2_4 _13681_ (.A(_06721_),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nor2_1 _13682_ (.A(_06594_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__xor2_1 _13683_ (.A(_06830_),
    .B(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__a21oi_2 _13684_ (.A1(_06768_),
    .A2(_06806_),
    .B1(_06764_),
    .Y(_06835_));
 sky130_fd_sc_hd__xnor2_1 _13685_ (.A(_06834_),
    .B(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__nand2_1 _13686_ (.A(_06814_),
    .B(_06817_),
    .Y(_06837_));
 sky130_fd_sc_hd__o21ai_1 _13687_ (.A1(_06815_),
    .A2(_06816_),
    .B1(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__or2_1 _13688_ (.A(_06803_),
    .B(_06804_),
    .X(_06839_));
 sky130_fd_sc_hd__or2b_1 _13689_ (.A(_06801_),
    .B_N(_06805_),
    .X(_06840_));
 sky130_fd_sc_hd__o2bb2a_1 _13690_ (.A1_N(_06700_),
    .A2_N(_06721_),
    .B1(_06725_),
    .B2(_06720_),
    .X(_06841_));
 sky130_fd_sc_hd__a31o_1 _13691_ (.A1(_06700_),
    .A2(_06721_),
    .A3(_06738_),
    .B1(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__a21oi_1 _13692_ (.A1(_06839_),
    .A2(_06840_),
    .B1(_06842_),
    .Y(_06843_));
 sky130_fd_sc_hd__and3_1 _13693_ (.A(_06839_),
    .B(_06840_),
    .C(_06842_),
    .X(_06844_));
 sky130_fd_sc_hd__or2_1 _13694_ (.A(_06843_),
    .B(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__xnor2_1 _13695_ (.A(_06838_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__xnor2_1 _13696_ (.A(_06836_),
    .B(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__xor2_1 _13697_ (.A(_06827_),
    .B(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__and2b_1 _13698_ (.A_N(_06818_),
    .B(_06813_),
    .X(_06849_));
 sky130_fd_sc_hd__a21o_1 _13699_ (.A1(_06811_),
    .A2(_06819_),
    .B1(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__or2_1 _13700_ (.A(_06723_),
    .B(_06702_),
    .X(_06851_));
 sky130_fd_sc_hd__or2_1 _13701_ (.A(_06749_),
    .B(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__nor2_1 _13702_ (.A(_06661_),
    .B(_06696_),
    .Y(_06853_));
 sky130_fd_sc_hd__xnor2_1 _13703_ (.A(_06851_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__xnor2_1 _13704_ (.A(_06852_),
    .B(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__xnor2_1 _13705_ (.A(_06850_),
    .B(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__or2_1 _13706_ (.A(_06748_),
    .B(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__nand2_1 _13707_ (.A(_06748_),
    .B(_06856_),
    .Y(_06858_));
 sky130_fd_sc_hd__nand2_1 _13708_ (.A(_06857_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__xor2_1 _13709_ (.A(_06848_),
    .B(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__xnor2_1 _13710_ (.A(_06825_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__xnor2_1 _13711_ (.A(_06759_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__xnor2_1 _13712_ (.A(_06788_),
    .B(_06790_),
    .Y(_06863_));
 sky130_fd_sc_hd__xnor2_1 _13713_ (.A(_06783_),
    .B(_06785_),
    .Y(_06864_));
 sky130_fd_sc_hd__or4b_1 _13714_ (.A(_06614_),
    .B(_06755_),
    .C(_06765_),
    .D_N(_06593_),
    .X(_06865_));
 sky130_fd_sc_hd__a22o_1 _13715_ (.A1(_06593_),
    .A2(_06769_),
    .B1(_06761_),
    .B2(_06700_),
    .X(_06866_));
 sky130_fd_sc_hd__nand4_1 _13716_ (.A(_06682_),
    .B(_06768_),
    .C(_06865_),
    .D(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__nand2_1 _13717_ (.A(_06865_),
    .B(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__xnor2_1 _13718_ (.A(_06864_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand2_1 _13719_ (.A(_06705_),
    .B(_06775_),
    .Y(_06870_));
 sky130_fd_sc_hd__a21o_1 _13720_ (.A1(_06704_),
    .A2(_06711_),
    .B1(_06720_),
    .X(_06871_));
 sky130_fd_sc_hd__xnor2_1 _13721_ (.A(_06715_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__xnor2_1 _13722_ (.A(_06870_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__and2b_1 _13723_ (.A_N(_06864_),
    .B(_06868_),
    .X(_06874_));
 sky130_fd_sc_hd__a21o_1 _13724_ (.A1(_06869_),
    .A2(_06873_),
    .B1(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__and2b_1 _13725_ (.A_N(_06863_),
    .B(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__xnor2_1 _13726_ (.A(_06863_),
    .B(_06875_),
    .Y(_06877_));
 sky130_fd_sc_hd__and3_1 _13727_ (.A(_06655_),
    .B(_06701_),
    .C(_06727_),
    .X(_06878_));
 sky130_fd_sc_hd__or3b_1 _13728_ (.A(_06667_),
    .B(_06726_),
    .C_N(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__nand2_4 _13729_ (.A(_06701_),
    .B(_06727_),
    .Y(_06880_));
 sky130_fd_sc_hd__o22ai_1 _13730_ (.A1(_06709_),
    .A2(_06726_),
    .B1(_06880_),
    .B2(_06723_),
    .Y(_06881_));
 sky130_fd_sc_hd__nand4_1 _13731_ (.A(_06632_),
    .B(_06738_),
    .C(_06879_),
    .D(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__nand2_1 _13732_ (.A(_06879_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__and3_1 _13733_ (.A(_06730_),
    .B(_06802_),
    .C(_06715_),
    .X(_06884_));
 sky130_fd_sc_hd__a31o_1 _13734_ (.A1(_06705_),
    .A2(_06775_),
    .A3(_06872_),
    .B1(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__a22o_1 _13735_ (.A1(_06655_),
    .A2(_06737_),
    .B1(_06736_),
    .B2(_06739_),
    .X(_06886_));
 sky130_fd_sc_hd__nand3_1 _13736_ (.A(_06740_),
    .B(_06885_),
    .C(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__a21o_1 _13737_ (.A1(_06740_),
    .A2(_06886_),
    .B1(_06885_),
    .X(_06888_));
 sky130_fd_sc_hd__nand3_1 _13738_ (.A(_06883_),
    .B(_06887_),
    .C(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__a21o_1 _13739_ (.A1(_06887_),
    .A2(_06888_),
    .B1(_06883_),
    .X(_06890_));
 sky130_fd_sc_hd__and3_1 _13740_ (.A(_06877_),
    .B(_06889_),
    .C(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__a21o_1 _13741_ (.A1(_06742_),
    .A2(_06795_),
    .B1(_06793_),
    .X(_06892_));
 sky130_fd_sc_hd__o211a_1 _13742_ (.A1(_06876_),
    .A2(_06891_),
    .B1(_06892_),
    .C1(_06796_),
    .X(_06893_));
 sky130_fd_sc_hd__a211oi_2 _13743_ (.A1(_06796_),
    .A2(_06892_),
    .B1(_06891_),
    .C1(_06876_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand2_1 _13744_ (.A(_06887_),
    .B(_06889_),
    .Y(_06895_));
 sky130_fd_sc_hd__or2_1 _13745_ (.A(_06755_),
    .B(_06695_),
    .X(_06896_));
 sky130_fd_sc_hd__or2_1 _13746_ (.A(_06750_),
    .B(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__xor2_1 _13747_ (.A(_06749_),
    .B(_06750_),
    .X(_06898_));
 sky130_fd_sc_hd__xnor2_1 _13748_ (.A(_06897_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__xnor2_1 _13749_ (.A(_06895_),
    .B(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__or3_1 _13750_ (.A(_06893_),
    .B(_06894_),
    .C(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__and2b_1 _13751_ (.A_N(_06893_),
    .B(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__xnor2_1 _13752_ (.A(_06822_),
    .B(_06823_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand2_1 _13753_ (.A(_06895_),
    .B(_06899_),
    .Y(_06904_));
 sky130_fd_sc_hd__xor2_1 _13754_ (.A(_06902_),
    .B(_06903_),
    .X(_06905_));
 sky130_fd_sc_hd__or2b_1 _13755_ (.A(_06904_),
    .B_N(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__o21a_1 _13756_ (.A1(_06902_),
    .A2(_06903_),
    .B1(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__xnor2_1 _13757_ (.A(_06862_),
    .B(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__a22o_1 _13758_ (.A1(_06682_),
    .A2(_06768_),
    .B1(_06865_),
    .B2(_06866_),
    .X(_06909_));
 sky130_fd_sc_hd__a22o_1 _13759_ (.A1(_06699_),
    .A2(_06769_),
    .B1(_06761_),
    .B2(_06682_),
    .X(_06910_));
 sky130_fd_sc_hd__nor2_1 _13760_ (.A(_06713_),
    .B(_06755_),
    .Y(_06911_));
 sky130_fd_sc_hd__and3_1 _13761_ (.A(_06699_),
    .B(_06761_),
    .C(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__a31o_1 _13762_ (.A1(_06730_),
    .A2(_06768_),
    .A3(_06910_),
    .B1(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__nand3_1 _13763_ (.A(_06867_),
    .B(_06909_),
    .C(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__a21o_1 _13764_ (.A1(_06867_),
    .A2(_06909_),
    .B1(_06913_),
    .X(_06915_));
 sky130_fd_sc_hd__nand2_1 _13765_ (.A(_06914_),
    .B(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__mux2_1 _13766_ (.A0(_06723_),
    .A1(_06714_),
    .S(_06730_),
    .X(_06917_));
 sky130_fd_sc_hd__xnor2_1 _13767_ (.A(_06916_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__and2b_1 _13768_ (.A_N(_06912_),
    .B(_06910_),
    .X(_06919_));
 sky130_fd_sc_hd__or3b_1 _13769_ (.A(_06720_),
    .B(_06798_),
    .C_N(_06919_),
    .X(_06920_));
 sky130_fd_sc_hd__a21o_1 _13770_ (.A1(_06730_),
    .A2(_06768_),
    .B1(_06919_),
    .X(_06921_));
 sky130_fd_sc_hd__nor2_1 _13771_ (.A(_06661_),
    .B(_06798_),
    .Y(_06922_));
 sky130_fd_sc_hd__and3_1 _13772_ (.A(_06676_),
    .B(_06761_),
    .C(_06911_),
    .X(_06923_));
 sky130_fd_sc_hd__a21oi_1 _13773_ (.A1(_06730_),
    .A2(_06761_),
    .B1(_06911_),
    .Y(_06924_));
 sky130_fd_sc_hd__nor2_1 _13774_ (.A(_06923_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__a21o_1 _13775_ (.A1(_06922_),
    .A2(_06925_),
    .B1(_06923_),
    .X(_06926_));
 sky130_fd_sc_hd__a21oi_1 _13776_ (.A1(_06920_),
    .A2(_06921_),
    .B1(_06926_),
    .Y(_06927_));
 sky130_fd_sc_hd__a211o_1 _13777_ (.A1(_06661_),
    .A2(_06723_),
    .B1(_06668_),
    .C1(_06656_),
    .X(_06928_));
 sky130_fd_sc_hd__o21a_1 _13778_ (.A1(_06709_),
    .A2(_06832_),
    .B1(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__and3_1 _13779_ (.A(_06920_),
    .B(_06921_),
    .C(_06926_),
    .X(_06930_));
 sky130_fd_sc_hd__o21bai_1 _13780_ (.A1(_06927_),
    .A2(_06929_),
    .B1_N(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__or2b_1 _13781_ (.A(_06918_),
    .B_N(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__xnor2_1 _13782_ (.A(_06918_),
    .B(_06931_),
    .Y(_06933_));
 sky130_fd_sc_hd__inv_2 _13783_ (.A(_06704_),
    .Y(_06934_));
 sky130_fd_sc_hd__or3b_2 _13784_ (.A(_06745_),
    .B(_06726_),
    .C_N(_06878_),
    .X(_06935_));
 sky130_fd_sc_hd__a21o_1 _13785_ (.A1(_06632_),
    .A2(_06731_),
    .B1(_06878_),
    .X(_06936_));
 sky130_fd_sc_hd__nand4_2 _13786_ (.A(_06769_),
    .B(_06738_),
    .C(_06935_),
    .D(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__a22o_1 _13787_ (.A1(_06769_),
    .A2(_06738_),
    .B1(_06935_),
    .B2(_06936_),
    .X(_06938_));
 sky130_fd_sc_hd__and3_1 _13788_ (.A(_06934_),
    .B(_06937_),
    .C(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__a21oi_1 _13789_ (.A1(_06937_),
    .A2(_06938_),
    .B1(_06934_),
    .Y(_06940_));
 sky130_fd_sc_hd__nor2_1 _13790_ (.A(_06745_),
    .B(_06880_),
    .Y(_06941_));
 sky130_fd_sc_hd__clkbuf_4 _13791_ (.A(_06726_),
    .X(_06942_));
 sky130_fd_sc_hd__nor2_1 _13792_ (.A(_06755_),
    .B(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__and2_1 _13793_ (.A(_06941_),
    .B(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__inv_2 _13794_ (.A(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__or3_1 _13795_ (.A(_06939_),
    .B(_06940_),
    .C(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__o21ai_1 _13796_ (.A1(_06939_),
    .A2(_06940_),
    .B1(_06945_),
    .Y(_06947_));
 sky130_fd_sc_hd__nand3_1 _13797_ (.A(_06933_),
    .B(_06946_),
    .C(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__a22o_1 _13798_ (.A1(_06632_),
    .A2(_06738_),
    .B1(_06879_),
    .B2(_06881_),
    .X(_06949_));
 sky130_fd_sc_hd__a21oi_1 _13799_ (.A1(_06882_),
    .A2(_06949_),
    .B1(_06721_),
    .Y(_06950_));
 sky130_fd_sc_hd__and3_1 _13800_ (.A(_06721_),
    .B(_06882_),
    .C(_06949_),
    .X(_06951_));
 sky130_fd_sc_hd__a211o_1 _13801_ (.A1(_06935_),
    .A2(_06937_),
    .B1(_06950_),
    .C1(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__nand2_1 _13802_ (.A(_06935_),
    .B(_06937_),
    .Y(_06953_));
 sky130_fd_sc_hd__o21bai_1 _13803_ (.A1(_06951_),
    .A2(_06950_),
    .B1_N(_06953_),
    .Y(_06954_));
 sky130_fd_sc_hd__xnor2_1 _13804_ (.A(_06869_),
    .B(_06873_),
    .Y(_06955_));
 sky130_fd_sc_hd__o21ai_1 _13805_ (.A1(_06916_),
    .A2(_06917_),
    .B1(_06914_),
    .Y(_06956_));
 sky130_fd_sc_hd__xnor2_1 _13806_ (.A(_06955_),
    .B(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__a21oi_1 _13807_ (.A1(_06952_),
    .A2(_06954_),
    .B1(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__and3_1 _13808_ (.A(_06952_),
    .B(_06957_),
    .C(_06954_),
    .X(_06959_));
 sky130_fd_sc_hd__a211oi_2 _13809_ (.A1(_06932_),
    .A2(_06948_),
    .B1(_06958_),
    .C1(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__o211a_1 _13810_ (.A1(_06959_),
    .A2(_06958_),
    .B1(_06948_),
    .C1(_06932_),
    .X(_06961_));
 sky130_fd_sc_hd__and2b_1 _13811_ (.A_N(_06939_),
    .B(_06946_),
    .X(_06962_));
 sky130_fd_sc_hd__xnor2_1 _13812_ (.A(_06896_),
    .B(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__nor3_1 _13813_ (.A(_06960_),
    .B(_06961_),
    .C(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__and2b_1 _13814_ (.A_N(_06955_),
    .B(_06956_),
    .X(_06965_));
 sky130_fd_sc_hd__a21o_1 _13815_ (.A1(_06889_),
    .A2(_06890_),
    .B1(_06877_),
    .X(_06966_));
 sky130_fd_sc_hd__nand3_1 _13816_ (.A(_06877_),
    .B(_06889_),
    .C(_06890_),
    .Y(_06967_));
 sky130_fd_sc_hd__o211a_1 _13817_ (.A1(_06965_),
    .A2(_06959_),
    .B1(_06966_),
    .C1(_06967_),
    .X(_06968_));
 sky130_fd_sc_hd__a211oi_2 _13818_ (.A1(_06967_),
    .A2(_06966_),
    .B1(_06959_),
    .C1(_06965_),
    .Y(_06969_));
 sky130_fd_sc_hd__a211oi_1 _13819_ (.A1(_06935_),
    .A2(_06937_),
    .B1(_06950_),
    .C1(_06951_),
    .Y(_06970_));
 sky130_fd_sc_hd__o21ai_1 _13820_ (.A1(_06755_),
    .A2(_06702_),
    .B1(_06746_),
    .Y(_06971_));
 sky130_fd_sc_hd__and2_1 _13821_ (.A(_06897_),
    .B(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__o21ai_1 _13822_ (.A1(_06951_),
    .A2(_06970_),
    .B1(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__or3_1 _13823_ (.A(_06951_),
    .B(_06970_),
    .C(_06972_),
    .X(_06974_));
 sky130_fd_sc_hd__nand2_1 _13824_ (.A(_06973_),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__o21ai_1 _13825_ (.A1(_06968_),
    .A2(_06969_),
    .B1(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__or3_1 _13826_ (.A(_06968_),
    .B(_06969_),
    .C(_06975_),
    .X(_06977_));
 sky130_fd_sc_hd__o211a_1 _13827_ (.A1(_06960_),
    .A2(_06964_),
    .B1(_06976_),
    .C1(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__or2_1 _13828_ (.A(_06896_),
    .B(_06962_),
    .X(_06979_));
 sky130_fd_sc_hd__a211oi_1 _13829_ (.A1(_06977_),
    .A2(_06976_),
    .B1(_06964_),
    .C1(_06960_),
    .Y(_06980_));
 sky130_fd_sc_hd__nor3_1 _13830_ (.A(_06979_),
    .B(_06978_),
    .C(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__nor3_1 _13831_ (.A(_06968_),
    .B(_06969_),
    .C(_06975_),
    .Y(_06982_));
 sky130_fd_sc_hd__o21ai_1 _13832_ (.A1(_06893_),
    .A2(_06894_),
    .B1(_06900_),
    .Y(_06983_));
 sky130_fd_sc_hd__o211a_1 _13833_ (.A1(_06968_),
    .A2(_06982_),
    .B1(_06983_),
    .C1(_06901_),
    .X(_06984_));
 sky130_fd_sc_hd__a211oi_1 _13834_ (.A1(_06901_),
    .A2(_06983_),
    .B1(_06982_),
    .C1(_06968_),
    .Y(_06985_));
 sky130_fd_sc_hd__or3_1 _13835_ (.A(_06973_),
    .B(_06984_),
    .C(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__o21ai_1 _13836_ (.A1(_06984_),
    .A2(_06985_),
    .B1(_06973_),
    .Y(_06987_));
 sky130_fd_sc_hd__o211ai_2 _13837_ (.A1(_06978_),
    .A2(_06981_),
    .B1(_06986_),
    .C1(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__xnor2_1 _13838_ (.A(_06904_),
    .B(_06905_),
    .Y(_06989_));
 sky130_fd_sc_hd__and2b_1 _13839_ (.A_N(_06984_),
    .B(_06986_),
    .X(_06990_));
 sky130_fd_sc_hd__xor2_1 _13840_ (.A(_06989_),
    .B(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__or2_1 _13841_ (.A(_06988_),
    .B(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__o21ai_1 _13842_ (.A1(_06978_),
    .A2(_06980_),
    .B1(_06979_),
    .Y(_06993_));
 sky130_fd_sc_hd__and2b_1 _13843_ (.A_N(_06981_),
    .B(_06993_),
    .X(_06994_));
 sky130_fd_sc_hd__xnor2_1 _13844_ (.A(_06922_),
    .B(_06925_),
    .Y(_06995_));
 sky130_fd_sc_hd__nand2_1 _13845_ (.A(_06730_),
    .B(_06761_),
    .Y(_06996_));
 sky130_fd_sc_hd__nand2_1 _13846_ (.A(_06705_),
    .B(_06769_),
    .Y(_06997_));
 sky130_fd_sc_hd__or2_1 _13847_ (.A(_06667_),
    .B(_06798_),
    .X(_06998_));
 sky130_fd_sc_hd__a22o_1 _13848_ (.A1(_06769_),
    .A2(_06730_),
    .B1(_06761_),
    .B2(_06705_),
    .X(_06999_));
 sky130_fd_sc_hd__o21ai_1 _13849_ (.A1(_06996_),
    .A2(_06997_),
    .B1(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__o22a_1 _13850_ (.A1(_06996_),
    .A2(_06997_),
    .B1(_06998_),
    .B2(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__nor2_1 _13851_ (.A(_06995_),
    .B(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__nand2_1 _13852_ (.A(_06632_),
    .B(_06775_),
    .Y(_07003_));
 sky130_fd_sc_hd__mux2_1 _13853_ (.A0(_06661_),
    .A1(_06708_),
    .S(_06709_),
    .X(_07004_));
 sky130_fd_sc_hd__xnor2_1 _13854_ (.A(_07003_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__xor2_1 _13855_ (.A(_06995_),
    .B(_07001_),
    .X(_07006_));
 sky130_fd_sc_hd__and2_1 _13856_ (.A(_07005_),
    .B(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__nor2_1 _13857_ (.A(_06930_),
    .B(_06927_),
    .Y(_07008_));
 sky130_fd_sc_hd__xnor2_1 _13858_ (.A(_07008_),
    .B(_06929_),
    .Y(_07009_));
 sky130_fd_sc_hd__o21a_1 _13859_ (.A1(_07002_),
    .A2(_07007_),
    .B1(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__xnor2_1 _13860_ (.A(_06941_),
    .B(_06943_),
    .Y(_07011_));
 sky130_fd_sc_hd__a32oi_1 _13861_ (.A1(_06632_),
    .A2(_06775_),
    .A3(_07004_),
    .B1(_06655_),
    .B2(_06668_),
    .Y(_07012_));
 sky130_fd_sc_hd__or2_2 _13862_ (.A(_07011_),
    .B(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__nand2_1 _13863_ (.A(_07011_),
    .B(_07012_),
    .Y(_07014_));
 sky130_fd_sc_hd__nand2_1 _13864_ (.A(_07013_),
    .B(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__nor3_1 _13865_ (.A(_07009_),
    .B(_07002_),
    .C(_07007_),
    .Y(_07016_));
 sky130_fd_sc_hd__or3_1 _13866_ (.A(_07010_),
    .B(_07015_),
    .C(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__or2b_1 _13867_ (.A(_07010_),
    .B_N(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__a21o_1 _13868_ (.A1(_06946_),
    .A2(_06947_),
    .B1(_06933_),
    .X(_07019_));
 sky130_fd_sc_hd__and2_1 _13869_ (.A(_06948_),
    .B(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__nand2_1 _13870_ (.A(_07018_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__xnor2_1 _13871_ (.A(_07018_),
    .B(_07020_),
    .Y(_07022_));
 sky130_fd_sc_hd__or2_1 _13872_ (.A(_07013_),
    .B(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__o21a_1 _13873_ (.A1(_06960_),
    .A2(_06961_),
    .B1(_06963_),
    .X(_07024_));
 sky130_fd_sc_hd__a211oi_1 _13874_ (.A1(_07021_),
    .A2(_07023_),
    .B1(_06964_),
    .C1(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__a211o_1 _13875_ (.A1(_06986_),
    .A2(_06987_),
    .B1(_06978_),
    .C1(_06981_),
    .X(_07026_));
 sky130_fd_sc_hd__nand4_1 _13876_ (.A(_06988_),
    .B(_06994_),
    .C(_07025_),
    .D(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__a22o_1 _13877_ (.A1(_06994_),
    .A2(_07025_),
    .B1(_07026_),
    .B2(_06988_),
    .X(_07028_));
 sky130_fd_sc_hd__o211ai_1 _13878_ (.A1(_06964_),
    .A2(_07024_),
    .B1(_07021_),
    .C1(_07023_),
    .Y(_07029_));
 sky130_fd_sc_hd__and3b_1 _13879_ (.A_N(_07025_),
    .B(_07029_),
    .C(_06994_),
    .X(_07030_));
 sky130_fd_sc_hd__xor2_1 _13880_ (.A(_07013_),
    .B(_07022_),
    .X(_07031_));
 sky130_fd_sc_hd__o21ai_1 _13881_ (.A1(_07010_),
    .A2(_07016_),
    .B1(_07015_),
    .Y(_07032_));
 sky130_fd_sc_hd__nand2_1 _13882_ (.A(_07017_),
    .B(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__nor2_1 _13883_ (.A(_07005_),
    .B(_07006_),
    .Y(_07034_));
 sky130_fd_sc_hd__or2_1 _13884_ (.A(_07007_),
    .B(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__and2_1 _13885_ (.A(_06704_),
    .B(_06711_),
    .X(_07036_));
 sky130_fd_sc_hd__nor2_1 _13886_ (.A(_06745_),
    .B(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__xnor2_1 _13887_ (.A(_06710_),
    .B(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__nor2_1 _13888_ (.A(_06755_),
    .B(_06832_),
    .Y(_07039_));
 sky130_fd_sc_hd__xnor2_1 _13889_ (.A(_07038_),
    .B(_07039_),
    .Y(_07040_));
 sky130_fd_sc_hd__xor2_1 _13890_ (.A(_06998_),
    .B(_07000_),
    .X(_07041_));
 sky130_fd_sc_hd__nor2_4 _13891_ (.A(_06745_),
    .B(_06755_),
    .Y(_07042_));
 sky130_fd_sc_hd__or2_1 _13892_ (.A(_07042_),
    .B(_06709_),
    .X(_07043_));
 sky130_fd_sc_hd__clkbuf_4 _13893_ (.A(_06765_),
    .X(_07044_));
 sky130_fd_sc_hd__o21a_1 _13894_ (.A1(_06723_),
    .A2(_07044_),
    .B1(_06997_),
    .X(_07045_));
 sky130_fd_sc_hd__a2bb2o_1 _13895_ (.A1_N(_07043_),
    .A2_N(_07045_),
    .B1(_07042_),
    .B2(_06668_),
    .X(_07046_));
 sky130_fd_sc_hd__and2_1 _13896_ (.A(_07041_),
    .B(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__nor2_1 _13897_ (.A(_07041_),
    .B(_07046_),
    .Y(_07048_));
 sky130_fd_sc_hd__nor2_1 _13898_ (.A(_07047_),
    .B(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__a21oi_1 _13899_ (.A1(_07040_),
    .A2(_07049_),
    .B1(_07047_),
    .Y(_07050_));
 sky130_fd_sc_hd__clkbuf_4 _13900_ (.A(_06755_),
    .X(_07051_));
 sky130_fd_sc_hd__nor2_1 _13901_ (.A(_07051_),
    .B(_06880_),
    .Y(_07052_));
 sky130_fd_sc_hd__or3_1 _13902_ (.A(_06755_),
    .B(_06832_),
    .C(_07038_),
    .X(_07053_));
 sky130_fd_sc_hd__a21bo_1 _13903_ (.A1(_06710_),
    .A2(_07037_),
    .B1_N(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__xnor2_1 _13904_ (.A(_07052_),
    .B(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__xnor2_1 _13905_ (.A(_07035_),
    .B(_07050_),
    .Y(_07056_));
 sky130_fd_sc_hd__nor2_1 _13906_ (.A(_07055_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__o21ba_1 _13907_ (.A1(_07035_),
    .A2(_07050_),
    .B1_N(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__nand2_1 _13908_ (.A(_07052_),
    .B(_07054_),
    .Y(_07059_));
 sky130_fd_sc_hd__xnor2_1 _13909_ (.A(_07033_),
    .B(_07058_),
    .Y(_07060_));
 sky130_fd_sc_hd__or2_1 _13910_ (.A(_07059_),
    .B(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__o21ai_2 _13911_ (.A1(_07033_),
    .A2(_07058_),
    .B1(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__and2_1 _13912_ (.A(_07031_),
    .B(_07062_),
    .X(_07063_));
 sky130_fd_sc_hd__a22o_1 _13913_ (.A1(_07027_),
    .A2(_07028_),
    .B1(_07030_),
    .B2(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__xnor2_1 _13914_ (.A(_07040_),
    .B(_07049_),
    .Y(_07065_));
 sky130_fd_sc_hd__clkbuf_4 _13915_ (.A(_06714_),
    .X(_07066_));
 sky130_fd_sc_hd__o22a_1 _13916_ (.A1(_07051_),
    .A2(_07036_),
    .B1(_07066_),
    .B2(_06745_),
    .X(_07067_));
 sky130_fd_sc_hd__a211o_1 _13917_ (.A1(_07043_),
    .A2(_07045_),
    .B1(_07046_),
    .C1(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__o2bb2a_1 _13918_ (.A1_N(_06661_),
    .A2_N(_06708_),
    .B1(_07065_),
    .B2(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__and2_1 _13919_ (.A(_07055_),
    .B(_07056_),
    .X(_07070_));
 sky130_fd_sc_hd__o21ba_1 _13920_ (.A1(_07057_),
    .A2(_07070_),
    .B1_N(_07042_),
    .X(_07071_));
 sky130_fd_sc_hd__a211oi_2 _13921_ (.A1(_07059_),
    .A2(_07060_),
    .B1(_07069_),
    .C1(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__o211a_1 _13922_ (.A1(_07031_),
    .A2(_07062_),
    .B1(_07072_),
    .C1(_07030_),
    .X(_07073_));
 sky130_fd_sc_hd__and4_1 _13923_ (.A(_07027_),
    .B(_07028_),
    .C(_07030_),
    .D(_07063_),
    .X(_07074_));
 sky130_fd_sc_hd__a21o_1 _13924_ (.A1(_07064_),
    .A2(_07073_),
    .B1(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__nand2_1 _13925_ (.A(_06988_),
    .B(_07027_),
    .Y(_07076_));
 sky130_fd_sc_hd__xnor2_1 _13926_ (.A(_06991_),
    .B(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__a2bb2o_1 _13927_ (.A1_N(_06991_),
    .A2_N(_07027_),
    .B1(_07075_),
    .B2(_07077_),
    .X(_07078_));
 sky130_fd_sc_hd__and2b_1 _13928_ (.A_N(_06990_),
    .B(_06989_),
    .X(_07079_));
 sky130_fd_sc_hd__and2b_1 _13929_ (.A_N(_07079_),
    .B(_06992_),
    .X(_07080_));
 sky130_fd_sc_hd__xor2_1 _13930_ (.A(_06908_),
    .B(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__a2bb2o_1 _13931_ (.A1_N(_06908_),
    .A2_N(_06992_),
    .B1(_07078_),
    .B2(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__a21bo_1 _13932_ (.A1(_06850_),
    .A2(_06855_),
    .B1_N(_06857_),
    .X(_07083_));
 sky130_fd_sc_hd__or2b_1 _13933_ (.A(_06847_),
    .B_N(_06827_),
    .X(_07084_));
 sky130_fd_sc_hd__o21ai_1 _13934_ (.A1(_06848_),
    .A2(_06859_),
    .B1(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__or2b_1 _13935_ (.A(_06835_),
    .B_N(_06834_),
    .X(_07086_));
 sky130_fd_sc_hd__nand2_1 _13936_ (.A(_06836_),
    .B(_06846_),
    .Y(_07087_));
 sky130_fd_sc_hd__nand2_1 _13937_ (.A(_07086_),
    .B(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__nor2_1 _13938_ (.A(_06484_),
    .B(_06832_),
    .Y(_07089_));
 sky130_fd_sc_hd__nand2_1 _13939_ (.A(_06828_),
    .B(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__a22o_1 _13940_ (.A1(_06558_),
    .A2(_06802_),
    .B1(_06775_),
    .B2(_06694_),
    .X(_07091_));
 sky130_fd_sc_hd__and2_1 _13941_ (.A(_07090_),
    .B(_07091_),
    .X(_07092_));
 sky130_fd_sc_hd__a22o_1 _13942_ (.A1(_06716_),
    .A2(_06828_),
    .B1(_06830_),
    .B2(_06833_),
    .X(_07093_));
 sky130_fd_sc_hd__o2bb2a_1 _13943_ (.A1_N(_06698_),
    .A2_N(_06880_),
    .B1(_06725_),
    .B2(_06682_),
    .X(_07094_));
 sky130_fd_sc_hd__xnor2_1 _13944_ (.A(_07093_),
    .B(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__o311a_1 _13945_ (.A1(_06698_),
    .A2(_06704_),
    .A3(_06720_),
    .B1(_06701_),
    .C1(_06700_),
    .X(_07096_));
 sky130_fd_sc_hd__xnor2_1 _13946_ (.A(_07095_),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__and2_1 _13947_ (.A(_07092_),
    .B(_07097_),
    .X(_07098_));
 sky130_fd_sc_hd__nor2_1 _13948_ (.A(_07092_),
    .B(_07097_),
    .Y(_07099_));
 sky130_fd_sc_hd__or2_1 _13949_ (.A(_07098_),
    .B(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__xnor2_1 _13950_ (.A(_07088_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__or3_1 _13951_ (.A(_06749_),
    .B(_06851_),
    .C(_06853_),
    .X(_07102_));
 sky130_fd_sc_hd__and2b_1 _13952_ (.A_N(_06845_),
    .B(_06838_),
    .X(_07103_));
 sky130_fd_sc_hd__or2_1 _13953_ (.A(_06843_),
    .B(_07103_),
    .X(_07104_));
 sky130_fd_sc_hd__or2_1 _13954_ (.A(_06661_),
    .B(_06702_),
    .X(_07105_));
 sky130_fd_sc_hd__or3_1 _13955_ (.A(_06723_),
    .B(_06696_),
    .C(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__or2_2 _13956_ (.A(_06720_),
    .B(_06696_),
    .X(_07107_));
 sky130_fd_sc_hd__xor2_1 _13957_ (.A(_07105_),
    .B(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__xnor2_1 _13958_ (.A(_07106_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__xnor2_1 _13959_ (.A(_07104_),
    .B(_07109_),
    .Y(_07110_));
 sky130_fd_sc_hd__xor2_1 _13960_ (.A(_07102_),
    .B(_07110_),
    .X(_07111_));
 sky130_fd_sc_hd__xnor2_1 _13961_ (.A(_07101_),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__xor2_1 _13962_ (.A(_07085_),
    .B(_07112_),
    .X(_07113_));
 sky130_fd_sc_hd__xor2_1 _13963_ (.A(_07083_),
    .B(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__and2b_1 _13964_ (.A_N(_06825_),
    .B(_06860_),
    .X(_07115_));
 sky130_fd_sc_hd__a21oi_1 _13965_ (.A1(_06759_),
    .A2(_06861_),
    .B1(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__xnor2_1 _13966_ (.A(_07114_),
    .B(_07116_),
    .Y(_07117_));
 sky130_fd_sc_hd__or2b_1 _13967_ (.A(_06908_),
    .B_N(_07079_),
    .X(_07118_));
 sky130_fd_sc_hd__o21ai_1 _13968_ (.A1(_06862_),
    .A2(_06907_),
    .B1(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__xnor2_1 _13969_ (.A(_07117_),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__xnor2_1 _13970_ (.A(_07082_),
    .B(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__xor2_1 _13971_ (.A(_07078_),
    .B(_07081_),
    .X(_07122_));
 sky130_fd_sc_hd__xnor2_1 _13972_ (.A(_07075_),
    .B(_07077_),
    .Y(_07123_));
 sky130_fd_sc_hd__and2b_1 _13973_ (.A_N(_07074_),
    .B(_07064_),
    .X(_07124_));
 sky130_fd_sc_hd__xnor2_2 _13974_ (.A(_07124_),
    .B(_07073_),
    .Y(_07125_));
 sky130_fd_sc_hd__nor2_1 _13975_ (.A(_07123_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__nor2_1 _13976_ (.A(_07122_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_1 _13977_ (.A(_07121_),
    .B(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__a2bb2o_1 _13978_ (.A1_N(_07117_),
    .A2_N(_07118_),
    .B1(_07120_),
    .B2(_07082_),
    .X(_07129_));
 sky130_fd_sc_hd__and2b_1 _13979_ (.A_N(_07112_),
    .B(_07085_),
    .X(_07130_));
 sky130_fd_sc_hd__and2b_1 _13980_ (.A_N(_07113_),
    .B(_07083_),
    .X(_07131_));
 sky130_fd_sc_hd__nor2_1 _13981_ (.A(_07130_),
    .B(_07131_),
    .Y(_07132_));
 sky130_fd_sc_hd__and2_1 _13982_ (.A(_07104_),
    .B(_07109_),
    .X(_07133_));
 sky130_fd_sc_hd__nor2_1 _13983_ (.A(_07102_),
    .B(_07110_),
    .Y(_07134_));
 sky130_fd_sc_hd__a21oi_2 _13984_ (.A1(_07086_),
    .A2(_07087_),
    .B1(_07100_),
    .Y(_07135_));
 sky130_fd_sc_hd__and2_1 _13985_ (.A(_07101_),
    .B(_07111_),
    .X(_07136_));
 sky130_fd_sc_hd__nand2_1 _13986_ (.A(_06700_),
    .B(_06738_),
    .Y(_07137_));
 sky130_fd_sc_hd__or2b_1 _13987_ (.A(_06880_),
    .B_N(_06694_),
    .X(_07138_));
 sky130_fd_sc_hd__nand2_1 _13988_ (.A(_06698_),
    .B(_06731_),
    .Y(_07139_));
 sky130_fd_sc_hd__xnor2_1 _13989_ (.A(_07138_),
    .B(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__xnor2_1 _13990_ (.A(_07137_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__xnor2_1 _13991_ (.A(_07090_),
    .B(_07141_),
    .Y(_07142_));
 sky130_fd_sc_hd__xnor2_1 _13992_ (.A(_06685_),
    .B(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__xnor2_1 _13993_ (.A(_07089_),
    .B(_07143_),
    .Y(_07144_));
 sky130_fd_sc_hd__nand2_1 _13994_ (.A(_07098_),
    .B(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__or2_1 _13995_ (.A(_07098_),
    .B(_07144_),
    .X(_07146_));
 sky130_fd_sc_hd__and2_1 _13996_ (.A(_07145_),
    .B(_07146_),
    .X(_07147_));
 sky130_fd_sc_hd__or4_1 _13997_ (.A(_06723_),
    .B(_06730_),
    .C(_06697_),
    .D(_07105_),
    .X(_07148_));
 sky130_fd_sc_hd__and2_1 _13998_ (.A(_07093_),
    .B(_07094_),
    .X(_07149_));
 sky130_fd_sc_hd__and2b_1 _13999_ (.A_N(_07095_),
    .B(_07096_),
    .X(_07150_));
 sky130_fd_sc_hd__or2_1 _14000_ (.A(_06720_),
    .B(_06702_),
    .X(_07151_));
 sky130_fd_sc_hd__or2_1 _14001_ (.A(_06713_),
    .B(_06696_),
    .X(_07152_));
 sky130_fd_sc_hd__xnor2_1 _14002_ (.A(_07151_),
    .B(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__or3_1 _14003_ (.A(_07105_),
    .B(_07107_),
    .C(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__o21ai_1 _14004_ (.A1(_07105_),
    .A2(_07107_),
    .B1(_07153_),
    .Y(_07155_));
 sky130_fd_sc_hd__and2_1 _14005_ (.A(_07154_),
    .B(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__o21ai_1 _14006_ (.A1(_07149_),
    .A2(_07150_),
    .B1(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__or3_1 _14007_ (.A(_07149_),
    .B(_07150_),
    .C(_07156_),
    .X(_07158_));
 sky130_fd_sc_hd__nand2_1 _14008_ (.A(_07157_),
    .B(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__xor2_1 _14009_ (.A(_07148_),
    .B(_07159_),
    .X(_07160_));
 sky130_fd_sc_hd__nand2_1 _14010_ (.A(_07147_),
    .B(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__or2_1 _14011_ (.A(_07147_),
    .B(_07160_),
    .X(_07162_));
 sky130_fd_sc_hd__o211ai_4 _14012_ (.A1(_07135_),
    .A2(_07136_),
    .B1(_07161_),
    .C1(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__a211o_1 _14013_ (.A1(_07161_),
    .A2(_07162_),
    .B1(_07135_),
    .C1(_07136_),
    .X(_07164_));
 sky130_fd_sc_hd__o211ai_2 _14014_ (.A1(_07133_),
    .A2(_07134_),
    .B1(_07163_),
    .C1(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__a211o_1 _14015_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07133_),
    .C1(_07134_),
    .X(_07166_));
 sky130_fd_sc_hd__and2_1 _14016_ (.A(_07165_),
    .B(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__xnor2_2 _14017_ (.A(_07132_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__nor2_1 _14018_ (.A(_07114_),
    .B(_07116_),
    .Y(_07169_));
 sky130_fd_sc_hd__or3_1 _14019_ (.A(_06862_),
    .B(_06907_),
    .C(_07117_),
    .X(_07170_));
 sky130_fd_sc_hd__and2b_1 _14020_ (.A_N(_07169_),
    .B(_07170_),
    .X(_07171_));
 sky130_fd_sc_hd__xnor2_1 _14021_ (.A(_07168_),
    .B(_07171_),
    .Y(_07172_));
 sky130_fd_sc_hd__xor2_2 _14022_ (.A(_07129_),
    .B(_07172_),
    .X(_07173_));
 sky130_fd_sc_hd__or2_2 _14023_ (.A(_07128_),
    .B(_07173_),
    .X(_07174_));
 sky130_fd_sc_hd__clkinv_2 _14024_ (.A(_07168_),
    .Y(_07175_));
 sky130_fd_sc_hd__a2bb2o_2 _14025_ (.A1_N(_07170_),
    .A2_N(_07175_),
    .B1(_07172_),
    .B2(_07129_),
    .X(_07176_));
 sky130_fd_sc_hd__nor2b_1 _14026_ (.A(_07132_),
    .B_N(_07167_),
    .Y(_07177_));
 sky130_fd_sc_hd__nand2_1 _14027_ (.A(_07145_),
    .B(_07161_),
    .Y(_07178_));
 sky130_fd_sc_hd__or3_1 _14028_ (.A(_06545_),
    .B(_06832_),
    .C(_07143_),
    .X(_07179_));
 sky130_fd_sc_hd__nand2_1 _14029_ (.A(_06694_),
    .B(_06731_),
    .Y(_07180_));
 sky130_fd_sc_hd__nand2_1 _14030_ (.A(_06880_),
    .B(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__o21a_1 _14031_ (.A1(_06942_),
    .A2(_07138_),
    .B1(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__xnor2_1 _14032_ (.A(_07179_),
    .B(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__nor2_1 _14033_ (.A(_07090_),
    .B(_07141_),
    .Y(_07184_));
 sky130_fd_sc_hd__nor2_1 _14034_ (.A(_06685_),
    .B(_07142_),
    .Y(_07185_));
 sky130_fd_sc_hd__or2_1 _14035_ (.A(_06713_),
    .B(_06702_),
    .X(_07186_));
 sky130_fd_sc_hd__or2_1 _14036_ (.A(_06614_),
    .B(_06696_),
    .X(_07187_));
 sky130_fd_sc_hd__nor2_1 _14037_ (.A(_07186_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__or3_1 _14038_ (.A(_07107_),
    .B(_07186_),
    .C(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__xnor2_1 _14039_ (.A(_07186_),
    .B(_07187_),
    .Y(_07190_));
 sky130_fd_sc_hd__o21ai_1 _14040_ (.A1(_07107_),
    .A2(_07186_),
    .B1(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__and2_1 _14041_ (.A(_07189_),
    .B(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__o21ai_1 _14042_ (.A1(_07184_),
    .A2(_07185_),
    .B1(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__or3_1 _14043_ (.A(_07184_),
    .B(_07185_),
    .C(_07192_),
    .X(_07194_));
 sky130_fd_sc_hd__nand2_1 _14044_ (.A(_07193_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__xor2_1 _14045_ (.A(_07154_),
    .B(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__and2_1 _14046_ (.A(_07183_),
    .B(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__nor2_1 _14047_ (.A(_07183_),
    .B(_07196_),
    .Y(_07198_));
 sky130_fd_sc_hd__or2_1 _14048_ (.A(_07197_),
    .B(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__xor2_1 _14049_ (.A(_07178_),
    .B(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__o21a_1 _14050_ (.A1(_07148_),
    .A2(_07159_),
    .B1(_07157_),
    .X(_07201_));
 sky130_fd_sc_hd__xnor2_1 _14051_ (.A(_07200_),
    .B(_07201_),
    .Y(_07202_));
 sky130_fd_sc_hd__a21oi_2 _14052_ (.A1(_07163_),
    .A2(_07165_),
    .B1(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__and3_1 _14053_ (.A(_07163_),
    .B(_07165_),
    .C(_07202_),
    .X(_07204_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_07203_),
    .B(_07204_),
    .Y(_07205_));
 sky130_fd_sc_hd__xor2_1 _14055_ (.A(_07177_),
    .B(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__and3_1 _14056_ (.A(_07169_),
    .B(_07168_),
    .C(_07206_),
    .X(_07207_));
 sky130_fd_sc_hd__a21oi_1 _14057_ (.A1(_07169_),
    .A2(_07168_),
    .B1(_07206_),
    .Y(_07208_));
 sky130_fd_sc_hd__nor2_2 _14058_ (.A(_07207_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__xor2_4 _14059_ (.A(_07176_),
    .B(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__nor2_2 _14060_ (.A(_07174_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__a21o_1 _14061_ (.A1(_07176_),
    .A2(_07209_),
    .B1(_07207_),
    .X(_07212_));
 sky130_fd_sc_hd__nand2_1 _14062_ (.A(_07177_),
    .B(_07205_),
    .Y(_07213_));
 sky130_fd_sc_hd__and2b_1 _14063_ (.A_N(_07199_),
    .B(_07178_),
    .X(_07214_));
 sky130_fd_sc_hd__nor2_1 _14064_ (.A(_07200_),
    .B(_07201_),
    .Y(_07215_));
 sky130_fd_sc_hd__and2b_1 _14065_ (.A_N(_07179_),
    .B(_07182_),
    .X(_07216_));
 sky130_fd_sc_hd__clkbuf_4 _14066_ (.A(_06880_),
    .X(_07217_));
 sky130_fd_sc_hd__a21o_1 _14067_ (.A1(_06880_),
    .A2(_07180_),
    .B1(_06685_),
    .X(_07218_));
 sky130_fd_sc_hd__o21ai_1 _14068_ (.A1(_07217_),
    .A2(_07180_),
    .B1(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__a22o_1 _14069_ (.A1(_06738_),
    .A2(_06694_),
    .B1(_06731_),
    .B2(_06558_),
    .X(_07220_));
 sky130_fd_sc_hd__or3_1 _14070_ (.A(_06484_),
    .B(_06725_),
    .C(_07180_),
    .X(_07221_));
 sky130_fd_sc_hd__and3_1 _14071_ (.A(_07219_),
    .B(_07220_),
    .C(_07221_),
    .X(_07222_));
 sky130_fd_sc_hd__a21oi_1 _14072_ (.A1(_07220_),
    .A2(_07221_),
    .B1(_07219_),
    .Y(_07223_));
 sky130_fd_sc_hd__or2_1 _14073_ (.A(_07222_),
    .B(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__o22a_1 _14074_ (.A1(_06614_),
    .A2(_06703_),
    .B1(_06696_),
    .B2(_06594_),
    .X(_07225_));
 sky130_fd_sc_hd__or4_1 _14075_ (.A(_06594_),
    .B(_06614_),
    .C(_06703_),
    .D(_06696_),
    .X(_07226_));
 sky130_fd_sc_hd__o21a_1 _14076_ (.A1(_06685_),
    .A2(_07182_),
    .B1(_07226_),
    .X(_07227_));
 sky130_fd_sc_hd__or3b_1 _14077_ (.A(_07188_),
    .B(_07225_),
    .C_N(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__xnor2_1 _14078_ (.A(_07189_),
    .B(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__or2_1 _14079_ (.A(_07224_),
    .B(_07229_),
    .X(_07230_));
 sky130_fd_sc_hd__nand2_1 _14080_ (.A(_07224_),
    .B(_07229_),
    .Y(_07231_));
 sky130_fd_sc_hd__and2_1 _14081_ (.A(_07230_),
    .B(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__o21a_1 _14082_ (.A1(_07216_),
    .A2(_07197_),
    .B1(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__or3_1 _14083_ (.A(_07216_),
    .B(_07197_),
    .C(_07232_),
    .X(_07234_));
 sky130_fd_sc_hd__and2b_1 _14084_ (.A_N(_07233_),
    .B(_07234_),
    .X(_07235_));
 sky130_fd_sc_hd__o21ai_1 _14085_ (.A1(_07154_),
    .A2(_07195_),
    .B1(_07193_),
    .Y(_07236_));
 sky130_fd_sc_hd__xor2_1 _14086_ (.A(_07235_),
    .B(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__o21a_1 _14087_ (.A1(_07214_),
    .A2(_07215_),
    .B1(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__nor3_1 _14088_ (.A(_07214_),
    .B(_07215_),
    .C(_07237_),
    .Y(_07239_));
 sky130_fd_sc_hd__nor2_1 _14089_ (.A(_07238_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__xor2_2 _14090_ (.A(_07203_),
    .B(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__xnor2_2 _14091_ (.A(_07213_),
    .B(_07241_),
    .Y(_07242_));
 sky130_fd_sc_hd__xnor2_4 _14092_ (.A(_07212_),
    .B(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__xnor2_4 _14093_ (.A(_07211_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__clkbuf_4 _14094_ (.A(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__nor2_1 _14095_ (.A(_06703_),
    .B(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__a21o_1 _14096_ (.A1(_07177_),
    .A2(_07205_),
    .B1(_07207_),
    .X(_07247_));
 sky130_fd_sc_hd__and3_1 _14097_ (.A(_06558_),
    .B(_06738_),
    .C(_07180_),
    .X(_07248_));
 sky130_fd_sc_hd__and3_1 _14098_ (.A(_06698_),
    .B(_07222_),
    .C(_07226_),
    .X(_07249_));
 sky130_fd_sc_hd__a21oi_1 _14099_ (.A1(_06698_),
    .A2(_07226_),
    .B1(_07222_),
    .Y(_07250_));
 sky130_fd_sc_hd__o21ba_1 _14100_ (.A1(_07249_),
    .A2(_07250_),
    .B1_N(_07188_),
    .X(_07251_));
 sky130_fd_sc_hd__xnor2_1 _14101_ (.A(_07248_),
    .B(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__o221a_1 _14102_ (.A1(_06685_),
    .A2(_07182_),
    .B1(_07189_),
    .B2(_07228_),
    .C1(_07230_),
    .X(_07253_));
 sky130_fd_sc_hd__xor2_1 _14103_ (.A(_07252_),
    .B(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__a211o_1 _14104_ (.A1(_07234_),
    .A2(_07236_),
    .B1(_07254_),
    .C1(_07233_),
    .X(_07255_));
 sky130_fd_sc_hd__o21ai_1 _14105_ (.A1(_07138_),
    .A2(_07139_),
    .B1(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__o2bb2a_1 _14106_ (.A1_N(_07203_),
    .A2_N(_07240_),
    .B1(_07256_),
    .B2(_07238_),
    .X(_07257_));
 sky130_fd_sc_hd__a21bo_1 _14107_ (.A1(_07238_),
    .A2(_07256_),
    .B1_N(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__and3_1 _14108_ (.A(_07176_),
    .B(_07209_),
    .C(_07242_),
    .X(_07259_));
 sky130_fd_sc_hd__a211oi_2 _14109_ (.A1(_07241_),
    .A2(_07247_),
    .B1(_07258_),
    .C1(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__a21oi_4 _14110_ (.A1(_07211_),
    .A2(_07243_),
    .B1(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__buf_2 _14111_ (.A(_07261_),
    .X(_07262_));
 sky130_fd_sc_hd__and3_1 _14112_ (.A(_06701_),
    .B(_06727_),
    .C(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__nand2_1 _14113_ (.A(_06731_),
    .B(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__clkbuf_4 _14114_ (.A(_07262_),
    .X(_07265_));
 sky130_fd_sc_hd__nand2_2 _14115_ (.A(_06738_),
    .B(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__nand2_1 _14116_ (.A(_06731_),
    .B(_07262_),
    .Y(_07267_));
 sky130_fd_sc_hd__xnor2_2 _14117_ (.A(_07267_),
    .B(_07263_),
    .Y(_07268_));
 sky130_fd_sc_hd__or2b_1 _14118_ (.A(_07266_),
    .B_N(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__or2_2 _14119_ (.A(_06545_),
    .B(_07261_),
    .X(_07270_));
 sky130_fd_sc_hd__o21a_1 _14120_ (.A1(_07217_),
    .A2(_07270_),
    .B1(_07267_),
    .X(_07271_));
 sky130_fd_sc_hd__nor2_2 _14121_ (.A(_07266_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__a21o_1 _14122_ (.A1(_07264_),
    .A2(_07269_),
    .B1(_07272_),
    .X(_07273_));
 sky130_fd_sc_hd__o211a_1 _14123_ (.A1(_06697_),
    .A2(_07246_),
    .B1(_07273_),
    .C1(_07265_),
    .X(_07274_));
 sky130_fd_sc_hd__o21a_1 _14124_ (.A1(_06942_),
    .A2(_07270_),
    .B1(_07266_),
    .X(_07275_));
 sky130_fd_sc_hd__nor2_1 _14125_ (.A(_07272_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__a21bo_1 _14126_ (.A1(_07274_),
    .A2(_07276_),
    .B1_N(_07273_),
    .X(_07277_));
 sky130_fd_sc_hd__buf_2 _14127_ (.A(_06725_),
    .X(_07278_));
 sky130_fd_sc_hd__mux2_1 _14128_ (.A0(_07278_),
    .A1(_07272_),
    .S(_07265_),
    .X(_07279_));
 sky130_fd_sc_hd__or2_1 _14129_ (.A(_07277_),
    .B(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__nand2_1 _14130_ (.A(_07266_),
    .B(_07271_),
    .Y(_07281_));
 sky130_fd_sc_hd__a21o_1 _14131_ (.A1(_07273_),
    .A2(_07281_),
    .B1(_06545_),
    .X(_07282_));
 sky130_fd_sc_hd__xnor2_4 _14132_ (.A(_07174_),
    .B(_07210_),
    .Y(_07283_));
 sky130_fd_sc_hd__clkbuf_4 _14133_ (.A(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__nor2_1 _14134_ (.A(_06697_),
    .B(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__inv_2 _14135_ (.A(_06697_),
    .Y(_07286_));
 sky130_fd_sc_hd__nand2_1 _14136_ (.A(_07286_),
    .B(_07265_),
    .Y(_07287_));
 sky130_fd_sc_hd__or2_1 _14137_ (.A(_07285_),
    .B(_07287_),
    .X(_07288_));
 sky130_fd_sc_hd__a21o_1 _14138_ (.A1(_07246_),
    .A2(_07288_),
    .B1(_07249_),
    .X(_07289_));
 sky130_fd_sc_hd__nand2_1 _14139_ (.A(_07282_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__a21oi_2 _14140_ (.A1(_07274_),
    .A2(_07276_),
    .B1(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__xor2_2 _14141_ (.A(_07280_),
    .B(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__nor2_1 _14142_ (.A(_07274_),
    .B(_07276_),
    .Y(_07293_));
 sky130_fd_sc_hd__o22a_1 _14143_ (.A1(_07246_),
    .A2(_07287_),
    .B1(_07291_),
    .B2(_07293_),
    .X(_07294_));
 sky130_fd_sc_hd__xnor2_2 _14144_ (.A(_07128_),
    .B(_07173_),
    .Y(_07295_));
 sky130_fd_sc_hd__clkbuf_4 _14145_ (.A(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__nor2_1 _14146_ (.A(_06703_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__nand2_1 _14147_ (.A(_07297_),
    .B(_07285_),
    .Y(_07298_));
 sky130_fd_sc_hd__or2_1 _14148_ (.A(_07121_),
    .B(_07127_),
    .X(_07299_));
 sky130_fd_sc_hd__nand2_2 _14149_ (.A(_07128_),
    .B(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__clkbuf_4 _14150_ (.A(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__nor2_1 _14151_ (.A(_06697_),
    .B(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__and3_1 _14152_ (.A(_07297_),
    .B(_07298_),
    .C(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__and3_1 _14153_ (.A(_06802_),
    .B(_06775_),
    .C(_07265_),
    .X(_07304_));
 sky130_fd_sc_hd__nor2_1 _14154_ (.A(_07278_),
    .B(_07245_),
    .Y(_07305_));
 sky130_fd_sc_hd__xor2_1 _14155_ (.A(_07268_),
    .B(_07305_),
    .X(_07306_));
 sky130_fd_sc_hd__nand2_1 _14156_ (.A(_07304_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__xnor2_1 _14157_ (.A(_07304_),
    .B(_07306_),
    .Y(_07308_));
 sky130_fd_sc_hd__nor2_1 _14158_ (.A(_07278_),
    .B(_07284_),
    .Y(_07309_));
 sky130_fd_sc_hd__or2_1 _14159_ (.A(_06942_),
    .B(_07245_),
    .X(_07310_));
 sky130_fd_sc_hd__xnor2_1 _14160_ (.A(_07263_),
    .B(_07310_),
    .Y(_07311_));
 sky130_fd_sc_hd__nand2_1 _14161_ (.A(_07309_),
    .B(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__o31a_1 _14162_ (.A1(_07217_),
    .A2(_07267_),
    .A3(_07245_),
    .B1(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__or2_1 _14163_ (.A(_07308_),
    .B(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__or2_1 _14164_ (.A(_06697_),
    .B(_07245_),
    .X(_07315_));
 sky130_fd_sc_hd__or2_1 _14165_ (.A(_06697_),
    .B(_07296_),
    .X(_07316_));
 sky130_fd_sc_hd__or3b_1 _14166_ (.A(_06703_),
    .B(_07284_),
    .C_N(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__xnor2_1 _14167_ (.A(_07315_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__a21oi_1 _14168_ (.A1(_07307_),
    .A2(_07314_),
    .B1(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__and3_1 _14169_ (.A(_07307_),
    .B(_07314_),
    .C(_07318_),
    .X(_07320_));
 sky130_fd_sc_hd__nor2_1 _14170_ (.A(_07319_),
    .B(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__a21o_1 _14171_ (.A1(_07303_),
    .A2(_07321_),
    .B1(_07319_),
    .X(_07322_));
 sky130_fd_sc_hd__or2_1 _14172_ (.A(_07282_),
    .B(_07289_),
    .X(_07323_));
 sky130_fd_sc_hd__nand2_1 _14173_ (.A(_07290_),
    .B(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__xor2_1 _14174_ (.A(_07303_),
    .B(_07321_),
    .X(_07325_));
 sky130_fd_sc_hd__clkbuf_4 _14175_ (.A(_07036_),
    .X(_07326_));
 sky130_fd_sc_hd__nand2_1 _14176_ (.A(_06775_),
    .B(_07265_),
    .Y(_07327_));
 sky130_fd_sc_hd__o21ai_2 _14177_ (.A1(_07326_),
    .A2(_07265_),
    .B1(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__xor2_1 _14178_ (.A(_07308_),
    .B(_07313_),
    .X(_07329_));
 sky130_fd_sc_hd__nand2_1 _14179_ (.A(_07328_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__clkbuf_4 _14180_ (.A(_06832_),
    .X(_07331_));
 sky130_fd_sc_hd__nand2_1 _14181_ (.A(_07268_),
    .B(_07305_),
    .Y(_07332_));
 sky130_fd_sc_hd__xor2_1 _14182_ (.A(_07266_),
    .B(_07268_),
    .X(_07333_));
 sky130_fd_sc_hd__a31o_1 _14183_ (.A1(_07264_),
    .A2(_07332_),
    .A3(_07333_),
    .B1(_07249_),
    .X(_07334_));
 sky130_fd_sc_hd__o21a_1 _14184_ (.A1(_07331_),
    .A2(_07265_),
    .B1(_07334_),
    .X(_07335_));
 sky130_fd_sc_hd__nor2_1 _14185_ (.A(_07330_),
    .B(_07335_),
    .Y(_07336_));
 sky130_fd_sc_hd__and2_1 _14186_ (.A(_07330_),
    .B(_07335_),
    .X(_07337_));
 sky130_fd_sc_hd__nor2_1 _14187_ (.A(_07336_),
    .B(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__a21oi_1 _14188_ (.A1(_07325_),
    .A2(_07338_),
    .B1(_07336_),
    .Y(_07339_));
 sky130_fd_sc_hd__xor2_1 _14189_ (.A(_07324_),
    .B(_07339_),
    .X(_07340_));
 sky130_fd_sc_hd__nor2_1 _14190_ (.A(_07324_),
    .B(_07339_),
    .Y(_07341_));
 sky130_fd_sc_hd__a21oi_1 _14191_ (.A1(_07322_),
    .A2(_07340_),
    .B1(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__nor2_1 _14192_ (.A(_07294_),
    .B(_07342_),
    .Y(_07343_));
 sky130_fd_sc_hd__and2b_1 _14193_ (.A_N(_07292_),
    .B(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__mux2_1 _14194_ (.A0(_07278_),
    .A1(_07286_),
    .S(_07265_),
    .X(_07345_));
 sky130_fd_sc_hd__nor2_1 _14195_ (.A(_07272_),
    .B(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__a2bb2o_1 _14196_ (.A1_N(_07290_),
    .A2_N(_07280_),
    .B1(_07346_),
    .B2(_07277_),
    .X(_07347_));
 sky130_fd_sc_hd__o21ba_1 _14197_ (.A1(_07277_),
    .A2(_07346_),
    .B1_N(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__xor2_1 _14198_ (.A(_07344_),
    .B(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__inv_2 _14199_ (.A(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__xnor2_1 _14200_ (.A(_07322_),
    .B(_07340_),
    .Y(_07351_));
 sky130_fd_sc_hd__nor2_1 _14201_ (.A(_06703_),
    .B(_07301_),
    .Y(_07352_));
 sky130_fd_sc_hd__and2_1 _14202_ (.A(_07122_),
    .B(_07126_),
    .X(_07353_));
 sky130_fd_sc_hd__or2_1 _14203_ (.A(_07127_),
    .B(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__clkbuf_4 _14204_ (.A(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__nor2_1 _14205_ (.A(_06697_),
    .B(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__and3_1 _14206_ (.A(_07316_),
    .B(_07352_),
    .C(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__or2_1 _14207_ (.A(_07297_),
    .B(_07285_),
    .X(_07358_));
 sky130_fd_sc_hd__a22o_1 _14208_ (.A1(_07297_),
    .A2(_07302_),
    .B1(_07358_),
    .B2(_07298_),
    .X(_07359_));
 sky130_fd_sc_hd__or2b_1 _14209_ (.A(_07303_),
    .B_N(_07359_),
    .X(_07360_));
 sky130_fd_sc_hd__or2_1 _14210_ (.A(_07278_),
    .B(_07296_),
    .X(_07361_));
 sky130_fd_sc_hd__o22a_1 _14211_ (.A1(_06942_),
    .A2(_07284_),
    .B1(_07245_),
    .B2(_07217_),
    .X(_07362_));
 sky130_fd_sc_hd__nor2_1 _14212_ (.A(_07361_),
    .B(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__and2_1 _14213_ (.A(_06716_),
    .B(_07261_),
    .X(_07364_));
 sky130_fd_sc_hd__clkbuf_2 _14214_ (.A(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__nand2_1 _14215_ (.A(_06802_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__nand2_1 _14216_ (.A(_06802_),
    .B(_07261_),
    .Y(_07367_));
 sky130_fd_sc_hd__xor2_2 _14217_ (.A(_07367_),
    .B(_07365_),
    .X(_07368_));
 sky130_fd_sc_hd__or2_1 _14218_ (.A(_07327_),
    .B(_07368_),
    .X(_07369_));
 sky130_fd_sc_hd__xnor2_1 _14219_ (.A(_07309_),
    .B(_07311_),
    .Y(_07370_));
 sky130_fd_sc_hd__a21o_1 _14220_ (.A1(_07366_),
    .A2(_07369_),
    .B1(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__nand3_1 _14221_ (.A(_07366_),
    .B(_07369_),
    .C(_07370_),
    .Y(_07372_));
 sky130_fd_sc_hd__and2_1 _14222_ (.A(_07371_),
    .B(_07372_),
    .X(_07373_));
 sky130_fd_sc_hd__a21bo_1 _14223_ (.A1(_07363_),
    .A2(_07373_),
    .B1_N(_07371_),
    .X(_07374_));
 sky130_fd_sc_hd__xnor2_1 _14224_ (.A(_07360_),
    .B(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__or2b_1 _14225_ (.A(_07360_),
    .B_N(_07374_),
    .X(_07376_));
 sky130_fd_sc_hd__a21bo_1 _14226_ (.A1(_07357_),
    .A2(_07375_),
    .B1_N(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__xnor2_1 _14227_ (.A(_07325_),
    .B(_07338_),
    .Y(_07378_));
 sky130_fd_sc_hd__xor2_1 _14228_ (.A(_07357_),
    .B(_07375_),
    .X(_07379_));
 sky130_fd_sc_hd__o211a_1 _14229_ (.A1(_07066_),
    .A2(_07270_),
    .B1(_07327_),
    .C1(_07367_),
    .X(_07380_));
 sky130_fd_sc_hd__nor2_1 _14230_ (.A(_07304_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__xor2_2 _14231_ (.A(_07363_),
    .B(_07373_),
    .X(_07382_));
 sky130_fd_sc_hd__xor2_1 _14232_ (.A(_07328_),
    .B(_07329_),
    .X(_07383_));
 sky130_fd_sc_hd__and3_1 _14233_ (.A(_07381_),
    .B(_07382_),
    .C(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__a21oi_1 _14234_ (.A1(_07381_),
    .A2(_07382_),
    .B1(_07383_),
    .Y(_07385_));
 sky130_fd_sc_hd__nor2_1 _14235_ (.A(_07384_),
    .B(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__a21oi_1 _14236_ (.A1(_07379_),
    .A2(_07386_),
    .B1(_07384_),
    .Y(_07387_));
 sky130_fd_sc_hd__nor2_1 _14237_ (.A(_07378_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__and2_1 _14238_ (.A(_07378_),
    .B(_07387_),
    .X(_07389_));
 sky130_fd_sc_hd__nor2_1 _14239_ (.A(_07388_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__a21oi_1 _14240_ (.A1(_07377_),
    .A2(_07390_),
    .B1(_07388_),
    .Y(_07391_));
 sky130_fd_sc_hd__nor2_1 _14241_ (.A(_07351_),
    .B(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__and2_1 _14242_ (.A(_07294_),
    .B(_07342_),
    .X(_07393_));
 sky130_fd_sc_hd__nor2_1 _14243_ (.A(_07343_),
    .B(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__a21oi_1 _14244_ (.A1(_07392_),
    .A2(_07394_),
    .B1(_07343_),
    .Y(_07395_));
 sky130_fd_sc_hd__xor2_1 _14245_ (.A(_07292_),
    .B(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__inv_2 _14246_ (.A(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__nand2_1 _14247_ (.A(_07392_),
    .B(_07394_),
    .Y(_07398_));
 sky130_fd_sc_hd__or2_1 _14248_ (.A(_07392_),
    .B(_07394_),
    .X(_07399_));
 sky130_fd_sc_hd__and2_1 _14249_ (.A(_07398_),
    .B(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__xnor2_1 _14250_ (.A(_07377_),
    .B(_07390_),
    .Y(_07401_));
 sky130_fd_sc_hd__and2_1 _14251_ (.A(_07123_),
    .B(_07125_),
    .X(_07402_));
 sky130_fd_sc_hd__nor2_1 _14252_ (.A(_07126_),
    .B(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__buf_2 _14253_ (.A(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__nor2_1 _14254_ (.A(_06703_),
    .B(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__nand2_1 _14255_ (.A(_07356_),
    .B(_07405_),
    .Y(_07406_));
 sky130_fd_sc_hd__nand2_1 _14256_ (.A(_07352_),
    .B(_07356_),
    .Y(_07407_));
 sky130_fd_sc_hd__nor2_1 _14257_ (.A(_06703_),
    .B(_07355_),
    .Y(_07408_));
 sky130_fd_sc_hd__or2_1 _14258_ (.A(_07302_),
    .B(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__a21oi_1 _14259_ (.A1(_07407_),
    .A2(_07409_),
    .B1(_06545_),
    .Y(_07410_));
 sky130_fd_sc_hd__nor2_1 _14260_ (.A(_07406_),
    .B(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__xnor2_1 _14261_ (.A(_07316_),
    .B(_07352_),
    .Y(_07412_));
 sky130_fd_sc_hd__a21oi_1 _14262_ (.A1(_07302_),
    .A2(_07408_),
    .B1(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__or2_1 _14263_ (.A(_07357_),
    .B(_07413_),
    .X(_07414_));
 sky130_fd_sc_hd__o31a_1 _14264_ (.A1(_07331_),
    .A2(_07245_),
    .A3(_07368_),
    .B1(_07366_),
    .X(_07415_));
 sky130_fd_sc_hd__and2_1 _14265_ (.A(_07361_),
    .B(_07362_),
    .X(_07416_));
 sky130_fd_sc_hd__or2_1 _14266_ (.A(_07363_),
    .B(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__xnor2_1 _14267_ (.A(_07415_),
    .B(_07417_),
    .Y(_07418_));
 sky130_fd_sc_hd__nor2_1 _14268_ (.A(_06942_),
    .B(_07295_),
    .Y(_07419_));
 sky130_fd_sc_hd__nor2_1 _14269_ (.A(_07217_),
    .B(_07283_),
    .Y(_07420_));
 sky130_fd_sc_hd__xor2_1 _14270_ (.A(_07419_),
    .B(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__or3b_1 _14271_ (.A(_07278_),
    .B(_07301_),
    .C_N(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__a21boi_1 _14272_ (.A1(_07419_),
    .A2(_07420_),
    .B1_N(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__or2_1 _14273_ (.A(_07415_),
    .B(_07417_),
    .X(_07424_));
 sky130_fd_sc_hd__o21a_1 _14274_ (.A1(_07418_),
    .A2(_07423_),
    .B1(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__nor2_1 _14275_ (.A(_07414_),
    .B(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__and2_1 _14276_ (.A(_07414_),
    .B(_07425_),
    .X(_07427_));
 sky130_fd_sc_hd__nor2_1 _14277_ (.A(_07426_),
    .B(_07427_),
    .Y(_07428_));
 sky130_fd_sc_hd__a21o_1 _14278_ (.A1(_07411_),
    .A2(_07428_),
    .B1(_07426_),
    .X(_07429_));
 sky130_fd_sc_hd__xnor2_1 _14279_ (.A(_07379_),
    .B(_07386_),
    .Y(_07430_));
 sky130_fd_sc_hd__xnor2_1 _14280_ (.A(_07411_),
    .B(_07428_),
    .Y(_07431_));
 sky130_fd_sc_hd__xnor2_1 _14281_ (.A(_07381_),
    .B(_07382_),
    .Y(_07432_));
 sky130_fd_sc_hd__or2_1 _14282_ (.A(_06799_),
    .B(_07265_),
    .X(_07433_));
 sky130_fd_sc_hd__nand2_1 _14283_ (.A(_07327_),
    .B(_07368_),
    .Y(_07434_));
 sky130_fd_sc_hd__nand2_1 _14284_ (.A(_07369_),
    .B(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__nor2_1 _14285_ (.A(_06832_),
    .B(_07245_),
    .Y(_07436_));
 sky130_fd_sc_hd__xnor2_2 _14286_ (.A(_07368_),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__and3_1 _14287_ (.A(_06761_),
    .B(_06768_),
    .C(_07262_),
    .X(_07438_));
 sky130_fd_sc_hd__nand2_1 _14288_ (.A(_06768_),
    .B(_07262_),
    .Y(_07439_));
 sky130_fd_sc_hd__o21a_1 _14289_ (.A1(_07044_),
    .A2(_07270_),
    .B1(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__nor2_1 _14290_ (.A(_07438_),
    .B(_07440_),
    .Y(_07441_));
 sky130_fd_sc_hd__a21oi_1 _14291_ (.A1(_07437_),
    .A2(_07441_),
    .B1(_07438_),
    .Y(_07442_));
 sky130_fd_sc_hd__a31o_1 _14292_ (.A1(_06558_),
    .A2(_07433_),
    .A3(_07435_),
    .B1(_07442_),
    .X(_07443_));
 sky130_fd_sc_hd__xor2_1 _14293_ (.A(_07418_),
    .B(_07423_),
    .X(_07444_));
 sky130_fd_sc_hd__nand4_1 _14294_ (.A(_06558_),
    .B(_07433_),
    .C(_07435_),
    .D(_07442_),
    .Y(_07445_));
 sky130_fd_sc_hd__and2_1 _14295_ (.A(_07443_),
    .B(_07445_),
    .X(_07446_));
 sky130_fd_sc_hd__nand2_1 _14296_ (.A(_07444_),
    .B(_07446_),
    .Y(_07447_));
 sky130_fd_sc_hd__and3_1 _14297_ (.A(_07432_),
    .B(_07443_),
    .C(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__a21o_1 _14298_ (.A1(_07443_),
    .A2(_07447_),
    .B1(_07432_),
    .X(_07449_));
 sky130_fd_sc_hd__o21a_1 _14299_ (.A1(_07431_),
    .A2(_07448_),
    .B1(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__nor2_1 _14300_ (.A(_07430_),
    .B(_07450_),
    .Y(_07451_));
 sky130_fd_sc_hd__and2_1 _14301_ (.A(_07430_),
    .B(_07450_),
    .X(_07452_));
 sky130_fd_sc_hd__nor2_1 _14302_ (.A(_07451_),
    .B(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__a21oi_1 _14303_ (.A1(_07429_),
    .A2(_07453_),
    .B1(_07451_),
    .Y(_07454_));
 sky130_fd_sc_hd__nor2_1 _14304_ (.A(_07401_),
    .B(_07454_),
    .Y(_07455_));
 sky130_fd_sc_hd__xor2_1 _14305_ (.A(_07351_),
    .B(_07391_),
    .X(_07456_));
 sky130_fd_sc_hd__and2_1 _14306_ (.A(_07455_),
    .B(_07456_),
    .X(_07457_));
 sky130_fd_sc_hd__xor2_1 _14307_ (.A(_07400_),
    .B(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__inv_2 _14308_ (.A(_07458_),
    .Y(_07459_));
 sky130_fd_sc_hd__nor2_1 _14309_ (.A(_07455_),
    .B(_07456_),
    .Y(_07460_));
 sky130_fd_sc_hd__nor2_1 _14310_ (.A(_07457_),
    .B(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__xnor2_2 _14311_ (.A(_07429_),
    .B(_07453_),
    .Y(_07462_));
 sky130_fd_sc_hd__nand3_1 _14312_ (.A(_07432_),
    .B(_07443_),
    .C(_07447_),
    .Y(_07463_));
 sky130_fd_sc_hd__nand2_1 _14313_ (.A(_07449_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__xnor2_1 _14314_ (.A(_07431_),
    .B(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__buf_2 _14315_ (.A(_07125_),
    .X(_07466_));
 sky130_fd_sc_hd__nor2_1 _14316_ (.A(_06697_),
    .B(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__and2_1 _14317_ (.A(_07405_),
    .B(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__nand2_1 _14318_ (.A(_07406_),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__and2_1 _14319_ (.A(_07406_),
    .B(_07410_),
    .X(_07470_));
 sky130_fd_sc_hd__or2_1 _14320_ (.A(_07411_),
    .B(_07470_),
    .X(_07471_));
 sky130_fd_sc_hd__nor2_1 _14321_ (.A(_07326_),
    .B(_07244_),
    .Y(_07472_));
 sky130_fd_sc_hd__xor2_1 _14322_ (.A(_07365_),
    .B(_07472_),
    .X(_07473_));
 sky130_fd_sc_hd__nor2_1 _14323_ (.A(_07331_),
    .B(_07284_),
    .Y(_07474_));
 sky130_fd_sc_hd__nand2_1 _14324_ (.A(_07365_),
    .B(_07472_),
    .Y(_07475_));
 sky130_fd_sc_hd__a21boi_2 _14325_ (.A1(_07473_),
    .A2(_07474_),
    .B1_N(_07475_),
    .Y(_07476_));
 sky130_fd_sc_hd__o21bai_1 _14326_ (.A1(_07278_),
    .A2(_07301_),
    .B1_N(_07421_),
    .Y(_07477_));
 sky130_fd_sc_hd__nand2_1 _14327_ (.A(_07422_),
    .B(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__xnor2_2 _14328_ (.A(_07476_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__nor2_1 _14329_ (.A(_07217_),
    .B(_07295_),
    .Y(_07480_));
 sky130_fd_sc_hd__nor2_2 _14330_ (.A(_06942_),
    .B(_07300_),
    .Y(_07481_));
 sky130_fd_sc_hd__or2_1 _14331_ (.A(_07278_),
    .B(_07354_),
    .X(_07482_));
 sky130_fd_sc_hd__xnor2_1 _14332_ (.A(_07480_),
    .B(_07481_),
    .Y(_07483_));
 sky130_fd_sc_hd__nor2_1 _14333_ (.A(_07482_),
    .B(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__a21oi_2 _14334_ (.A1(_07480_),
    .A2(_07481_),
    .B1(_07484_),
    .Y(_07485_));
 sky130_fd_sc_hd__or2_1 _14335_ (.A(_07476_),
    .B(_07478_),
    .X(_07486_));
 sky130_fd_sc_hd__o21a_1 _14336_ (.A1(_07479_),
    .A2(_07485_),
    .B1(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__nor2_1 _14337_ (.A(_07471_),
    .B(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__and2_1 _14338_ (.A(_07471_),
    .B(_07487_),
    .X(_07489_));
 sky130_fd_sc_hd__nor2_1 _14339_ (.A(_07488_),
    .B(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__xnor2_1 _14340_ (.A(_07469_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__xnor2_1 _14341_ (.A(_07444_),
    .B(_07446_),
    .Y(_07492_));
 sky130_fd_sc_hd__xor2_2 _14342_ (.A(_07479_),
    .B(_07485_),
    .X(_07493_));
 sky130_fd_sc_hd__xor2_2 _14343_ (.A(_07437_),
    .B(_07441_),
    .X(_07494_));
 sky130_fd_sc_hd__nand2_1 _14344_ (.A(_06761_),
    .B(_07262_),
    .Y(_07495_));
 sky130_fd_sc_hd__o211a_1 _14345_ (.A1(_07051_),
    .A2(_07270_),
    .B1(_07439_),
    .C1(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__xnor2_1 _14346_ (.A(_07473_),
    .B(_07474_),
    .Y(_07497_));
 sky130_fd_sc_hd__nand2_1 _14347_ (.A(_07042_),
    .B(_07262_),
    .Y(_07498_));
 sky130_fd_sc_hd__or3b_1 _14348_ (.A(_06632_),
    .B(_06799_),
    .C_N(_07261_),
    .X(_07499_));
 sky130_fd_sc_hd__a21oi_1 _14349_ (.A1(_07498_),
    .A2(_07499_),
    .B1(_07438_),
    .Y(_07500_));
 sky130_fd_sc_hd__o21ba_1 _14350_ (.A1(_07496_),
    .A2(_07497_),
    .B1_N(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__xnor2_2 _14351_ (.A(_07494_),
    .B(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__or2b_1 _14352_ (.A(_07501_),
    .B_N(_07494_),
    .X(_07503_));
 sky130_fd_sc_hd__a21boi_1 _14353_ (.A1(_07493_),
    .A2(_07502_),
    .B1_N(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__xor2_1 _14354_ (.A(_07492_),
    .B(_07504_),
    .X(_07505_));
 sky130_fd_sc_hd__nor2_1 _14355_ (.A(_07492_),
    .B(_07504_),
    .Y(_07506_));
 sky130_fd_sc_hd__a21oi_1 _14356_ (.A1(_07491_),
    .A2(_07505_),
    .B1(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__xnor2_1 _14357_ (.A(_07465_),
    .B(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__a31o_1 _14358_ (.A1(_07406_),
    .A2(_07468_),
    .A3(_07490_),
    .B1(_07488_),
    .X(_07509_));
 sky130_fd_sc_hd__or2b_1 _14359_ (.A(_07508_),
    .B_N(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__o21a_1 _14360_ (.A1(_07465_),
    .A2(_07507_),
    .B1(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__nor2_1 _14361_ (.A(_07462_),
    .B(_07511_),
    .Y(_07512_));
 sky130_fd_sc_hd__and2_1 _14362_ (.A(_07401_),
    .B(_07454_),
    .X(_07513_));
 sky130_fd_sc_hd__nor2_1 _14363_ (.A(_07455_),
    .B(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__and3_1 _14364_ (.A(_07461_),
    .B(_07512_),
    .C(_07514_),
    .X(_07515_));
 sky130_fd_sc_hd__a21oi_1 _14365_ (.A1(_07512_),
    .A2(_07514_),
    .B1(_07461_),
    .Y(_07516_));
 sky130_fd_sc_hd__nor2_1 _14366_ (.A(_07515_),
    .B(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__inv_2 _14367_ (.A(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__xor2_1 _14368_ (.A(_07509_),
    .B(_07508_),
    .X(_07519_));
 sky130_fd_sc_hd__or2_1 _14369_ (.A(_07066_),
    .B(_07283_),
    .X(_07520_));
 sky130_fd_sc_hd__or3_1 _14370_ (.A(_07326_),
    .B(_07244_),
    .C(_07520_),
    .X(_07521_));
 sky130_fd_sc_hd__nor2_1 _14371_ (.A(_07326_),
    .B(_07283_),
    .Y(_07522_));
 sky130_fd_sc_hd__o21ba_1 _14372_ (.A1(_07066_),
    .A2(_07244_),
    .B1_N(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__or4b_1 _14373_ (.A(_06832_),
    .B(_07523_),
    .C(_07296_),
    .D_N(_07521_),
    .X(_07524_));
 sky130_fd_sc_hd__xnor2_1 _14374_ (.A(_07482_),
    .B(_07483_),
    .Y(_07525_));
 sky130_fd_sc_hd__a21oi_1 _14375_ (.A1(_07521_),
    .A2(_07524_),
    .B1(_07525_),
    .Y(_07526_));
 sky130_fd_sc_hd__and3_1 _14376_ (.A(_07521_),
    .B(_07524_),
    .C(_07525_),
    .X(_07527_));
 sky130_fd_sc_hd__or2_1 _14377_ (.A(_07526_),
    .B(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__or2_1 _14378_ (.A(_07217_),
    .B(_07354_),
    .X(_07529_));
 sky130_fd_sc_hd__inv_2 _14379_ (.A(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__or2_1 _14380_ (.A(_07278_),
    .B(_07403_),
    .X(_07531_));
 sky130_fd_sc_hd__o22a_1 _14381_ (.A1(_07217_),
    .A2(_07301_),
    .B1(_07355_),
    .B2(_06942_),
    .X(_07532_));
 sky130_fd_sc_hd__a21o_1 _14382_ (.A1(_07481_),
    .A2(_07530_),
    .B1(_07532_),
    .X(_07533_));
 sky130_fd_sc_hd__o2bb2a_1 _14383_ (.A1_N(_07481_),
    .A2_N(_07530_),
    .B1(_07531_),
    .B2(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__nor2_1 _14384_ (.A(_07528_),
    .B(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__or2_1 _14385_ (.A(_07406_),
    .B(_07468_),
    .X(_07536_));
 sky130_fd_sc_hd__o211a_1 _14386_ (.A1(_07356_),
    .A2(_07405_),
    .B1(_07469_),
    .C1(_07536_),
    .X(_07537_));
 sky130_fd_sc_hd__o21a_1 _14387_ (.A1(_07526_),
    .A2(_07535_),
    .B1(_07537_),
    .X(_07538_));
 sky130_fd_sc_hd__xnor2_1 _14388_ (.A(_07491_),
    .B(_07505_),
    .Y(_07539_));
 sky130_fd_sc_hd__nor3_1 _14389_ (.A(_07526_),
    .B(_07535_),
    .C(_07537_),
    .Y(_07540_));
 sky130_fd_sc_hd__nor2_1 _14390_ (.A(_07538_),
    .B(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__xnor2_2 _14391_ (.A(_07493_),
    .B(_07502_),
    .Y(_07542_));
 sky130_fd_sc_hd__xor2_1 _14392_ (.A(_07528_),
    .B(_07534_),
    .X(_07543_));
 sky130_fd_sc_hd__or2_1 _14393_ (.A(_07496_),
    .B(_07500_),
    .X(_07544_));
 sky130_fd_sc_hd__xnor2_1 _14394_ (.A(_07497_),
    .B(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__nor2_1 _14395_ (.A(_07066_),
    .B(_07284_),
    .Y(_07546_));
 sky130_fd_sc_hd__a21oi_1 _14396_ (.A1(_07472_),
    .A2(_07546_),
    .B1(_07523_),
    .Y(_07547_));
 sky130_fd_sc_hd__nor2_1 _14397_ (.A(_07331_),
    .B(_07296_),
    .Y(_07548_));
 sky130_fd_sc_hd__xnor2_1 _14398_ (.A(_07547_),
    .B(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__o21a_1 _14399_ (.A1(_06745_),
    .A2(_06768_),
    .B1(_07262_),
    .X(_07550_));
 sky130_fd_sc_hd__nand2_1 _14400_ (.A(_07499_),
    .B(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__and2_1 _14401_ (.A(_06745_),
    .B(_07262_),
    .X(_07552_));
 sky130_fd_sc_hd__nor2_1 _14402_ (.A(_06799_),
    .B(_07245_),
    .Y(_07553_));
 sky130_fd_sc_hd__a21bo_1 _14403_ (.A1(_07552_),
    .A2(_07553_),
    .B1_N(_07498_),
    .X(_07554_));
 sky130_fd_sc_hd__xor2_1 _14404_ (.A(_07551_),
    .B(_07554_),
    .X(_07555_));
 sky130_fd_sc_hd__or2b_1 _14405_ (.A(_07551_),
    .B_N(_07554_),
    .X(_07556_));
 sky130_fd_sc_hd__o21ai_1 _14406_ (.A1(_07549_),
    .A2(_07555_),
    .B1(_07556_),
    .Y(_07557_));
 sky130_fd_sc_hd__xnor2_1 _14407_ (.A(_07545_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__or2b_1 _14408_ (.A(_07545_),
    .B_N(_07557_),
    .X(_07559_));
 sky130_fd_sc_hd__a21boi_2 _14409_ (.A1(_07543_),
    .A2(_07558_),
    .B1_N(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__xor2_2 _14410_ (.A(_07542_),
    .B(_07560_),
    .X(_07561_));
 sky130_fd_sc_hd__nor2_1 _14411_ (.A(_07542_),
    .B(_07560_),
    .Y(_07562_));
 sky130_fd_sc_hd__a21oi_1 _14412_ (.A1(_07541_),
    .A2(_07561_),
    .B1(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__xor2_1 _14413_ (.A(_07539_),
    .B(_07563_),
    .X(_07564_));
 sky130_fd_sc_hd__nor2_1 _14414_ (.A(_07539_),
    .B(_07563_),
    .Y(_07565_));
 sky130_fd_sc_hd__a21oi_1 _14415_ (.A1(_07538_),
    .A2(_07564_),
    .B1(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__nor2_1 _14416_ (.A(_07519_),
    .B(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__xor2_2 _14417_ (.A(_07462_),
    .B(_07511_),
    .X(_07568_));
 sky130_fd_sc_hd__and2_1 _14418_ (.A(_07567_),
    .B(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__xnor2_1 _14419_ (.A(_07538_),
    .B(_07564_),
    .Y(_07570_));
 sky130_fd_sc_hd__nor2_1 _14420_ (.A(_07066_),
    .B(_07296_),
    .Y(_07571_));
 sky130_fd_sc_hd__nand2_1 _14421_ (.A(_07522_),
    .B(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__nor2_1 _14422_ (.A(_07326_),
    .B(_07296_),
    .Y(_07573_));
 sky130_fd_sc_hd__xnor2_1 _14423_ (.A(_07520_),
    .B(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__nor2_1 _14424_ (.A(_06832_),
    .B(_07301_),
    .Y(_07575_));
 sky130_fd_sc_hd__nand2_1 _14425_ (.A(_07574_),
    .B(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__xnor2_1 _14426_ (.A(_07531_),
    .B(_07533_),
    .Y(_07577_));
 sky130_fd_sc_hd__a21o_1 _14427_ (.A1(_07572_),
    .A2(_07576_),
    .B1(_07577_),
    .X(_07578_));
 sky130_fd_sc_hd__nand3_1 _14428_ (.A(_07572_),
    .B(_07576_),
    .C(_07577_),
    .Y(_07579_));
 sky130_fd_sc_hd__nand2_1 _14429_ (.A(_07578_),
    .B(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__nor2_1 _14430_ (.A(_07278_),
    .B(_07466_),
    .Y(_07581_));
 sky130_fd_sc_hd__nor2_1 _14431_ (.A(_06942_),
    .B(_07403_),
    .Y(_07582_));
 sky130_fd_sc_hd__inv_2 _14432_ (.A(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__nor2_1 _14433_ (.A(_07529_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__nor2_1 _14434_ (.A(_07530_),
    .B(_07582_),
    .Y(_07585_));
 sky130_fd_sc_hd__nor2_1 _14435_ (.A(_07584_),
    .B(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__a21oi_1 _14436_ (.A1(_07581_),
    .A2(_07586_),
    .B1(_07584_),
    .Y(_07587_));
 sky130_fd_sc_hd__or2_1 _14437_ (.A(_07580_),
    .B(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__o22a_1 _14438_ (.A1(_06703_),
    .A2(_07466_),
    .B1(_07404_),
    .B2(_06697_),
    .X(_07589_));
 sky130_fd_sc_hd__or2_1 _14439_ (.A(_07468_),
    .B(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__a21oi_2 _14440_ (.A1(_07578_),
    .A2(_07588_),
    .B1(_07590_),
    .Y(_07591_));
 sky130_fd_sc_hd__xnor2_2 _14441_ (.A(_07541_),
    .B(_07561_),
    .Y(_07592_));
 sky130_fd_sc_hd__and3_1 _14442_ (.A(_07578_),
    .B(_07588_),
    .C(_07590_),
    .X(_07593_));
 sky130_fd_sc_hd__nor2_1 _14443_ (.A(_07591_),
    .B(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__xnor2_1 _14444_ (.A(_07543_),
    .B(_07558_),
    .Y(_07595_));
 sky130_fd_sc_hd__xor2_1 _14445_ (.A(_07580_),
    .B(_07587_),
    .X(_07596_));
 sky130_fd_sc_hd__xnor2_1 _14446_ (.A(_07549_),
    .B(_07555_),
    .Y(_07597_));
 sky130_fd_sc_hd__or2_1 _14447_ (.A(_07574_),
    .B(_07575_),
    .X(_07598_));
 sky130_fd_sc_hd__and2_1 _14448_ (.A(_07576_),
    .B(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__xnor2_1 _14449_ (.A(_07552_),
    .B(_07553_),
    .Y(_07600_));
 sky130_fd_sc_hd__nor2_1 _14450_ (.A(_06799_),
    .B(_07284_),
    .Y(_07601_));
 sky130_fd_sc_hd__a2bb2o_1 _14451_ (.A1_N(_07244_),
    .A2_N(_07044_),
    .B1(_06769_),
    .B2(_07262_),
    .X(_07602_));
 sky130_fd_sc_hd__or4b_1 _14452_ (.A(_07051_),
    .B(_07244_),
    .C(_07044_),
    .D_N(_07261_),
    .X(_07603_));
 sky130_fd_sc_hd__a21bo_1 _14453_ (.A1(_07601_),
    .A2(_07602_),
    .B1_N(_07603_),
    .X(_07604_));
 sky130_fd_sc_hd__xnor2_1 _14454_ (.A(_07600_),
    .B(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__and2b_1 _14455_ (.A_N(_07600_),
    .B(_07604_),
    .X(_07606_));
 sky130_fd_sc_hd__a21oi_1 _14456_ (.A1(_07599_),
    .A2(_07605_),
    .B1(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__xor2_1 _14457_ (.A(_07597_),
    .B(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__nor2_1 _14458_ (.A(_07597_),
    .B(_07607_),
    .Y(_07609_));
 sky130_fd_sc_hd__a21oi_1 _14459_ (.A1(_07596_),
    .A2(_07608_),
    .B1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__xor2_1 _14460_ (.A(_07595_),
    .B(_07610_),
    .X(_07611_));
 sky130_fd_sc_hd__nor2_1 _14461_ (.A(_07595_),
    .B(_07610_),
    .Y(_07612_));
 sky130_fd_sc_hd__a21oi_2 _14462_ (.A1(_07594_),
    .A2(_07611_),
    .B1(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__xor2_2 _14463_ (.A(_07592_),
    .B(_07613_),
    .X(_07614_));
 sky130_fd_sc_hd__nor2_1 _14464_ (.A(_07592_),
    .B(_07613_),
    .Y(_07615_));
 sky130_fd_sc_hd__a21oi_1 _14465_ (.A1(_07591_),
    .A2(_07614_),
    .B1(_07615_),
    .Y(_07616_));
 sky130_fd_sc_hd__nor2_1 _14466_ (.A(_07570_),
    .B(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__xor2_1 _14467_ (.A(_07519_),
    .B(_07566_),
    .X(_07618_));
 sky130_fd_sc_hd__and2_1 _14468_ (.A(_07617_),
    .B(_07618_),
    .X(_07619_));
 sky130_fd_sc_hd__xnor2_2 _14469_ (.A(_07591_),
    .B(_07614_),
    .Y(_07620_));
 sky130_fd_sc_hd__nor2_1 _14470_ (.A(_07326_),
    .B(_07300_),
    .Y(_07621_));
 sky130_fd_sc_hd__nand2_1 _14471_ (.A(_07571_),
    .B(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__or2_1 _14472_ (.A(_07571_),
    .B(_07621_),
    .X(_07623_));
 sky130_fd_sc_hd__nand2_1 _14473_ (.A(_07622_),
    .B(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__or3_1 _14474_ (.A(_07331_),
    .B(_07355_),
    .C(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__xnor2_1 _14475_ (.A(_07581_),
    .B(_07586_),
    .Y(_07626_));
 sky130_fd_sc_hd__a21o_1 _14476_ (.A1(_07622_),
    .A2(_07625_),
    .B1(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__nand3_1 _14477_ (.A(_07622_),
    .B(_07625_),
    .C(_07626_),
    .Y(_07628_));
 sky130_fd_sc_hd__nand2_1 _14478_ (.A(_07627_),
    .B(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__or2_1 _14479_ (.A(_07217_),
    .B(_07466_),
    .X(_07630_));
 sky130_fd_sc_hd__o31a_1 _14480_ (.A1(_07583_),
    .A2(_07629_),
    .A3(_07630_),
    .B1(_07627_),
    .X(_07631_));
 sky130_fd_sc_hd__nor2b_1 _14481_ (.A(_07631_),
    .B_N(_07467_),
    .Y(_07632_));
 sky130_fd_sc_hd__xnor2_1 _14482_ (.A(_07594_),
    .B(_07611_),
    .Y(_07633_));
 sky130_fd_sc_hd__and2b_1 _14483_ (.A_N(_07467_),
    .B(_07631_),
    .X(_07634_));
 sky130_fd_sc_hd__nor2_1 _14484_ (.A(_07632_),
    .B(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__xnor2_1 _14485_ (.A(_07596_),
    .B(_07608_),
    .Y(_07636_));
 sky130_fd_sc_hd__nor2_1 _14486_ (.A(_07583_),
    .B(_07630_),
    .Y(_07637_));
 sky130_fd_sc_hd__xnor2_1 _14487_ (.A(_07629_),
    .B(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__xnor2_1 _14488_ (.A(_07599_),
    .B(_07605_),
    .Y(_07639_));
 sky130_fd_sc_hd__nor2_1 _14489_ (.A(_07331_),
    .B(_07355_),
    .Y(_07640_));
 sky130_fd_sc_hd__xnor2_1 _14490_ (.A(_07624_),
    .B(_07640_),
    .Y(_07641_));
 sky130_fd_sc_hd__nand3_1 _14491_ (.A(_07603_),
    .B(_07601_),
    .C(_07602_),
    .Y(_07642_));
 sky130_fd_sc_hd__a21o_1 _14492_ (.A1(_07603_),
    .A2(_07602_),
    .B1(_07601_),
    .X(_07643_));
 sky130_fd_sc_hd__nor2_1 _14493_ (.A(_06799_),
    .B(_07296_),
    .Y(_07644_));
 sky130_fd_sc_hd__o22ai_2 _14494_ (.A1(_07044_),
    .A2(_07284_),
    .B1(_07245_),
    .B2(_07051_),
    .Y(_07645_));
 sky130_fd_sc_hd__or4_1 _14495_ (.A(_07051_),
    .B(_07044_),
    .C(_07284_),
    .D(_07244_),
    .X(_07646_));
 sky130_fd_sc_hd__a21bo_1 _14496_ (.A1(_07644_),
    .A2(_07645_),
    .B1_N(_07646_),
    .X(_07647_));
 sky130_fd_sc_hd__a21o_1 _14497_ (.A1(_07642_),
    .A2(_07643_),
    .B1(_07647_),
    .X(_07648_));
 sky130_fd_sc_hd__nand3_1 _14498_ (.A(_07642_),
    .B(_07643_),
    .C(_07647_),
    .Y(_07649_));
 sky130_fd_sc_hd__a21boi_1 _14499_ (.A1(_07641_),
    .A2(_07648_),
    .B1_N(_07649_),
    .Y(_07650_));
 sky130_fd_sc_hd__xor2_1 _14500_ (.A(_07639_),
    .B(_07650_),
    .X(_07651_));
 sky130_fd_sc_hd__nor2_1 _14501_ (.A(_07639_),
    .B(_07650_),
    .Y(_07652_));
 sky130_fd_sc_hd__a21o_1 _14502_ (.A1(_07638_),
    .A2(_07651_),
    .B1(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__xnor2_1 _14503_ (.A(_07636_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__or2b_1 _14504_ (.A(_07636_),
    .B_N(_07653_),
    .X(_07655_));
 sky130_fd_sc_hd__a21boi_1 _14505_ (.A1(_07635_),
    .A2(_07654_),
    .B1_N(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__xor2_1 _14506_ (.A(_07633_),
    .B(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__nor2_1 _14507_ (.A(_07633_),
    .B(_07656_),
    .Y(_07658_));
 sky130_fd_sc_hd__a21oi_2 _14508_ (.A1(_07632_),
    .A2(_07657_),
    .B1(_07658_),
    .Y(_07659_));
 sky130_fd_sc_hd__nor2_1 _14509_ (.A(_07620_),
    .B(_07659_),
    .Y(_07660_));
 sky130_fd_sc_hd__xor2_1 _14510_ (.A(_07570_),
    .B(_07616_),
    .X(_07661_));
 sky130_fd_sc_hd__and2_1 _14511_ (.A(_07660_),
    .B(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__xor2_2 _14512_ (.A(_07620_),
    .B(_07659_),
    .X(_07663_));
 sky130_fd_sc_hd__nor2_1 _14513_ (.A(_07066_),
    .B(_07355_),
    .Y(_07664_));
 sky130_fd_sc_hd__nand2_1 _14514_ (.A(_07621_),
    .B(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__o22a_1 _14515_ (.A1(_07066_),
    .A2(_07301_),
    .B1(_07355_),
    .B2(_07326_),
    .X(_07666_));
 sky130_fd_sc_hd__a21o_1 _14516_ (.A1(_07621_),
    .A2(_07664_),
    .B1(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__or3_1 _14517_ (.A(_07331_),
    .B(_07404_),
    .C(_07667_),
    .X(_07668_));
 sky130_fd_sc_hd__o22a_1 _14518_ (.A1(_06942_),
    .A2(_07466_),
    .B1(_07404_),
    .B2(_07217_),
    .X(_07669_));
 sky130_fd_sc_hd__or2_1 _14519_ (.A(_07637_),
    .B(_07669_),
    .X(_07670_));
 sky130_fd_sc_hd__a21oi_2 _14520_ (.A1(_07665_),
    .A2(_07668_),
    .B1(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__xnor2_1 _14521_ (.A(_07638_),
    .B(_07651_),
    .Y(_07672_));
 sky130_fd_sc_hd__and3_1 _14522_ (.A(_07665_),
    .B(_07668_),
    .C(_07670_),
    .X(_07673_));
 sky130_fd_sc_hd__nor2_1 _14523_ (.A(_07671_),
    .B(_07673_),
    .Y(_07674_));
 sky130_fd_sc_hd__nand3_1 _14524_ (.A(_07649_),
    .B(_07641_),
    .C(_07648_),
    .Y(_07675_));
 sky130_fd_sc_hd__a21o_1 _14525_ (.A1(_07649_),
    .A2(_07648_),
    .B1(_07641_),
    .X(_07676_));
 sky130_fd_sc_hd__nand3_1 _14526_ (.A(_07646_),
    .B(_07644_),
    .C(_07645_),
    .Y(_07677_));
 sky130_fd_sc_hd__a21o_1 _14527_ (.A1(_07646_),
    .A2(_07645_),
    .B1(_07644_),
    .X(_07678_));
 sky130_fd_sc_hd__nor2_1 _14528_ (.A(_07044_),
    .B(_07296_),
    .Y(_07679_));
 sky130_fd_sc_hd__and3b_1 _14529_ (.A_N(_07283_),
    .B(_07679_),
    .C(_06769_),
    .X(_07680_));
 sky130_fd_sc_hd__or2_1 _14530_ (.A(_06799_),
    .B(_07301_),
    .X(_07681_));
 sky130_fd_sc_hd__o21ba_1 _14531_ (.A1(_07051_),
    .A2(_07284_),
    .B1_N(_07679_),
    .X(_07682_));
 sky130_fd_sc_hd__or3_1 _14532_ (.A(_07680_),
    .B(_07681_),
    .C(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__or2b_1 _14533_ (.A(_07680_),
    .B_N(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__nand3_1 _14534_ (.A(_07677_),
    .B(_07678_),
    .C(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__nor2_1 _14535_ (.A(_07331_),
    .B(_07404_),
    .Y(_07686_));
 sky130_fd_sc_hd__xnor2_1 _14536_ (.A(_07667_),
    .B(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__a21o_1 _14537_ (.A1(_07677_),
    .A2(_07678_),
    .B1(_07684_),
    .X(_07688_));
 sky130_fd_sc_hd__and3_1 _14538_ (.A(_07685_),
    .B(_07687_),
    .C(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__a31o_1 _14539_ (.A1(_07677_),
    .A2(_07678_),
    .A3(_07684_),
    .B1(_07689_),
    .X(_07690_));
 sky130_fd_sc_hd__and3_1 _14540_ (.A(_07675_),
    .B(_07676_),
    .C(_07690_),
    .X(_07691_));
 sky130_fd_sc_hd__a21oi_1 _14541_ (.A1(_07675_),
    .A2(_07676_),
    .B1(_07690_),
    .Y(_07692_));
 sky130_fd_sc_hd__nor2_1 _14542_ (.A(_07691_),
    .B(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__a21oi_1 _14543_ (.A1(_07674_),
    .A2(_07693_),
    .B1(_07691_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand2_1 _14544_ (.A(_07672_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__nor2_1 _14545_ (.A(_07672_),
    .B(_07694_),
    .Y(_07696_));
 sky130_fd_sc_hd__a21oi_2 _14546_ (.A1(_07671_),
    .A2(_07695_),
    .B1(_07696_),
    .Y(_07697_));
 sky130_fd_sc_hd__xnor2_1 _14547_ (.A(_07635_),
    .B(_07654_),
    .Y(_07698_));
 sky130_fd_sc_hd__xor2_1 _14548_ (.A(_07632_),
    .B(_07657_),
    .X(_07699_));
 sky130_fd_sc_hd__nor3b_2 _14549_ (.A(_07697_),
    .B(_07698_),
    .C_N(_07699_),
    .Y(_07700_));
 sky130_fd_sc_hd__and2_1 _14550_ (.A(_07663_),
    .B(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__xor2_2 _14551_ (.A(_07663_),
    .B(_07700_),
    .X(_07702_));
 sky130_fd_sc_hd__and2b_1 _14552_ (.A_N(_07696_),
    .B(_07695_),
    .X(_07703_));
 sky130_fd_sc_hd__xor2_1 _14553_ (.A(_07671_),
    .B(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__xnor2_1 _14554_ (.A(_07674_),
    .B(_07693_),
    .Y(_07705_));
 sky130_fd_sc_hd__nor2_1 _14555_ (.A(_07326_),
    .B(_07404_),
    .Y(_07706_));
 sky130_fd_sc_hd__nand2_1 _14556_ (.A(_07664_),
    .B(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__or2_1 _14557_ (.A(_07664_),
    .B(_07706_),
    .X(_07708_));
 sky130_fd_sc_hd__nand2_1 _14558_ (.A(_07707_),
    .B(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__o31a_1 _14559_ (.A1(_07331_),
    .A2(_07466_),
    .A3(_07709_),
    .B1(_07707_),
    .X(_07710_));
 sky130_fd_sc_hd__nor2_1 _14560_ (.A(_07630_),
    .B(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__and2_1 _14561_ (.A(_07630_),
    .B(_07710_),
    .X(_07712_));
 sky130_fd_sc_hd__nor2_1 _14562_ (.A(_07711_),
    .B(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__a21oi_1 _14563_ (.A1(_07685_),
    .A2(_07688_),
    .B1(_07687_),
    .Y(_07714_));
 sky130_fd_sc_hd__nor2_1 _14564_ (.A(_07331_),
    .B(_07466_),
    .Y(_07715_));
 sky130_fd_sc_hd__xnor2_1 _14565_ (.A(_07709_),
    .B(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__o21ai_1 _14566_ (.A1(_07680_),
    .A2(_07682_),
    .B1(_07681_),
    .Y(_07717_));
 sky130_fd_sc_hd__nor2_1 _14567_ (.A(_07051_),
    .B(_07301_),
    .Y(_07718_));
 sky130_fd_sc_hd__nor2_1 _14568_ (.A(_06799_),
    .B(_07355_),
    .Y(_07719_));
 sky130_fd_sc_hd__o22a_1 _14569_ (.A1(_07051_),
    .A2(_07296_),
    .B1(_07301_),
    .B2(_07044_),
    .X(_07720_));
 sky130_fd_sc_hd__a21oi_1 _14570_ (.A1(_07679_),
    .A2(_07718_),
    .B1(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__a22o_1 _14571_ (.A1(_07679_),
    .A2(_07718_),
    .B1(_07719_),
    .B2(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__a21o_1 _14572_ (.A1(_07683_),
    .A2(_07717_),
    .B1(_07722_),
    .X(_07723_));
 sky130_fd_sc_hd__and3_1 _14573_ (.A(_07683_),
    .B(_07717_),
    .C(_07722_),
    .X(_07724_));
 sky130_fd_sc_hd__a21oi_1 _14574_ (.A1(_07716_),
    .A2(_07723_),
    .B1(_07724_),
    .Y(_07725_));
 sky130_fd_sc_hd__o21ai_1 _14575_ (.A1(_07689_),
    .A2(_07714_),
    .B1(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__or3_1 _14576_ (.A(_07689_),
    .B(_07714_),
    .C(_07725_),
    .X(_07727_));
 sky130_fd_sc_hd__a21boi_1 _14577_ (.A1(_07713_),
    .A2(_07726_),
    .B1_N(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__xor2_1 _14578_ (.A(_07705_),
    .B(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__nand2_1 _14579_ (.A(_07711_),
    .B(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__o21ai_1 _14580_ (.A1(_07705_),
    .A2(_07728_),
    .B1(_07730_),
    .Y(_07731_));
 sky130_fd_sc_hd__xor2_1 _14581_ (.A(_07698_),
    .B(_07697_),
    .X(_07732_));
 sky130_fd_sc_hd__and4_1 _14582_ (.A(_07699_),
    .B(_07704_),
    .C(_07731_),
    .D(_07732_),
    .X(_07733_));
 sky130_fd_sc_hd__xor2_2 _14583_ (.A(_07702_),
    .B(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__or2_1 _14584_ (.A(_07704_),
    .B(_07731_),
    .X(_07735_));
 sky130_fd_sc_hd__and2b_1 _14585_ (.A_N(_07724_),
    .B(_07723_),
    .X(_07736_));
 sky130_fd_sc_hd__xnor2_1 _14586_ (.A(_07716_),
    .B(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__xnor2_1 _14587_ (.A(_07719_),
    .B(_07721_),
    .Y(_07738_));
 sky130_fd_sc_hd__nor2_1 _14588_ (.A(_07044_),
    .B(_07355_),
    .Y(_07739_));
 sky130_fd_sc_hd__or2_1 _14589_ (.A(_06799_),
    .B(_07404_),
    .X(_07740_));
 sky130_fd_sc_hd__xnor2_1 _14590_ (.A(_07718_),
    .B(_07739_),
    .Y(_07741_));
 sky130_fd_sc_hd__or2_1 _14591_ (.A(_07740_),
    .B(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__a21bo_1 _14592_ (.A1(_07718_),
    .A2(_07739_),
    .B1_N(_07742_),
    .X(_07743_));
 sky130_fd_sc_hd__or2b_1 _14593_ (.A(_07738_),
    .B_N(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__or2_1 _14594_ (.A(_07066_),
    .B(_07466_),
    .X(_07745_));
 sky130_fd_sc_hd__nor3_1 _14595_ (.A(_07326_),
    .B(_07404_),
    .C(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__o22a_1 _14596_ (.A1(_07326_),
    .A2(_07466_),
    .B1(_07404_),
    .B2(_07066_),
    .X(_07747_));
 sky130_fd_sc_hd__nor2_1 _14597_ (.A(_07746_),
    .B(_07747_),
    .Y(_07748_));
 sky130_fd_sc_hd__xnor2_1 _14598_ (.A(_07738_),
    .B(_07743_),
    .Y(_07749_));
 sky130_fd_sc_hd__nand2_1 _14599_ (.A(_07748_),
    .B(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__nand2_1 _14600_ (.A(_07740_),
    .B(_07741_),
    .Y(_07751_));
 sky130_fd_sc_hd__and2_1 _14601_ (.A(_07742_),
    .B(_07751_),
    .X(_07752_));
 sky130_fd_sc_hd__or2_1 _14602_ (.A(_06799_),
    .B(_07466_),
    .X(_07753_));
 sky130_fd_sc_hd__or2_1 _14603_ (.A(_07051_),
    .B(_07355_),
    .X(_07754_));
 sky130_fd_sc_hd__or2_1 _14604_ (.A(_07044_),
    .B(_07404_),
    .X(_07755_));
 sky130_fd_sc_hd__xnor2_1 _14605_ (.A(_07754_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__nand2_1 _14606_ (.A(_07753_),
    .B(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__or2_1 _14607_ (.A(_07753_),
    .B(_07756_),
    .X(_07758_));
 sky130_fd_sc_hd__and4_1 _14608_ (.A(_07042_),
    .B(_07126_),
    .C(_07757_),
    .D(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__and2_1 _14609_ (.A(_07752_),
    .B(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__o21a_1 _14610_ (.A1(_07754_),
    .A2(_07755_),
    .B1(_07758_),
    .X(_07761_));
 sky130_fd_sc_hd__nand2_1 _14611_ (.A(_07745_),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__nor2_1 _14612_ (.A(_07745_),
    .B(_07761_),
    .Y(_07763_));
 sky130_fd_sc_hd__or3_1 _14613_ (.A(_07752_),
    .B(_07759_),
    .C(_07763_),
    .X(_07764_));
 sky130_fd_sc_hd__or2_1 _14614_ (.A(_07748_),
    .B(_07749_),
    .X(_07765_));
 sky130_fd_sc_hd__a22o_1 _14615_ (.A1(_07750_),
    .A2(_07765_),
    .B1(_07760_),
    .B2(_07763_),
    .X(_07766_));
 sky130_fd_sc_hd__o211a_1 _14616_ (.A1(_07760_),
    .A2(_07762_),
    .B1(_07764_),
    .C1(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__nor2_1 _14617_ (.A(_07746_),
    .B(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__a31o_1 _14618_ (.A1(_07737_),
    .A2(_07744_),
    .A3(_07750_),
    .B1(_07768_),
    .X(_07769_));
 sky130_fd_sc_hd__a21o_1 _14619_ (.A1(_07744_),
    .A2(_07750_),
    .B1(_07737_),
    .X(_07770_));
 sky130_fd_sc_hd__nand2_1 _14620_ (.A(_07746_),
    .B(_07767_),
    .Y(_07771_));
 sky130_fd_sc_hd__a21oi_1 _14621_ (.A1(_07727_),
    .A2(_07726_),
    .B1(_07713_),
    .Y(_07772_));
 sky130_fd_sc_hd__and3_1 _14622_ (.A(_07727_),
    .B(_07713_),
    .C(_07726_),
    .X(_07773_));
 sky130_fd_sc_hd__a311o_1 _14623_ (.A1(_07769_),
    .A2(_07770_),
    .A3(_07771_),
    .B1(_07772_),
    .C1(_07773_),
    .X(_07774_));
 sky130_fd_sc_hd__or2_1 _14624_ (.A(_07711_),
    .B(_07729_),
    .X(_07775_));
 sky130_fd_sc_hd__and3b_1 _14625_ (.A_N(_07774_),
    .B(_07775_),
    .C(_07730_),
    .X(_07776_));
 sky130_fd_sc_hd__and4_1 _14626_ (.A(_07699_),
    .B(_07732_),
    .C(_07735_),
    .D(_07776_),
    .X(_07777_));
 sky130_fd_sc_hd__and2_1 _14627_ (.A(_07702_),
    .B(_07733_),
    .X(_07778_));
 sky130_fd_sc_hd__a21o_1 _14628_ (.A1(_07734_),
    .A2(_07777_),
    .B1(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__nor2_1 _14629_ (.A(_07660_),
    .B(_07701_),
    .Y(_07780_));
 sky130_fd_sc_hd__xnor2_1 _14630_ (.A(_07661_),
    .B(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__a22o_1 _14631_ (.A1(_07701_),
    .A2(_07661_),
    .B1(_07779_),
    .B2(_07781_),
    .X(_07782_));
 sky130_fd_sc_hd__nor2_1 _14632_ (.A(_07617_),
    .B(_07662_),
    .Y(_07783_));
 sky130_fd_sc_hd__xnor2_1 _14633_ (.A(_07618_),
    .B(_07783_),
    .Y(_07784_));
 sky130_fd_sc_hd__a22o_1 _14634_ (.A1(_07618_),
    .A2(_07662_),
    .B1(_07782_),
    .B2(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__nor3_1 _14635_ (.A(_07567_),
    .B(_07568_),
    .C(_07619_),
    .Y(_07786_));
 sky130_fd_sc_hd__a211oi_2 _14636_ (.A1(_07568_),
    .A2(_07619_),
    .B1(_07786_),
    .C1(_07569_),
    .Y(_07787_));
 sky130_fd_sc_hd__a22o_1 _14637_ (.A1(_07568_),
    .A2(_07619_),
    .B1(_07785_),
    .B2(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__nor2_1 _14638_ (.A(_07512_),
    .B(_07569_),
    .Y(_07789_));
 sky130_fd_sc_hd__xnor2_1 _14639_ (.A(_07514_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__a22oi_2 _14640_ (.A1(_07514_),
    .A2(_07569_),
    .B1(_07788_),
    .B2(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__o21a_1 _14641_ (.A1(_07457_),
    .A2(_07515_),
    .B1(_07400_),
    .X(_07792_));
 sky130_fd_sc_hd__inv_2 _14642_ (.A(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__o31a_2 _14643_ (.A1(_07459_),
    .A2(_07518_),
    .A3(_07791_),
    .B1(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__nor2_1 _14644_ (.A(_07292_),
    .B(_07398_),
    .Y(_07795_));
 sky130_fd_sc_hd__o21bai_2 _14645_ (.A1(_07397_),
    .A2(_07794_),
    .B1_N(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__xnor2_2 _14646_ (.A(_07350_),
    .B(_07796_),
    .Y(_07797_));
 sky130_fd_sc_hd__xnor2_1 _14647_ (.A(_07397_),
    .B(_07794_),
    .Y(_07798_));
 sky130_fd_sc_hd__nor2_1 _14648_ (.A(_06555_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__or2_1 _14649_ (.A(_06547_),
    .B(_06565_),
    .X(_07800_));
 sky130_fd_sc_hd__buf_2 _14650_ (.A(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__a211o_1 _14651_ (.A1(_06555_),
    .A2(_07797_),
    .B1(_07799_),
    .C1(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__buf_2 _14652_ (.A(_06628_),
    .X(_07803_));
 sky130_fd_sc_hd__or3b_1 _14653_ (.A(_07292_),
    .B(_07395_),
    .C_N(_07348_),
    .X(_07804_));
 sky130_fd_sc_hd__o31a_2 _14654_ (.A1(_07397_),
    .A2(_07794_),
    .A3(_07350_),
    .B1(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__o21ai_2 _14655_ (.A1(_06703_),
    .A2(_07270_),
    .B1(_07287_),
    .Y(_07806_));
 sky130_fd_sc_hd__nor4_4 _14656_ (.A(_06545_),
    .B(_07272_),
    .C(_07347_),
    .D(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__xor2_2 _14657_ (.A(_07805_),
    .B(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__nor3_2 _14658_ (.A(_07803_),
    .B(_07805_),
    .C(_07807_),
    .Y(_07809_));
 sky130_fd_sc_hd__a211o_1 _14659_ (.A1(_07803_),
    .A2(_07808_),
    .B1(_07809_),
    .C1(_06566_),
    .X(_07810_));
 sky130_fd_sc_hd__buf_2 _14660_ (.A(_06644_),
    .X(_07811_));
 sky130_fd_sc_hd__a21oi_1 _14661_ (.A1(_07802_),
    .A2(_07810_),
    .B1(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__xnor2_2 _14662_ (.A(_07785_),
    .B(_07787_),
    .Y(_07813_));
 sky130_fd_sc_hd__xnor2_1 _14663_ (.A(_07788_),
    .B(_07790_),
    .Y(_07814_));
 sky130_fd_sc_hd__nor2_1 _14664_ (.A(_06628_),
    .B(_07814_),
    .Y(_07815_));
 sky130_fd_sc_hd__o21ba_1 _14665_ (.A1(_06554_),
    .A2(_07813_),
    .B1_N(_07815_),
    .X(_07816_));
 sky130_fd_sc_hd__clkinv_2 _14666_ (.A(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__o21bai_1 _14667_ (.A1(_07518_),
    .A2(_07791_),
    .B1_N(_07515_),
    .Y(_07818_));
 sky130_fd_sc_hd__xnor2_2 _14668_ (.A(_07459_),
    .B(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__xnor2_1 _14669_ (.A(_07517_),
    .B(_07791_),
    .Y(_07820_));
 sky130_fd_sc_hd__mux2_1 _14670_ (.A0(_07819_),
    .A1(_07820_),
    .S(_06628_),
    .X(_07821_));
 sky130_fd_sc_hd__mux2_1 _14671_ (.A0(_07817_),
    .A1(_07821_),
    .S(_07801_),
    .X(_07822_));
 sky130_fd_sc_hd__xnor2_2 _14672_ (.A(_07734_),
    .B(_07777_),
    .Y(_07823_));
 sky130_fd_sc_hd__or2_1 _14673_ (.A(_07803_),
    .B(_07823_),
    .X(_07824_));
 sky130_fd_sc_hd__xnor2_1 _14674_ (.A(_07782_),
    .B(_07784_),
    .Y(_07825_));
 sky130_fd_sc_hd__or2_1 _14675_ (.A(_06628_),
    .B(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__xor2_1 _14676_ (.A(_07779_),
    .B(_07781_),
    .X(_07827_));
 sky130_fd_sc_hd__nand2_1 _14677_ (.A(_06628_),
    .B(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__and2_1 _14678_ (.A(_07826_),
    .B(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__mux2_1 _14679_ (.A0(_07824_),
    .A1(_07829_),
    .S(_07801_),
    .X(_07830_));
 sky130_fd_sc_hd__nand2_1 _14680_ (.A(_06549_),
    .B(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__o211ai_1 _14681_ (.A1(_06549_),
    .A2(_07822_),
    .B1(_07831_),
    .C1(_06544_),
    .Y(_07832_));
 sky130_fd_sc_hd__o31ai_1 _14682_ (.A1(_06544_),
    .A2(_06550_),
    .A3(_07812_),
    .B1(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__clkbuf_4 _14683_ (.A(_06602_),
    .X(_07834_));
 sky130_fd_sc_hd__a21o_1 _14684_ (.A1(_06461_),
    .A2(_07833_),
    .B1(_07834_),
    .X(_07835_));
 sky130_fd_sc_hd__and4b_1 _14685_ (.A_N(_04472_),
    .B(_04471_),
    .C(_04468_),
    .D(_06157_),
    .X(_07836_));
 sky130_fd_sc_hd__buf_2 _14686_ (.A(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__clkbuf_4 _14687_ (.A(_07837_),
    .X(_07838_));
 sky130_fd_sc_hd__mux2_1 _14688_ (.A0(\rbzero.wall_tracer.stepDistY[-11] ),
    .A1(_07835_),
    .S(_07838_),
    .X(_07839_));
 sky130_fd_sc_hd__clkbuf_1 _14689_ (.A(_07839_),
    .X(_00391_));
 sky130_fd_sc_hd__nor3_2 _14690_ (.A(_06555_),
    .B(_07805_),
    .C(_07807_),
    .Y(_07840_));
 sky130_fd_sc_hd__mux2_1 _14691_ (.A0(_07808_),
    .A1(_07797_),
    .S(_07803_),
    .X(_07841_));
 sky130_fd_sc_hd__mux2_1 _14692_ (.A0(_07840_),
    .A1(_07841_),
    .S(_06566_),
    .X(_07842_));
 sky130_fd_sc_hd__a21oi_1 _14693_ (.A1(_06549_),
    .A2(_07842_),
    .B1(_06544_),
    .Y(_07843_));
 sky130_fd_sc_hd__and2_1 _14694_ (.A(_06523_),
    .B(_06543_),
    .X(_07844_));
 sky130_fd_sc_hd__or2_2 _14695_ (.A(_06527_),
    .B(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__nor2_1 _14696_ (.A(_06554_),
    .B(_07814_),
    .Y(_07846_));
 sky130_fd_sc_hd__and2_1 _14697_ (.A(_06554_),
    .B(_07820_),
    .X(_07847_));
 sky130_fd_sc_hd__or2_1 _14698_ (.A(_07846_),
    .B(_07847_),
    .X(_07848_));
 sky130_fd_sc_hd__xnor2_1 _14699_ (.A(_07396_),
    .B(_07794_),
    .Y(_07849_));
 sky130_fd_sc_hd__mux2_1 _14700_ (.A0(_07849_),
    .A1(_07819_),
    .S(_06628_),
    .X(_07850_));
 sky130_fd_sc_hd__mux2_1 _14701_ (.A0(_07848_),
    .A1(_07850_),
    .S(_07801_),
    .X(_07851_));
 sky130_fd_sc_hd__nor2_1 _14702_ (.A(_06628_),
    .B(_07813_),
    .Y(_07852_));
 sky130_fd_sc_hd__nor2_1 _14703_ (.A(_06554_),
    .B(_07825_),
    .Y(_07853_));
 sky130_fd_sc_hd__nor2_1 _14704_ (.A(_07852_),
    .B(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__and2_1 _14705_ (.A(_06554_),
    .B(_07827_),
    .X(_07855_));
 sky130_fd_sc_hd__o21bai_1 _14706_ (.A1(_06554_),
    .A2(_07823_),
    .B1_N(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__nor2_1 _14707_ (.A(_07801_),
    .B(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__a21oi_2 _14708_ (.A1(_07801_),
    .A2(_07854_),
    .B1(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__or2_1 _14709_ (.A(_06644_),
    .B(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__o21a_1 _14710_ (.A1(_06549_),
    .A2(_07851_),
    .B1(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__nor2_1 _14711_ (.A(_07845_),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__nor2_2 _14712_ (.A(_06545_),
    .B(_06494_),
    .Y(_07862_));
 sky130_fd_sc_hd__buf_4 _14713_ (.A(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__o31ai_4 _14714_ (.A1(_06669_),
    .A2(_07843_),
    .A3(_07861_),
    .B1(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__mux2_1 _14715_ (.A0(\rbzero.wall_tracer.stepDistY[-10] ),
    .A1(_07864_),
    .S(_07838_),
    .X(_07865_));
 sky130_fd_sc_hd__clkbuf_1 _14716_ (.A(_07865_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _14717_ (.A0(_07808_),
    .A1(_07797_),
    .S(_06555_),
    .X(_07866_));
 sky130_fd_sc_hd__or3_1 _14718_ (.A(_06545_),
    .B(_06687_),
    .C(_07809_),
    .X(_07867_));
 sky130_fd_sc_hd__o211a_1 _14719_ (.A1(_06587_),
    .A2(_07866_),
    .B1(_07867_),
    .C1(_06603_),
    .X(_07868_));
 sky130_fd_sc_hd__buf_2 _14720_ (.A(_06587_),
    .X(_07869_));
 sky130_fd_sc_hd__mux2_1 _14721_ (.A0(_07849_),
    .A1(_07819_),
    .S(_06555_),
    .X(_07870_));
 sky130_fd_sc_hd__a21oi_1 _14722_ (.A1(_07803_),
    .A2(_07820_),
    .B1(_07815_),
    .Y(_07871_));
 sky130_fd_sc_hd__nor2_1 _14723_ (.A(_06587_),
    .B(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__buf_2 _14724_ (.A(_06603_),
    .X(_07873_));
 sky130_fd_sc_hd__a211o_1 _14725_ (.A1(_07869_),
    .A2(_07870_),
    .B1(_07872_),
    .C1(_07873_),
    .X(_07874_));
 sky130_fd_sc_hd__o21ai_1 _14726_ (.A1(_06555_),
    .A2(_07813_),
    .B1(_07826_),
    .Y(_07875_));
 sky130_fd_sc_hd__or2_1 _14727_ (.A(_06638_),
    .B(_07875_),
    .X(_07876_));
 sky130_fd_sc_hd__or2_1 _14728_ (.A(_06669_),
    .B(_06523_),
    .X(_07877_));
 sky130_fd_sc_hd__a31oi_1 _14729_ (.A1(_06573_),
    .A2(_07828_),
    .A3(_07824_),
    .B1(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__a31o_1 _14730_ (.A1(_07874_),
    .A2(_07876_),
    .A3(_07878_),
    .B1(_07834_),
    .X(_07879_));
 sky130_fd_sc_hd__a21o_2 _14731_ (.A1(_06508_),
    .A2(_07868_),
    .B1(_07879_),
    .X(_07880_));
 sky130_fd_sc_hd__mux2_1 _14732_ (.A0(\rbzero.wall_tracer.stepDistY[-9] ),
    .A1(_07880_),
    .S(_07838_),
    .X(_07881_));
 sky130_fd_sc_hd__clkbuf_1 _14733_ (.A(_07881_),
    .X(_00393_));
 sky130_fd_sc_hd__nor2_1 _14734_ (.A(_07803_),
    .B(_07798_),
    .Y(_07882_));
 sky130_fd_sc_hd__a21oi_1 _14735_ (.A1(_07803_),
    .A2(_07797_),
    .B1(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__a21oi_1 _14736_ (.A1(_07803_),
    .A2(_07819_),
    .B1(_07847_),
    .Y(_07884_));
 sky130_fd_sc_hd__and2_1 _14737_ (.A(_06687_),
    .B(_07884_),
    .X(_07885_));
 sky130_fd_sc_hd__a211o_1 _14738_ (.A1(_07869_),
    .A2(_07883_),
    .B1(_07885_),
    .C1(_07873_),
    .X(_07886_));
 sky130_fd_sc_hd__or2_1 _14739_ (.A(_07846_),
    .B(_07852_),
    .X(_07887_));
 sky130_fd_sc_hd__inv_2 _14740_ (.A(_07887_),
    .Y(_07888_));
 sky130_fd_sc_hd__nor2_1 _14741_ (.A(_07853_),
    .B(_07855_),
    .Y(_07889_));
 sky130_fd_sc_hd__o221a_1 _14742_ (.A1(_06638_),
    .A2(_07888_),
    .B1(_07889_),
    .B2(_06619_),
    .C1(_06595_),
    .X(_07890_));
 sky130_fd_sc_hd__a21o_1 _14743_ (.A1(_06555_),
    .A2(_07808_),
    .B1(_07840_),
    .X(_07891_));
 sky130_fd_sc_hd__a21oi_1 _14744_ (.A1(_06573_),
    .A2(_07891_),
    .B1(_06595_),
    .Y(_07892_));
 sky130_fd_sc_hd__a211o_1 _14745_ (.A1(_07886_),
    .A2(_07890_),
    .B1(_07892_),
    .C1(_06669_),
    .X(_07893_));
 sky130_fd_sc_hd__and2_1 _14746_ (.A(_07801_),
    .B(_07856_),
    .X(_07894_));
 sky130_fd_sc_hd__nand2_1 _14747_ (.A(_07811_),
    .B(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__o21a_1 _14748_ (.A1(_06556_),
    .A2(_07895_),
    .B1(_07863_),
    .X(_07896_));
 sky130_fd_sc_hd__nand2_1 _14749_ (.A(_07893_),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__mux2_1 _14750_ (.A0(\rbzero.wall_tracer.stepDistY[-8] ),
    .A1(_07897_),
    .S(_07838_),
    .X(_07898_));
 sky130_fd_sc_hd__clkbuf_1 _14751_ (.A(_07898_),
    .X(_00394_));
 sky130_fd_sc_hd__or2_1 _14752_ (.A(_06545_),
    .B(_07809_),
    .X(_07899_));
 sky130_fd_sc_hd__and2_1 _14753_ (.A(_06573_),
    .B(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__nand2_1 _14754_ (.A(_07869_),
    .B(_07871_),
    .Y(_07901_));
 sky130_fd_sc_hd__o211a_1 _14755_ (.A1(_07869_),
    .A2(_07875_),
    .B1(_07901_),
    .C1(_07873_),
    .X(_07902_));
 sky130_fd_sc_hd__nor2_1 _14756_ (.A(_06523_),
    .B(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__xnor2_1 _14757_ (.A(_07805_),
    .B(_07807_),
    .Y(_07904_));
 sky130_fd_sc_hd__xnor2_1 _14758_ (.A(_07349_),
    .B(_07796_),
    .Y(_07905_));
 sky130_fd_sc_hd__mux2_1 _14759_ (.A0(_07904_),
    .A1(_07905_),
    .S(_06555_),
    .X(_07906_));
 sky130_fd_sc_hd__nor2_1 _14760_ (.A(_07869_),
    .B(_07870_),
    .Y(_07907_));
 sky130_fd_sc_hd__a211o_1 _14761_ (.A1(_07869_),
    .A2(_07906_),
    .B1(_07907_),
    .C1(_07873_),
    .X(_07908_));
 sky130_fd_sc_hd__a2bb2o_1 _14762_ (.A1_N(_06595_),
    .A2_N(_07900_),
    .B1(_07903_),
    .B2(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__o31a_1 _14763_ (.A1(_06461_),
    .A2(_06549_),
    .A3(_07830_),
    .B1(_07863_),
    .X(_07910_));
 sky130_fd_sc_hd__o21a_2 _14764_ (.A1(_06669_),
    .A2(_07909_),
    .B1(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__nor2_1 _14765_ (.A(\rbzero.wall_tracer.stepDistY[-7] ),
    .B(_07838_),
    .Y(_07912_));
 sky130_fd_sc_hd__a21oi_1 _14766_ (.A1(_07838_),
    .A2(_07911_),
    .B1(_07912_),
    .Y(_00395_));
 sky130_fd_sc_hd__a211o_1 _14767_ (.A1(_06555_),
    .A2(_07808_),
    .B1(_07840_),
    .C1(_06687_),
    .X(_07913_));
 sky130_fd_sc_hd__a211o_1 _14768_ (.A1(_07803_),
    .A2(_07797_),
    .B1(_07882_),
    .C1(_06587_),
    .X(_07914_));
 sky130_fd_sc_hd__a21o_1 _14769_ (.A1(_07913_),
    .A2(_07914_),
    .B1(_07873_),
    .X(_07915_));
 sky130_fd_sc_hd__mux2_1 _14770_ (.A0(_07888_),
    .A1(_07884_),
    .S(_07869_),
    .X(_07916_));
 sky130_fd_sc_hd__a21oi_1 _14771_ (.A1(_07873_),
    .A2(_07916_),
    .B1(_07877_),
    .Y(_07917_));
 sky130_fd_sc_hd__and3_1 _14772_ (.A(_06612_),
    .B(_07811_),
    .C(_07858_),
    .X(_07918_));
 sky130_fd_sc_hd__a21oi_2 _14773_ (.A1(_07915_),
    .A2(_07917_),
    .B1(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__nand2_1 _14774_ (.A(_07863_),
    .B(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__mux2_1 _14775_ (.A0(\rbzero.wall_tracer.stepDistY[-6] ),
    .A1(_07920_),
    .S(_07838_),
    .X(_07921_));
 sky130_fd_sc_hd__clkbuf_1 _14776_ (.A(_07921_),
    .X(_00396_));
 sky130_fd_sc_hd__o21a_1 _14777_ (.A1(_06545_),
    .A2(_07809_),
    .B1(_07869_),
    .X(_07922_));
 sky130_fd_sc_hd__a211o_1 _14778_ (.A1(_06687_),
    .A2(_07866_),
    .B1(_07922_),
    .C1(_07873_),
    .X(_07923_));
 sky130_fd_sc_hd__nor2_1 _14779_ (.A(_06669_),
    .B(_06523_),
    .Y(_07924_));
 sky130_fd_sc_hd__a211o_1 _14780_ (.A1(_07869_),
    .A2(_07870_),
    .B1(_07872_),
    .C1(_06585_),
    .X(_07925_));
 sky130_fd_sc_hd__and2_1 _14781_ (.A(_07924_),
    .B(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__mux2_1 _14782_ (.A0(_07829_),
    .A1(_07816_),
    .S(_07801_),
    .X(_07927_));
 sky130_fd_sc_hd__or2_1 _14783_ (.A(_06566_),
    .B(_07824_),
    .X(_07928_));
 sky130_fd_sc_hd__mux2_1 _14784_ (.A0(_07927_),
    .A1(_07928_),
    .S(_06548_),
    .X(_07929_));
 sky130_fd_sc_hd__o21ai_1 _14785_ (.A1(_06556_),
    .A2(_07929_),
    .B1(_07862_),
    .Y(_07930_));
 sky130_fd_sc_hd__a21oi_4 _14786_ (.A1(_07923_),
    .A2(_07926_),
    .B1(_07930_),
    .Y(_07931_));
 sky130_fd_sc_hd__nor2_1 _14787_ (.A(\rbzero.wall_tracer.stepDistY[-5] ),
    .B(_07838_),
    .Y(_07932_));
 sky130_fd_sc_hd__a21oi_1 _14788_ (.A1(_07838_),
    .A2(_07931_),
    .B1(_07932_),
    .Y(_00397_));
 sky130_fd_sc_hd__a21o_1 _14789_ (.A1(_07869_),
    .A2(_07883_),
    .B1(_07885_),
    .X(_07933_));
 sky130_fd_sc_hd__a21oi_1 _14790_ (.A1(_06687_),
    .A2(_07891_),
    .B1(_07873_),
    .Y(_07934_));
 sky130_fd_sc_hd__a211o_1 _14791_ (.A1(_07873_),
    .A2(_07933_),
    .B1(_07934_),
    .C1(_07877_),
    .X(_07935_));
 sky130_fd_sc_hd__nand2_1 _14792_ (.A(_06566_),
    .B(_07854_),
    .Y(_07936_));
 sky130_fd_sc_hd__o21a_1 _14793_ (.A1(_06566_),
    .A2(_07848_),
    .B1(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__mux2_1 _14794_ (.A0(_07894_),
    .A1(_07937_),
    .S(_07811_),
    .X(_07938_));
 sky130_fd_sc_hd__a21oi_1 _14795_ (.A1(_06612_),
    .A2(_07938_),
    .B1(_07834_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_1 _14796_ (.A(_07935_),
    .B(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__mux2_1 _14797_ (.A0(\rbzero.wall_tracer.stepDistY[-4] ),
    .A1(_07940_),
    .S(_07838_),
    .X(_07941_));
 sky130_fd_sc_hd__clkbuf_1 _14798_ (.A(_07941_),
    .X(_00398_));
 sky130_fd_sc_hd__o21ai_2 _14799_ (.A1(_06549_),
    .A2(_07822_),
    .B1(_07831_),
    .Y(_07942_));
 sky130_fd_sc_hd__or2_1 _14800_ (.A(_06556_),
    .B(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__a21oi_1 _14801_ (.A1(_06687_),
    .A2(_07899_),
    .B1(_07873_),
    .Y(_07944_));
 sky130_fd_sc_hd__nand2_1 _14802_ (.A(_06687_),
    .B(_07870_),
    .Y(_07945_));
 sky130_fd_sc_hd__o211a_1 _14803_ (.A1(_06687_),
    .A2(_07906_),
    .B1(_07945_),
    .C1(_06603_),
    .X(_07946_));
 sky130_fd_sc_hd__o31a_1 _14804_ (.A1(_07877_),
    .A2(_07944_),
    .A3(_07946_),
    .B1(_07862_),
    .X(_07947_));
 sky130_fd_sc_hd__nand2_2 _14805_ (.A(_07943_),
    .B(_07947_),
    .Y(_07948_));
 sky130_fd_sc_hd__buf_4 _14806_ (.A(_07837_),
    .X(_07949_));
 sky130_fd_sc_hd__mux2_1 _14807_ (.A0(\rbzero.wall_tracer.stepDistY[-3] ),
    .A1(_07948_),
    .S(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__clkbuf_1 _14808_ (.A(_07950_),
    .X(_00399_));
 sky130_fd_sc_hd__and3_1 _14809_ (.A(_06603_),
    .B(_07913_),
    .C(_07914_),
    .X(_07951_));
 sky130_fd_sc_hd__o211a_1 _14810_ (.A1(_06548_),
    .A2(_07851_),
    .B1(_07859_),
    .C1(_06612_),
    .X(_07952_));
 sky130_fd_sc_hd__a211o_4 _14811_ (.A1(_07924_),
    .A2(_07951_),
    .B1(_07952_),
    .C1(_06602_),
    .X(_07953_));
 sky130_fd_sc_hd__mux2_1 _14812_ (.A0(\rbzero.wall_tracer.stepDistY[-2] ),
    .A1(_07953_),
    .S(_07949_),
    .X(_07954_));
 sky130_fd_sc_hd__clkbuf_1 _14813_ (.A(_07954_),
    .X(_00400_));
 sky130_fd_sc_hd__or2_1 _14814_ (.A(_07801_),
    .B(_07821_),
    .X(_07955_));
 sky130_fd_sc_hd__a211o_1 _14815_ (.A1(_06555_),
    .A2(_07797_),
    .B1(_07799_),
    .C1(_06566_),
    .X(_07956_));
 sky130_fd_sc_hd__nor2_1 _14816_ (.A(_06644_),
    .B(_07927_),
    .Y(_07957_));
 sky130_fd_sc_hd__a311o_1 _14817_ (.A1(_06644_),
    .A2(_07955_),
    .A3(_07956_),
    .B1(_07957_),
    .C1(_06544_),
    .X(_07958_));
 sky130_fd_sc_hd__a22oi_2 _14818_ (.A1(_06595_),
    .A2(_07868_),
    .B1(_07958_),
    .B2(_06612_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_4 _14819_ (.A(_07863_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__mux2_1 _14820_ (.A0(\rbzero.wall_tracer.stepDistY[-1] ),
    .A1(_07960_),
    .S(_07949_),
    .X(_07961_));
 sky130_fd_sc_hd__clkbuf_1 _14821_ (.A(_07961_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _14822_ (.A0(_07841_),
    .A1(_07850_),
    .S(_06566_),
    .X(_07962_));
 sky130_fd_sc_hd__mux2_1 _14823_ (.A0(_07937_),
    .A1(_07962_),
    .S(_06644_),
    .X(_07963_));
 sky130_fd_sc_hd__nor2_1 _14824_ (.A(_06575_),
    .B(_07895_),
    .Y(_07964_));
 sky130_fd_sc_hd__a31o_1 _14825_ (.A1(_06595_),
    .A2(_06573_),
    .A3(_07891_),
    .B1(_07834_),
    .X(_07965_));
 sky130_fd_sc_hd__a211o_4 _14826_ (.A1(_06612_),
    .A2(_07963_),
    .B1(_07964_),
    .C1(_07965_),
    .X(_07966_));
 sky130_fd_sc_hd__mux2_1 _14827_ (.A0(\rbzero.wall_tracer.stepDistY[0] ),
    .A1(_07966_),
    .S(_07949_),
    .X(_07967_));
 sky130_fd_sc_hd__clkbuf_1 _14828_ (.A(_07967_),
    .X(_00402_));
 sky130_fd_sc_hd__nand2_1 _14829_ (.A(_07802_),
    .B(_07810_),
    .Y(_07968_));
 sky130_fd_sc_hd__nor2_1 _14830_ (.A(_06644_),
    .B(_07822_),
    .Y(_07969_));
 sky130_fd_sc_hd__a21oi_1 _14831_ (.A1(_07811_),
    .A2(_07968_),
    .B1(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__a221o_4 _14832_ (.A1(_06595_),
    .A2(_07900_),
    .B1(_07970_),
    .B2(_06612_),
    .C1(_07834_),
    .X(_07971_));
 sky130_fd_sc_hd__mux2_1 _14833_ (.A0(\rbzero.wall_tracer.stepDistY[1] ),
    .A1(_07971_),
    .S(_07949_),
    .X(_07972_));
 sky130_fd_sc_hd__clkbuf_1 _14834_ (.A(_07972_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _14835_ (.A0(_07842_),
    .A1(_07851_),
    .S(_06549_),
    .X(_07973_));
 sky130_fd_sc_hd__nor2_2 _14836_ (.A(_06461_),
    .B(_07844_),
    .Y(_07974_));
 sky130_fd_sc_hd__a31o_1 _14837_ (.A1(_07811_),
    .A2(_07974_),
    .A3(_07858_),
    .B1(_07834_),
    .X(_07975_));
 sky130_fd_sc_hd__a21o_2 _14838_ (.A1(_06612_),
    .A2(_07973_),
    .B1(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__mux2_1 _14839_ (.A0(\rbzero.wall_tracer.stepDistY[2] ),
    .A1(_07976_),
    .S(_07949_),
    .X(_07977_));
 sky130_fd_sc_hd__clkbuf_1 _14840_ (.A(_07977_),
    .X(_00404_));
 sky130_fd_sc_hd__nand2_1 _14841_ (.A(_06544_),
    .B(_07929_),
    .Y(_07978_));
 sky130_fd_sc_hd__a21oi_1 _14842_ (.A1(_07803_),
    .A2(_07808_),
    .B1(_07809_),
    .Y(_07979_));
 sky130_fd_sc_hd__nor2_1 _14843_ (.A(_07801_),
    .B(_07979_),
    .Y(_07980_));
 sky130_fd_sc_hd__a31o_1 _14844_ (.A1(_06549_),
    .A2(_07955_),
    .A3(_07956_),
    .B1(_06544_),
    .X(_07981_));
 sky130_fd_sc_hd__a21o_1 _14845_ (.A1(_07811_),
    .A2(_07980_),
    .B1(_07981_),
    .X(_07982_));
 sky130_fd_sc_hd__a31o_2 _14846_ (.A1(_06669_),
    .A2(_07978_),
    .A3(_07982_),
    .B1(_07834_),
    .X(_07983_));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(\rbzero.wall_tracer.stepDistY[3] ),
    .A1(_07983_),
    .S(_07949_),
    .X(_07984_));
 sky130_fd_sc_hd__clkbuf_1 _14848_ (.A(_07984_),
    .X(_00405_));
 sky130_fd_sc_hd__a31o_1 _14849_ (.A1(_06687_),
    .A2(_07811_),
    .A3(_07840_),
    .B1(_06544_),
    .X(_07985_));
 sky130_fd_sc_hd__a21oi_1 _14850_ (.A1(_06549_),
    .A2(_07962_),
    .B1(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__nor2_1 _14851_ (.A(_07845_),
    .B(_07938_),
    .Y(_07987_));
 sky130_fd_sc_hd__o31ai_2 _14852_ (.A1(_06461_),
    .A2(_07986_),
    .A3(_07987_),
    .B1(_07863_),
    .Y(_07988_));
 sky130_fd_sc_hd__buf_2 _14853_ (.A(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__mux2_1 _14854_ (.A0(\rbzero.wall_tracer.stepDistY[4] ),
    .A1(_07989_),
    .S(_07949_),
    .X(_07990_));
 sky130_fd_sc_hd__clkbuf_1 _14855_ (.A(_07990_),
    .X(_00406_));
 sky130_fd_sc_hd__or3_1 _14856_ (.A(_06461_),
    .B(_07811_),
    .C(_07968_),
    .X(_07991_));
 sky130_fd_sc_hd__o211ai_4 _14857_ (.A1(_06575_),
    .A2(_07942_),
    .B1(_07991_),
    .C1(_07862_),
    .Y(_07992_));
 sky130_fd_sc_hd__mux2_1 _14858_ (.A0(\rbzero.wall_tracer.stepDistY[5] ),
    .A1(_07992_),
    .S(_07949_),
    .X(_07993_));
 sky130_fd_sc_hd__clkbuf_1 _14859_ (.A(_07993_),
    .X(_00407_));
 sky130_fd_sc_hd__a221o_1 _14860_ (.A1(_06686_),
    .A2(_07842_),
    .B1(_07860_),
    .B2(_07974_),
    .C1(_07834_),
    .X(_07994_));
 sky130_fd_sc_hd__mux2_1 _14861_ (.A0(\rbzero.wall_tracer.stepDistY[6] ),
    .A1(_07994_),
    .S(_07949_),
    .X(_07995_));
 sky130_fd_sc_hd__clkbuf_1 _14862_ (.A(_07995_),
    .X(_00408_));
 sky130_fd_sc_hd__a31o_1 _14863_ (.A1(_07811_),
    .A2(_07955_),
    .A3(_07956_),
    .B1(_07957_),
    .X(_07996_));
 sky130_fd_sc_hd__nor2_1 _14864_ (.A(_07845_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__a21oi_1 _14865_ (.A1(_06686_),
    .A2(_07980_),
    .B1(_07974_),
    .Y(_07998_));
 sky130_fd_sc_hd__o21ai_2 _14866_ (.A1(_07997_),
    .A2(_07998_),
    .B1(_07863_),
    .Y(_07999_));
 sky130_fd_sc_hd__mux2_1 _14867_ (.A0(\rbzero.wall_tracer.stepDistY[7] ),
    .A1(_07999_),
    .S(_07837_),
    .X(_08000_));
 sky130_fd_sc_hd__clkbuf_1 _14868_ (.A(_08000_),
    .X(_00409_));
 sky130_fd_sc_hd__a31o_1 _14869_ (.A1(_06669_),
    .A2(_06573_),
    .A3(_07840_),
    .B1(_07974_),
    .X(_08001_));
 sky130_fd_sc_hd__o21ai_1 _14870_ (.A1(_07845_),
    .A2(_07963_),
    .B1(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__nand2_1 _14871_ (.A(_07863_),
    .B(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__mux2_1 _14872_ (.A0(\rbzero.wall_tracer.stepDistY[8] ),
    .A1(_08003_),
    .S(_07837_),
    .X(_08004_));
 sky130_fd_sc_hd__clkbuf_1 _14873_ (.A(_08004_),
    .X(_00410_));
 sky130_fd_sc_hd__a21o_1 _14874_ (.A1(_07974_),
    .A2(_07970_),
    .B1(_07834_),
    .X(_08005_));
 sky130_fd_sc_hd__mux2_1 _14875_ (.A0(\rbzero.wall_tracer.stepDistY[9] ),
    .A1(_08005_),
    .S(_07837_),
    .X(_08006_));
 sky130_fd_sc_hd__clkbuf_1 _14876_ (.A(_08006_),
    .X(_00411_));
 sky130_fd_sc_hd__and2b_1 _14877_ (.A_N(_06455_),
    .B(_06519_),
    .X(_08007_));
 sky130_fd_sc_hd__and4_1 _14878_ (.A(_07863_),
    .B(_08007_),
    .C(_06544_),
    .D(_07973_),
    .X(_08008_));
 sky130_fd_sc_hd__mux2_1 _14879_ (.A0(\rbzero.wall_tracer.stepDistY[10] ),
    .A1(_08008_),
    .S(_07837_),
    .X(_08009_));
 sky130_fd_sc_hd__clkbuf_1 _14880_ (.A(_08009_),
    .X(_00412_));
 sky130_fd_sc_hd__or2_1 _14881_ (.A(_06101_),
    .B(_06202_),
    .X(_08010_));
 sky130_fd_sc_hd__buf_2 _14882_ (.A(_08010_),
    .X(_08011_));
 sky130_fd_sc_hd__clkbuf_4 _14883_ (.A(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__buf_4 _14884_ (.A(_06251_),
    .X(_08013_));
 sky130_fd_sc_hd__mux2_1 _14885_ (.A0(\rbzero.wall_tracer.trackDistY[-11] ),
    .A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .S(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__clkbuf_4 _14886_ (.A(_06203_),
    .X(_08015_));
 sky130_fd_sc_hd__or2_1 _14887_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__buf_4 _14888_ (.A(_04478_),
    .X(_01622_));
 sky130_fd_sc_hd__o211a_1 _14889_ (.A1(_08012_),
    .A2(_08014_),
    .B1(_08016_),
    .C1(_01622_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _14890_ (.A0(\rbzero.wall_tracer.trackDistY[-10] ),
    .A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .S(_08013_),
    .X(_08017_));
 sky130_fd_sc_hd__inv_2 _14891_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .Y(_08018_));
 sky130_fd_sc_hd__nand2_1 _14892_ (.A(_08018_),
    .B(_08011_),
    .Y(_08019_));
 sky130_fd_sc_hd__o211a_1 _14893_ (.A1(_08012_),
    .A2(_08017_),
    .B1(_08019_),
    .C1(_01622_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _14894_ (.A0(\rbzero.wall_tracer.trackDistY[-9] ),
    .A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .S(_08013_),
    .X(_08020_));
 sky130_fd_sc_hd__or2_1 _14895_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(_08015_),
    .X(_08021_));
 sky130_fd_sc_hd__o211a_1 _14896_ (.A1(_08012_),
    .A2(_08020_),
    .B1(_08021_),
    .C1(_01622_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _14897_ (.A0(\rbzero.wall_tracer.trackDistY[-8] ),
    .A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .S(_08013_),
    .X(_08022_));
 sky130_fd_sc_hd__or2_1 _14898_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_08015_),
    .X(_08023_));
 sky130_fd_sc_hd__o211a_1 _14899_ (.A1(_08012_),
    .A2(_08022_),
    .B1(_08023_),
    .C1(_01622_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _14900_ (.A0(\rbzero.wall_tracer.trackDistY[-7] ),
    .A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .S(_08013_),
    .X(_08024_));
 sky130_fd_sc_hd__or2_1 _14901_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(_08015_),
    .X(_08025_));
 sky130_fd_sc_hd__o211a_1 _14902_ (.A1(_08012_),
    .A2(_08024_),
    .B1(_08025_),
    .C1(_01622_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _14903_ (.A0(\rbzero.wall_tracer.trackDistY[-6] ),
    .A1(\rbzero.wall_tracer.trackDistX[-6] ),
    .S(_08013_),
    .X(_08026_));
 sky130_fd_sc_hd__or2_1 _14904_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(_08015_),
    .X(_08027_));
 sky130_fd_sc_hd__o211a_1 _14905_ (.A1(_08012_),
    .A2(_08026_),
    .B1(_08027_),
    .C1(_01622_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _14906_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .S(_08013_),
    .X(_08028_));
 sky130_fd_sc_hd__or2_1 _14907_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_08015_),
    .X(_08029_));
 sky130_fd_sc_hd__o211a_1 _14908_ (.A1(_08012_),
    .A2(_08028_),
    .B1(_08029_),
    .C1(_01622_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _14909_ (.A0(\rbzero.wall_tracer.trackDistY[-4] ),
    .A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .S(_08013_),
    .X(_08030_));
 sky130_fd_sc_hd__or2_1 _14910_ (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .B(_08015_),
    .X(_08031_));
 sky130_fd_sc_hd__o211a_1 _14911_ (.A1(_08012_),
    .A2(_08030_),
    .B1(_08031_),
    .C1(_01622_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _14912_ (.A0(\rbzero.wall_tracer.trackDistY[-3] ),
    .A1(\rbzero.wall_tracer.trackDistX[-3] ),
    .S(_08013_),
    .X(_08032_));
 sky130_fd_sc_hd__clkbuf_2 _14913_ (.A(_06203_),
    .X(_08033_));
 sky130_fd_sc_hd__or2_1 _14914_ (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .B(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__buf_2 _14915_ (.A(_04478_),
    .X(_08035_));
 sky130_fd_sc_hd__o211a_1 _14916_ (.A1(_08012_),
    .A2(_08032_),
    .B1(_08034_),
    .C1(_08035_),
    .X(_00421_));
 sky130_fd_sc_hd__clkbuf_4 _14917_ (.A(_06251_),
    .X(_08036_));
 sky130_fd_sc_hd__mux2_1 _14918_ (.A0(\rbzero.wall_tracer.trackDistY[-2] ),
    .A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .S(_08036_),
    .X(_08037_));
 sky130_fd_sc_hd__or2_1 _14919_ (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .B(_08033_),
    .X(_08038_));
 sky130_fd_sc_hd__o211a_1 _14920_ (.A1(_08012_),
    .A2(_08037_),
    .B1(_08038_),
    .C1(_08035_),
    .X(_00422_));
 sky130_fd_sc_hd__buf_2 _14921_ (.A(_08011_),
    .X(_08039_));
 sky130_fd_sc_hd__mux2_1 _14922_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .S(_08036_),
    .X(_08040_));
 sky130_fd_sc_hd__or2_1 _14923_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(_08033_),
    .X(_08041_));
 sky130_fd_sc_hd__o211a_1 _14924_ (.A1(_08039_),
    .A2(_08040_),
    .B1(_08041_),
    .C1(_08035_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _14925_ (.A0(\rbzero.wall_tracer.trackDistY[0] ),
    .A1(\rbzero.wall_tracer.trackDistX[0] ),
    .S(_08036_),
    .X(_08042_));
 sky130_fd_sc_hd__inv_2 _14926_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .Y(_08043_));
 sky130_fd_sc_hd__nand2_1 _14927_ (.A(_08043_),
    .B(_08011_),
    .Y(_08044_));
 sky130_fd_sc_hd__o211a_1 _14928_ (.A1(_08039_),
    .A2(_08042_),
    .B1(_08044_),
    .C1(_08035_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _14929_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(\rbzero.wall_tracer.trackDistX[1] ),
    .S(_08036_),
    .X(_08045_));
 sky130_fd_sc_hd__or2_1 _14930_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08033_),
    .X(_08046_));
 sky130_fd_sc_hd__o211a_1 _14931_ (.A1(_08039_),
    .A2(_08045_),
    .B1(_08046_),
    .C1(_08035_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _14932_ (.A0(\rbzero.wall_tracer.trackDistY[2] ),
    .A1(\rbzero.wall_tracer.trackDistX[2] ),
    .S(_08036_),
    .X(_08047_));
 sky130_fd_sc_hd__or2_1 _14933_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08033_),
    .X(_08048_));
 sky130_fd_sc_hd__o211a_1 _14934_ (.A1(_08039_),
    .A2(_08047_),
    .B1(_08048_),
    .C1(_08035_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _14935_ (.A0(\rbzero.wall_tracer.trackDistY[3] ),
    .A1(\rbzero.wall_tracer.trackDistX[3] ),
    .S(_08036_),
    .X(_08049_));
 sky130_fd_sc_hd__or2_1 _14936_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08033_),
    .X(_08050_));
 sky130_fd_sc_hd__o211a_1 _14937_ (.A1(_08039_),
    .A2(_08049_),
    .B1(_08050_),
    .C1(_08035_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _14938_ (.A0(\rbzero.wall_tracer.trackDistY[4] ),
    .A1(\rbzero.wall_tracer.trackDistX[4] ),
    .S(_08036_),
    .X(_08051_));
 sky130_fd_sc_hd__or2_1 _14939_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08033_),
    .X(_08052_));
 sky130_fd_sc_hd__o211a_1 _14940_ (.A1(_08039_),
    .A2(_08051_),
    .B1(_08052_),
    .C1(_08035_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _14941_ (.A0(\rbzero.wall_tracer.trackDistY[5] ),
    .A1(\rbzero.wall_tracer.trackDistX[5] ),
    .S(_08036_),
    .X(_08053_));
 sky130_fd_sc_hd__or2_1 _14942_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08033_),
    .X(_08054_));
 sky130_fd_sc_hd__o211a_1 _14943_ (.A1(_08039_),
    .A2(_08053_),
    .B1(_08054_),
    .C1(_08035_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _14944_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(\rbzero.wall_tracer.trackDistX[6] ),
    .S(_08036_),
    .X(_08055_));
 sky130_fd_sc_hd__or2_1 _14945_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08033_),
    .X(_08056_));
 sky130_fd_sc_hd__o211a_1 _14946_ (.A1(_08039_),
    .A2(_08055_),
    .B1(_08056_),
    .C1(_08035_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _14947_ (.A0(\rbzero.wall_tracer.trackDistY[7] ),
    .A1(\rbzero.wall_tracer.trackDistX[7] ),
    .S(_08036_),
    .X(_08057_));
 sky130_fd_sc_hd__or2_1 _14948_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08033_),
    .X(_08058_));
 sky130_fd_sc_hd__buf_4 _14949_ (.A(_04478_),
    .X(_08059_));
 sky130_fd_sc_hd__o211a_1 _14950_ (.A1(_08039_),
    .A2(_08057_),
    .B1(_08058_),
    .C1(_08059_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(\rbzero.wall_tracer.trackDistY[8] ),
    .A1(\rbzero.wall_tracer.trackDistX[8] ),
    .S(_06251_),
    .X(_08060_));
 sky130_fd_sc_hd__or2_1 _14952_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_06203_),
    .X(_08061_));
 sky130_fd_sc_hd__o211a_1 _14953_ (.A1(_08039_),
    .A2(_08060_),
    .B1(_08061_),
    .C1(_08059_),
    .X(_00432_));
 sky130_fd_sc_hd__a211oi_1 _14954_ (.A1(_06204_),
    .A2(\rbzero.wall_tracer.trackDistY[10] ),
    .B1(_06205_),
    .C1(_06250_),
    .Y(_08062_));
 sky130_fd_sc_hd__a211o_1 _14955_ (.A1(\rbzero.wall_tracer.trackDistX[9] ),
    .A2(_08013_),
    .B1(_08062_),
    .C1(_08011_),
    .X(_08063_));
 sky130_fd_sc_hd__o211a_1 _14956_ (.A1(\rbzero.wall_tracer.visualWallDist[9] ),
    .A2(_08015_),
    .B1(_08063_),
    .C1(_08059_),
    .X(_00433_));
 sky130_fd_sc_hd__a21o_1 _14957_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(\rbzero.wall_tracer.trackDistY[10] ),
    .B1(_08011_),
    .X(_08064_));
 sky130_fd_sc_hd__o211a_1 _14958_ (.A1(\rbzero.wall_tracer.visualWallDist[10] ),
    .A2(_08015_),
    .B1(_08064_),
    .C1(_08059_),
    .X(_00434_));
 sky130_fd_sc_hd__and4b_1 _14959_ (.A_N(_04471_),
    .B(_04469_),
    .C(_04475_),
    .D(_04472_),
    .X(_08065_));
 sky130_fd_sc_hd__clkbuf_4 _14960_ (.A(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__clkbuf_4 _14961_ (.A(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(\rbzero.wall_tracer.stepDistX[-11] ),
    .A1(_07835_),
    .S(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__clkbuf_1 _14963_ (.A(_08068_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _14964_ (.A0(\rbzero.wall_tracer.stepDistX[-10] ),
    .A1(_07864_),
    .S(_08067_),
    .X(_08069_));
 sky130_fd_sc_hd__clkbuf_1 _14965_ (.A(_08069_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _14966_ (.A0(\rbzero.wall_tracer.stepDistX[-9] ),
    .A1(_07880_),
    .S(_08067_),
    .X(_08070_));
 sky130_fd_sc_hd__clkbuf_1 _14967_ (.A(_08070_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _14968_ (.A0(\rbzero.wall_tracer.stepDistX[-8] ),
    .A1(_07897_),
    .S(_08067_),
    .X(_08071_));
 sky130_fd_sc_hd__clkbuf_1 _14969_ (.A(_08071_),
    .X(_00438_));
 sky130_fd_sc_hd__nor2_1 _14970_ (.A(\rbzero.wall_tracer.stepDistX[-7] ),
    .B(_08067_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21oi_1 _14971_ (.A1(_07911_),
    .A2(_08067_),
    .B1(_08072_),
    .Y(_00439_));
 sky130_fd_sc_hd__mux2_1 _14972_ (.A0(\rbzero.wall_tracer.stepDistX[-6] ),
    .A1(_07920_),
    .S(_08067_),
    .X(_08073_));
 sky130_fd_sc_hd__clkbuf_1 _14973_ (.A(_08073_),
    .X(_00440_));
 sky130_fd_sc_hd__nor2_1 _14974_ (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(_08067_),
    .Y(_08074_));
 sky130_fd_sc_hd__a21oi_1 _14975_ (.A1(_07931_),
    .A2(_08067_),
    .B1(_08074_),
    .Y(_00441_));
 sky130_fd_sc_hd__mux2_1 _14976_ (.A0(\rbzero.wall_tracer.stepDistX[-4] ),
    .A1(_07940_),
    .S(_08067_),
    .X(_08075_));
 sky130_fd_sc_hd__clkbuf_1 _14977_ (.A(_08075_),
    .X(_00442_));
 sky130_fd_sc_hd__buf_4 _14978_ (.A(_08066_),
    .X(_08076_));
 sky130_fd_sc_hd__mux2_1 _14979_ (.A0(\rbzero.wall_tracer.stepDistX[-3] ),
    .A1(_07948_),
    .S(_08076_),
    .X(_08077_));
 sky130_fd_sc_hd__clkbuf_1 _14980_ (.A(_08077_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _14981_ (.A0(\rbzero.wall_tracer.stepDistX[-2] ),
    .A1(_07953_),
    .S(_08076_),
    .X(_08078_));
 sky130_fd_sc_hd__clkbuf_1 _14982_ (.A(_08078_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _14983_ (.A0(\rbzero.wall_tracer.stepDistX[-1] ),
    .A1(_07960_),
    .S(_08076_),
    .X(_08079_));
 sky130_fd_sc_hd__clkbuf_1 _14984_ (.A(_08079_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _14985_ (.A0(\rbzero.wall_tracer.stepDistX[0] ),
    .A1(_07966_),
    .S(_08076_),
    .X(_08080_));
 sky130_fd_sc_hd__clkbuf_1 _14986_ (.A(_08080_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _14987_ (.A0(\rbzero.wall_tracer.stepDistX[1] ),
    .A1(_07971_),
    .S(_08076_),
    .X(_08081_));
 sky130_fd_sc_hd__clkbuf_1 _14988_ (.A(_08081_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _14989_ (.A0(\rbzero.wall_tracer.stepDistX[2] ),
    .A1(_07976_),
    .S(_08076_),
    .X(_08082_));
 sky130_fd_sc_hd__clkbuf_1 _14990_ (.A(_08082_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _14991_ (.A0(\rbzero.wall_tracer.stepDistX[3] ),
    .A1(_07983_),
    .S(_08076_),
    .X(_08083_));
 sky130_fd_sc_hd__clkbuf_1 _14992_ (.A(_08083_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14993_ (.A0(\rbzero.wall_tracer.stepDistX[4] ),
    .A1(_07989_),
    .S(_08076_),
    .X(_08084_));
 sky130_fd_sc_hd__clkbuf_1 _14994_ (.A(_08084_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _14995_ (.A0(\rbzero.wall_tracer.stepDistX[5] ),
    .A1(_07992_),
    .S(_08076_),
    .X(_08085_));
 sky130_fd_sc_hd__clkbuf_1 _14996_ (.A(_08085_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _14997_ (.A0(\rbzero.wall_tracer.stepDistX[6] ),
    .A1(_07994_),
    .S(_08076_),
    .X(_08086_));
 sky130_fd_sc_hd__clkbuf_1 _14998_ (.A(_08086_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _14999_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_07999_),
    .S(_08066_),
    .X(_08087_));
 sky130_fd_sc_hd__clkbuf_1 _15000_ (.A(_08087_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _15001_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_08003_),
    .S(_08066_),
    .X(_08088_));
 sky130_fd_sc_hd__clkbuf_1 _15002_ (.A(_08088_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _15003_ (.A0(\rbzero.wall_tracer.stepDistX[9] ),
    .A1(_08005_),
    .S(_08066_),
    .X(_08089_));
 sky130_fd_sc_hd__clkbuf_1 _15004_ (.A(_08089_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _15005_ (.A0(\rbzero.wall_tracer.stepDistX[10] ),
    .A1(_08008_),
    .S(_08066_),
    .X(_08090_));
 sky130_fd_sc_hd__clkbuf_1 _15006_ (.A(_08090_),
    .X(_00456_));
 sky130_fd_sc_hd__buf_4 _15007_ (.A(_04015_),
    .X(_08091_));
 sky130_fd_sc_hd__clkbuf_8 _15008_ (.A(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__buf_4 _15009_ (.A(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__and2_1 _15010_ (.A(_08093_),
    .B(_05081_),
    .X(_08094_));
 sky130_fd_sc_hd__clkbuf_1 _15011_ (.A(_08094_),
    .X(_00457_));
 sky130_fd_sc_hd__nor2_1 _15012_ (.A(net65),
    .B(_05316_),
    .Y(_00458_));
 sky130_fd_sc_hd__and2_1 _15013_ (.A(_08093_),
    .B(_05399_),
    .X(_08095_));
 sky130_fd_sc_hd__clkbuf_1 _15014_ (.A(_08095_),
    .X(_00459_));
 sky130_fd_sc_hd__and2_1 _15015_ (.A(_08093_),
    .B(_05492_),
    .X(_08096_));
 sky130_fd_sc_hd__clkbuf_1 _15016_ (.A(_08096_),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _15017_ (.A(_08093_),
    .B(_05582_),
    .X(_08097_));
 sky130_fd_sc_hd__clkbuf_1 _15018_ (.A(_08097_),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _15019_ (.A(_08093_),
    .B(_05671_),
    .X(_08098_));
 sky130_fd_sc_hd__clkbuf_1 _15020_ (.A(_08098_),
    .X(_00462_));
 sky130_fd_sc_hd__nor2_4 _15021_ (.A(_04465_),
    .B(_04473_),
    .Y(_08099_));
 sky130_fd_sc_hd__buf_6 _15022_ (.A(_08099_),
    .X(_08100_));
 sky130_fd_sc_hd__buf_8 _15023_ (.A(_08100_),
    .X(_08101_));
 sky130_fd_sc_hd__nand2_1 _15024_ (.A(_08101_),
    .B(_06202_),
    .Y(_08102_));
 sky130_fd_sc_hd__or2_1 _15025_ (.A(_06137_),
    .B(_06200_),
    .X(_08103_));
 sky130_fd_sc_hd__or3b_1 _15026_ (.A(_06145_),
    .B(_06180_),
    .C_N(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__a21bo_1 _15027_ (.A1(\rbzero.mapdyw[0] ),
    .A2(_06145_),
    .B1_N(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__mux2_1 _15028_ (.A0(_08105_),
    .A1(\rbzero.mapdxw[0] ),
    .S(_06154_),
    .X(_08106_));
 sky130_fd_sc_hd__a21o_1 _15029_ (.A1(_08101_),
    .A2(_06202_),
    .B1(\rbzero.wall_hot[0] ),
    .X(_08107_));
 sky130_fd_sc_hd__o211a_1 _15030_ (.A1(_08102_),
    .A2(_08106_),
    .B1(_08107_),
    .C1(_08059_),
    .X(_00463_));
 sky130_fd_sc_hd__nor2_1 _15031_ (.A(_06145_),
    .B(_06187_),
    .Y(_08108_));
 sky130_fd_sc_hd__a22o_1 _15032_ (.A1(\rbzero.mapdyw[1] ),
    .A2(_06145_),
    .B1(_08103_),
    .B2(_08108_),
    .X(_08109_));
 sky130_fd_sc_hd__mux2_1 _15033_ (.A0(_08109_),
    .A1(\rbzero.mapdxw[1] ),
    .S(_06154_),
    .X(_08110_));
 sky130_fd_sc_hd__buf_6 _15034_ (.A(_04467_),
    .X(_08111_));
 sky130_fd_sc_hd__clkbuf_4 _15035_ (.A(_08111_),
    .X(_08112_));
 sky130_fd_sc_hd__buf_6 _15036_ (.A(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__a21oi_1 _15037_ (.A1(_04494_),
    .A2(_08102_),
    .B1(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__o21a_1 _15038_ (.A1(_08102_),
    .A2(_08110_),
    .B1(_08114_),
    .X(_00464_));
 sky130_fd_sc_hd__buf_4 _15039_ (.A(_04511_),
    .X(_08115_));
 sky130_fd_sc_hd__o211a_1 _15040_ (.A1(_08115_),
    .A2(_08015_),
    .B1(_06252_),
    .C1(_08059_),
    .X(_00465_));
 sky130_fd_sc_hd__nand2_1 _15041_ (.A(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .Y(_08116_));
 sky130_fd_sc_hd__nor2_1 _15042_ (.A(_04465_),
    .B(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__buf_2 _15043_ (.A(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__buf_4 _15044_ (.A(_08118_),
    .X(_08119_));
 sky130_fd_sc_hd__buf_4 _15045_ (.A(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__and2b_1 _15046_ (.A_N(_04511_),
    .B(\rbzero.debug_overlay.playerY[-6] ),
    .X(_08121_));
 sky130_fd_sc_hd__a21oi_1 _15047_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_08115_),
    .B1(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__buf_4 _15048_ (.A(_06158_),
    .X(_08123_));
 sky130_fd_sc_hd__buf_6 _15049_ (.A(_08123_),
    .X(_08124_));
 sky130_fd_sc_hd__nand2_4 _15050_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__buf_2 _15051_ (.A(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__buf_4 _15052_ (.A(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__or2_1 _15053_ (.A(\rbzero.trace_state[0] ),
    .B(_06158_),
    .X(_08128_));
 sky130_fd_sc_hd__clkbuf_8 _15054_ (.A(_08128_),
    .X(_08129_));
 sky130_fd_sc_hd__buf_8 _15055_ (.A(_08129_),
    .X(_08130_));
 sky130_fd_sc_hd__or2_1 _15056_ (.A(_04465_),
    .B(_08116_),
    .X(_08131_));
 sky130_fd_sc_hd__buf_4 _15057_ (.A(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__mux2_1 _15058_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(_04510_),
    .X(_08133_));
 sky130_fd_sc_hd__and3_1 _15059_ (.A(_04472_),
    .B(\rbzero.trace_state[0] ),
    .C(_06157_),
    .X(_08134_));
 sky130_fd_sc_hd__buf_4 _15060_ (.A(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__a21o_1 _15061_ (.A1(_08119_),
    .A2(_08133_),
    .B1(_08135_),
    .X(_08136_));
 sky130_fd_sc_hd__a21o_2 _15062_ (.A1(_07835_),
    .A2(_08132_),
    .B1(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__o211ai_4 _15063_ (.A1(\rbzero.wall_tracer.stepDistY[-11] ),
    .A2(_08124_),
    .B1(_08130_),
    .C1(_08137_),
    .Y(_08138_));
 sky130_fd_sc_hd__mux2_1 _15064_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(_04510_),
    .X(_08139_));
 sky130_fd_sc_hd__or2_1 _15065_ (.A(_08132_),
    .B(_08139_),
    .X(_08140_));
 sky130_fd_sc_hd__and2_1 _15066_ (.A(\rbzero.trace_state[1] ),
    .B(_06157_),
    .X(_08141_));
 sky130_fd_sc_hd__buf_4 _15067_ (.A(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__nand2_4 _15068_ (.A(\rbzero.trace_state[0] ),
    .B(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__buf_6 _15069_ (.A(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__o211a_4 _15070_ (.A1(_07864_),
    .A2(_08119_),
    .B1(_08140_),
    .C1(_08144_),
    .X(_08145_));
 sky130_fd_sc_hd__a21o_2 _15071_ (.A1(\rbzero.wall_tracer.stepDistY[-10] ),
    .A2(_08142_),
    .B1(_06160_),
    .X(_08146_));
 sky130_fd_sc_hd__nor2_4 _15072_ (.A(_08145_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__nand2_8 _15073_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08124_),
    .Y(_08148_));
 sky130_fd_sc_hd__or2_1 _15074_ (.A(_08147_),
    .B(_08148_),
    .X(_08149_));
 sky130_fd_sc_hd__or3_2 _15075_ (.A(_08127_),
    .B(_08138_),
    .C(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__a21o_1 _15076_ (.A1(_07943_),
    .A2(_07947_),
    .B1(_08117_),
    .X(_08151_));
 sky130_fd_sc_hd__nand2_1 _15077_ (.A(\rbzero.side_hot ),
    .B(_06345_),
    .Y(_08152_));
 sky130_fd_sc_hd__o211a_1 _15078_ (.A1(_04509_),
    .A2(_06048_),
    .B1(_08117_),
    .C1(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__nor2_1 _15079_ (.A(_08142_),
    .B(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__a2bb2o_1 _15080_ (.A1_N(\rbzero.wall_tracer.stepDistY[-3] ),
    .A2_N(_08143_),
    .B1(_08151_),
    .B2(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__o21bai_4 _15081_ (.A1(\rbzero.wall_tracer.stepDistX[-3] ),
    .A2(_08129_),
    .B1_N(_08155_),
    .Y(_08156_));
 sky130_fd_sc_hd__xor2_1 _15082_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(\rbzero.debug_overlay.playerY[-9] ),
    .X(_08157_));
 sky130_fd_sc_hd__mux2_1 _15083_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(_08157_),
    .S(_06074_),
    .X(_08158_));
 sky130_fd_sc_hd__mux2_1 _15084_ (.A0(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A1(_08158_),
    .S(_08134_),
    .X(_08159_));
 sky130_fd_sc_hd__nor2_1 _15085_ (.A(_06390_),
    .B(_06391_),
    .Y(_08160_));
 sky130_fd_sc_hd__or3b_1 _15086_ (.A(\rbzero.wall_tracer.rayAddendX[-2] ),
    .B(_06376_),
    .C_N(_06366_),
    .X(_08161_));
 sky130_fd_sc_hd__or4_1 _15087_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .B(_06381_),
    .C(_06360_),
    .D(_08161_),
    .X(_08162_));
 sky130_fd_sc_hd__nand4_1 _15088_ (.A(_06341_),
    .B(_06345_),
    .C(_06350_),
    .D(_06354_),
    .Y(_08163_));
 sky130_fd_sc_hd__or4b_1 _15089_ (.A(_08160_),
    .B(_08162_),
    .C(_08163_),
    .D_N(_06396_),
    .X(_08164_));
 sky130_fd_sc_hd__nor2_1 _15090_ (.A(_06331_),
    .B(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__a21bo_2 _15091_ (.A1(_06327_),
    .A2(_08165_),
    .B1_N(_06413_),
    .X(_08166_));
 sky130_fd_sc_hd__xnor2_2 _15092_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_08167_));
 sky130_fd_sc_hd__or2_1 _15093_ (.A(_08166_),
    .B(_08167_),
    .X(_08168_));
 sky130_fd_sc_hd__a21oi_1 _15094_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(_08166_),
    .B1(_08128_),
    .Y(_08169_));
 sky130_fd_sc_hd__a2bb2o_2 _15095_ (.A1_N(_06159_),
    .A2_N(_08159_),
    .B1(_08168_),
    .B2(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__buf_4 _15096_ (.A(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__a21o_1 _15097_ (.A1(_07935_),
    .A2(_07939_),
    .B1(_08118_),
    .X(_08172_));
 sky130_fd_sc_hd__nand2_1 _15098_ (.A(_04509_),
    .B(_06350_),
    .Y(_08173_));
 sky130_fd_sc_hd__o211a_1 _15099_ (.A1(_04509_),
    .A2(_06052_),
    .B1(_08118_),
    .C1(_08173_),
    .X(_08174_));
 sky130_fd_sc_hd__nor2_1 _15100_ (.A(_08142_),
    .B(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__a2bb2o_4 _15101_ (.A1_N(\rbzero.wall_tracer.stepDistY[-4] ),
    .A2_N(_08144_),
    .B1(_08172_),
    .B2(_08175_),
    .X(_08176_));
 sky130_fd_sc_hd__o21bai_4 _15102_ (.A1(\rbzero.wall_tracer.stepDistX[-4] ),
    .A2(_08129_),
    .B1_N(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__buf_4 _15103_ (.A(_08166_),
    .X(_08178_));
 sky130_fd_sc_hd__or3_1 _15104_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(\rbzero.debug_overlay.playerX[-8] ),
    .C(\rbzero.debug_overlay.playerX[-9] ),
    .X(_08179_));
 sky130_fd_sc_hd__o21ai_1 _15105_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(\rbzero.debug_overlay.playerX[-9] ),
    .B1(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_08180_));
 sky130_fd_sc_hd__nand2_1 _15106_ (.A(_08179_),
    .B(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__nor2_1 _15107_ (.A(_08178_),
    .B(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__a21o_1 _15108_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_08166_),
    .B1(_08128_),
    .X(_08183_));
 sky130_fd_sc_hd__or3_1 _15109_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(\rbzero.debug_overlay.playerY[-8] ),
    .C(\rbzero.debug_overlay.playerY[-9] ),
    .X(_08184_));
 sky130_fd_sc_hd__o21ai_1 _15110_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(\rbzero.debug_overlay.playerY[-9] ),
    .B1(\rbzero.debug_overlay.playerY[-7] ),
    .Y(_08185_));
 sky130_fd_sc_hd__nand2_1 _15111_ (.A(_08184_),
    .B(_08185_),
    .Y(_08186_));
 sky130_fd_sc_hd__nand2_1 _15112_ (.A(_06074_),
    .B(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__o211a_1 _15113_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_06074_),
    .B1(_08134_),
    .C1(_08187_),
    .X(_08188_));
 sky130_fd_sc_hd__a211o_1 _15114_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_08143_),
    .B1(_08188_),
    .C1(_06160_),
    .X(_08189_));
 sky130_fd_sc_hd__o21ai_4 _15115_ (.A1(_08182_),
    .A2(_08183_),
    .B1(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__clkbuf_4 _15116_ (.A(_08190_),
    .X(_08191_));
 sky130_fd_sc_hd__o22ai_1 _15117_ (.A1(_08156_),
    .A2(_08171_),
    .B1(_08177_),
    .B2(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__or2_1 _15118_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08184_),
    .X(_08193_));
 sky130_fd_sc_hd__nand2_1 _15119_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08184_),
    .Y(_08194_));
 sky130_fd_sc_hd__nand2_1 _15120_ (.A(_08193_),
    .B(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__nor2_1 _15121_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_06075_),
    .Y(_08196_));
 sky130_fd_sc_hd__a211o_1 _15122_ (.A1(_06075_),
    .A2(_08195_),
    .B1(_08196_),
    .C1(_08144_),
    .X(_08197_));
 sky130_fd_sc_hd__a21oi_1 _15123_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_08123_),
    .B1(_06160_),
    .Y(_08198_));
 sky130_fd_sc_hd__or2_1 _15124_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08179_),
    .X(_08199_));
 sky130_fd_sc_hd__nand2_1 _15125_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08179_),
    .Y(_08200_));
 sky130_fd_sc_hd__nand2_1 _15126_ (.A(_08199_),
    .B(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__clkinv_2 _15127_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .Y(_08202_));
 sky130_fd_sc_hd__mux2_1 _15128_ (.A0(_08201_),
    .A1(_08202_),
    .S(_08178_),
    .X(_08203_));
 sky130_fd_sc_hd__a22o_4 _15129_ (.A1(_08197_),
    .A2(_08198_),
    .B1(_08203_),
    .B2(_06161_),
    .X(_08204_));
 sky130_fd_sc_hd__nor2_1 _15130_ (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(_08129_),
    .Y(_08205_));
 sky130_fd_sc_hd__nor2_1 _15131_ (.A(_04509_),
    .B(_06054_),
    .Y(_08206_));
 sky130_fd_sc_hd__a211o_1 _15132_ (.A1(_04509_),
    .A2(_06354_),
    .B1(_08132_),
    .C1(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__o21a_1 _15133_ (.A1(_07931_),
    .A2(_08118_),
    .B1(_08207_),
    .X(_08208_));
 sky130_fd_sc_hd__a2bb2o_4 _15134_ (.A1_N(\rbzero.wall_tracer.stepDistY[-5] ),
    .A2_N(_08143_),
    .B1(_08208_),
    .B2(_06158_),
    .X(_08209_));
 sky130_fd_sc_hd__or2_1 _15135_ (.A(_08205_),
    .B(_08209_),
    .X(_08210_));
 sky130_fd_sc_hd__buf_2 _15136_ (.A(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__nor2_1 _15137_ (.A(_08204_),
    .B(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__or4_1 _15138_ (.A(_08156_),
    .B(_08191_),
    .C(_08171_),
    .D(_08177_),
    .X(_08213_));
 sky130_fd_sc_hd__a21bo_1 _15139_ (.A1(_08192_),
    .A2(_08212_),
    .B1_N(_08213_),
    .X(_08214_));
 sky130_fd_sc_hd__xnor2_1 _15140_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_08193_),
    .Y(_08215_));
 sky130_fd_sc_hd__nor2_1 _15141_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_06074_),
    .Y(_08216_));
 sky130_fd_sc_hd__a211o_1 _15142_ (.A1(_06074_),
    .A2(_08215_),
    .B1(_08216_),
    .C1(_08143_),
    .X(_08217_));
 sky130_fd_sc_hd__a21oi_1 _15143_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_08123_),
    .B1(_06160_),
    .Y(_08218_));
 sky130_fd_sc_hd__xnor2_2 _15144_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_08199_),
    .Y(_08219_));
 sky130_fd_sc_hd__inv_2 _15145_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .Y(_08220_));
 sky130_fd_sc_hd__mux2_1 _15146_ (.A0(_08219_),
    .A1(_08220_),
    .S(_08166_),
    .X(_08221_));
 sky130_fd_sc_hd__a22o_2 _15147_ (.A1(_08217_),
    .A2(_08218_),
    .B1(_08221_),
    .B2(_06160_),
    .X(_08222_));
 sky130_fd_sc_hd__buf_2 _15148_ (.A(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__nor2_1 _15149_ (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .B(_08129_),
    .Y(_08224_));
 sky130_fd_sc_hd__a21o_1 _15150_ (.A1(_07863_),
    .A2(_07919_),
    .B1(_08118_),
    .X(_08225_));
 sky130_fd_sc_hd__mux2_1 _15151_ (.A0(_06058_),
    .A1(_06360_),
    .S(_04509_),
    .X(_08226_));
 sky130_fd_sc_hd__a21oi_1 _15152_ (.A1(_08118_),
    .A2(_08226_),
    .B1(_08142_),
    .Y(_08227_));
 sky130_fd_sc_hd__a2bb2o_2 _15153_ (.A1_N(\rbzero.wall_tracer.stepDistY[-6] ),
    .A2_N(_08143_),
    .B1(_08225_),
    .B2(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__or2_1 _15154_ (.A(_08224_),
    .B(_08228_),
    .X(_08229_));
 sky130_fd_sc_hd__buf_2 _15155_ (.A(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__or3_1 _15156_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .C(_08193_),
    .X(_08231_));
 sky130_fd_sc_hd__o21ai_1 _15157_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_08193_),
    .B1(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_08232_));
 sky130_fd_sc_hd__nand2_1 _15158_ (.A(_08231_),
    .B(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand2_1 _15159_ (.A(_06074_),
    .B(_08233_),
    .Y(_08234_));
 sky130_fd_sc_hd__o211a_1 _15160_ (.A1(\rbzero.debug_overlay.playerY[-4] ),
    .A2(_06074_),
    .B1(_08134_),
    .C1(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__a21oi_1 _15161_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_08143_),
    .B1(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__or3_1 _15162_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(\rbzero.debug_overlay.playerX[-5] ),
    .C(_08199_),
    .X(_08237_));
 sky130_fd_sc_hd__o21ai_1 _15163_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_08199_),
    .B1(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_08238_));
 sky130_fd_sc_hd__nand2_1 _15164_ (.A(_08237_),
    .B(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__or2_1 _15165_ (.A(_08166_),
    .B(_08239_),
    .X(_08240_));
 sky130_fd_sc_hd__a21oi_1 _15166_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_08166_),
    .B1(_08129_),
    .Y(_08241_));
 sky130_fd_sc_hd__a22o_4 _15167_ (.A1(_08129_),
    .A2(_08236_),
    .B1(_08240_),
    .B2(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__clkbuf_4 _15168_ (.A(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__or4_1 _15169_ (.A(_08211_),
    .B(_08223_),
    .C(_08230_),
    .D(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__clkbuf_4 _15170_ (.A(_08228_),
    .X(_08245_));
 sky130_fd_sc_hd__nor2_1 _15171_ (.A(_08224_),
    .B(_08245_),
    .Y(_08246_));
 sky130_fd_sc_hd__clkinv_4 _15172_ (.A(_08242_),
    .Y(_08247_));
 sky130_fd_sc_hd__a2bb2o_1 _15173_ (.A1_N(_08211_),
    .A2_N(_08223_),
    .B1(_08246_),
    .B2(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__nand2_1 _15174_ (.A(_08244_),
    .B(_08248_),
    .Y(_08249_));
 sky130_fd_sc_hd__or2_2 _15175_ (.A(\rbzero.wall_tracer.stepDistX[-7] ),
    .B(_08129_),
    .X(_08250_));
 sky130_fd_sc_hd__nor2_1 _15176_ (.A(_04510_),
    .B(_06060_),
    .Y(_08251_));
 sky130_fd_sc_hd__a211o_1 _15177_ (.A1(_04510_),
    .A2(_06366_),
    .B1(_08132_),
    .C1(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__o211ai_4 _15178_ (.A1(_07911_),
    .A2(_08119_),
    .B1(_08252_),
    .C1(_08123_),
    .Y(_08253_));
 sky130_fd_sc_hd__o211ai_4 _15179_ (.A1(\rbzero.wall_tracer.stepDistY[-7] ),
    .A2(_08144_),
    .B1(_08250_),
    .C1(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__clkbuf_4 _15180_ (.A(_08254_),
    .X(_08255_));
 sky130_fd_sc_hd__or2_1 _15181_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08231_),
    .X(_08256_));
 sky130_fd_sc_hd__nand2_1 _15182_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08231_),
    .Y(_08257_));
 sky130_fd_sc_hd__nand2_1 _15183_ (.A(_08256_),
    .B(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__nor2_1 _15184_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_06075_),
    .Y(_08259_));
 sky130_fd_sc_hd__a211o_1 _15185_ (.A1(_06075_),
    .A2(_08258_),
    .B1(_08259_),
    .C1(_08144_),
    .X(_08260_));
 sky130_fd_sc_hd__a21oi_1 _15186_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_08123_),
    .B1(_06161_),
    .Y(_08261_));
 sky130_fd_sc_hd__or2_1 _15187_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08237_),
    .X(_08262_));
 sky130_fd_sc_hd__nand2_1 _15188_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08237_),
    .Y(_08263_));
 sky130_fd_sc_hd__nand2_1 _15189_ (.A(_08262_),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__mux2_1 _15190_ (.A0(_08264_),
    .A1(_05059_),
    .S(_08178_),
    .X(_08265_));
 sky130_fd_sc_hd__a22o_2 _15191_ (.A1(_08260_),
    .A2(_08261_),
    .B1(_08265_),
    .B2(_06161_),
    .X(_08266_));
 sky130_fd_sc_hd__clkbuf_4 _15192_ (.A(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__nor2_1 _15193_ (.A(_08255_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__xnor2_1 _15194_ (.A(_08249_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__xnor2_1 _15195_ (.A(_08214_),
    .B(_08269_),
    .Y(_08270_));
 sky130_fd_sc_hd__or4_1 _15196_ (.A(_08222_),
    .B(_08229_),
    .C(_08242_),
    .D(_08254_),
    .X(_08271_));
 sky130_fd_sc_hd__o22ai_1 _15197_ (.A1(_08222_),
    .A2(_08230_),
    .B1(_08243_),
    .B2(_08254_),
    .Y(_08272_));
 sky130_fd_sc_hd__nand2_1 _15198_ (.A(_08271_),
    .B(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__nor2_1 _15199_ (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .B(_08129_),
    .Y(_08274_));
 sky130_fd_sc_hd__a21o_1 _15200_ (.A1(_07893_),
    .A2(_07896_),
    .B1(_08118_),
    .X(_08275_));
 sky130_fd_sc_hd__mux2_1 _15201_ (.A0(_06062_),
    .A1(_06381_),
    .S(_04509_),
    .X(_08276_));
 sky130_fd_sc_hd__a21oi_1 _15202_ (.A1(_08118_),
    .A2(_08276_),
    .B1(_08142_),
    .Y(_08277_));
 sky130_fd_sc_hd__a2bb2o_4 _15203_ (.A1_N(\rbzero.wall_tracer.stepDistY[-8] ),
    .A2_N(_08143_),
    .B1(_08275_),
    .B2(_08277_),
    .X(_08278_));
 sky130_fd_sc_hd__or2_1 _15204_ (.A(_08274_),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__clkbuf_4 _15205_ (.A(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__or3_1 _15206_ (.A(_08266_),
    .B(_08273_),
    .C(_08280_),
    .X(_08281_));
 sky130_fd_sc_hd__nand2_1 _15207_ (.A(_08271_),
    .B(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__or2b_1 _15208_ (.A(_08270_),
    .B_N(_08282_),
    .X(_08283_));
 sky130_fd_sc_hd__a21bo_1 _15209_ (.A1(_08214_),
    .A2(_08269_),
    .B1_N(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__clkbuf_4 _15210_ (.A(_08147_),
    .X(_08285_));
 sky130_fd_sc_hd__buf_4 _15211_ (.A(_08148_),
    .X(_08286_));
 sky130_fd_sc_hd__o22ai_2 _15212_ (.A1(_08127_),
    .A2(_08285_),
    .B1(_08286_),
    .B2(_08138_),
    .Y(_08287_));
 sky130_fd_sc_hd__nand2_1 _15213_ (.A(_08150_),
    .B(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__xnor2_1 _15214_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_08256_),
    .Y(_08289_));
 sky130_fd_sc_hd__nor2_1 _15215_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_06075_),
    .Y(_08290_));
 sky130_fd_sc_hd__a211o_1 _15216_ (.A1(_06075_),
    .A2(_08289_),
    .B1(_08290_),
    .C1(_08144_),
    .X(_08291_));
 sky130_fd_sc_hd__a21oi_1 _15217_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_08123_),
    .B1(_06160_),
    .Y(_08292_));
 sky130_fd_sc_hd__xnor2_1 _15218_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_08262_),
    .Y(_08293_));
 sky130_fd_sc_hd__mux2_1 _15219_ (.A0(_08293_),
    .A1(_05055_),
    .S(_08178_),
    .X(_08294_));
 sky130_fd_sc_hd__a22o_2 _15220_ (.A1(_08291_),
    .A2(_08292_),
    .B1(_08294_),
    .B2(_06160_),
    .X(_08295_));
 sky130_fd_sc_hd__clkbuf_4 _15221_ (.A(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__nor2_1 _15222_ (.A(_08255_),
    .B(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__or3_4 _15223_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .C(_08256_),
    .X(_08298_));
 sky130_fd_sc_hd__o21ai_1 _15224_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_08256_),
    .B1(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_08299_));
 sky130_fd_sc_hd__and2_1 _15225_ (.A(_08298_),
    .B(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__mux2_1 _15226_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(_08300_),
    .S(_06074_),
    .X(_08301_));
 sky130_fd_sc_hd__mux2_1 _15227_ (.A0(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A1(_08301_),
    .S(_08135_),
    .X(_08302_));
 sky130_fd_sc_hd__or3_4 _15228_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .B(\rbzero.debug_overlay.playerX[-2] ),
    .C(_08262_),
    .X(_08303_));
 sky130_fd_sc_hd__o21ai_1 _15229_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_08262_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_08304_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_08303_),
    .B(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__or2_1 _15231_ (.A(_08178_),
    .B(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__a21oi_1 _15232_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_08178_),
    .B1(_08130_),
    .Y(_08307_));
 sky130_fd_sc_hd__a2bb2o_4 _15233_ (.A1_N(_06161_),
    .A2_N(_08302_),
    .B1(_08306_),
    .B2(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__nor2_1 _15234_ (.A(_08280_),
    .B(_08308_),
    .Y(_08309_));
 sky130_fd_sc_hd__xnor2_1 _15235_ (.A(_08297_),
    .B(_08309_),
    .Y(_08310_));
 sky130_fd_sc_hd__inv_2 _15236_ (.A(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_08311_));
 sky130_fd_sc_hd__mux2_1 _15237_ (.A0(_06063_),
    .A1(_06376_),
    .S(_04509_),
    .X(_08312_));
 sky130_fd_sc_hd__and2_1 _15238_ (.A(_08118_),
    .B(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__a21oi_2 _15239_ (.A1(_07880_),
    .A2(_08132_),
    .B1(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__nor2_1 _15240_ (.A(\rbzero.wall_tracer.stepDistX[-9] ),
    .B(_08129_),
    .Y(_08315_));
 sky130_fd_sc_hd__a221o_2 _15241_ (.A1(_08311_),
    .A2(_08135_),
    .B1(_08314_),
    .B2(_08123_),
    .C1(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__clkbuf_4 _15242_ (.A(_08316_),
    .X(_08317_));
 sky130_fd_sc_hd__buf_4 _15243_ (.A(_08144_),
    .X(_08318_));
 sky130_fd_sc_hd__buf_4 _15244_ (.A(_08142_),
    .X(_08319_));
 sky130_fd_sc_hd__o32a_1 _15245_ (.A1(_06081_),
    .A2(_08318_),
    .A3(_08298_),
    .B1(_08319_),
    .B2(_08043_),
    .X(_08320_));
 sky130_fd_sc_hd__o31a_4 _15246_ (.A1(_08130_),
    .A2(_08178_),
    .A3(_08303_),
    .B1(_08320_),
    .X(_08321_));
 sky130_fd_sc_hd__or2_1 _15247_ (.A(_08317_),
    .B(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__xnor2_1 _15248_ (.A(_08310_),
    .B(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__or2_1 _15249_ (.A(_08279_),
    .B(_08296_),
    .X(_08324_));
 sky130_fd_sc_hd__clkbuf_4 _15250_ (.A(_08308_),
    .X(_08325_));
 sky130_fd_sc_hd__o22ai_4 _15251_ (.A1(\rbzero.wall_tracer.stepDistX[-10] ),
    .A2(_08130_),
    .B1(_08145_),
    .B2(_08146_),
    .Y(_08326_));
 sky130_fd_sc_hd__nor2_1 _15252_ (.A(_08321_),
    .B(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__nor2_1 _15253_ (.A(_08308_),
    .B(_08316_),
    .Y(_08328_));
 sky130_fd_sc_hd__xnor2_1 _15254_ (.A(_08324_),
    .B(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__nand2_1 _15255_ (.A(_08327_),
    .B(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__o31a_1 _15256_ (.A1(_08324_),
    .A2(_08325_),
    .A3(_08317_),
    .B1(_08330_),
    .X(_08331_));
 sky130_fd_sc_hd__nor2_1 _15257_ (.A(_08323_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__and2_1 _15258_ (.A(_08323_),
    .B(_08331_),
    .X(_08333_));
 sky130_fd_sc_hd__nor2_1 _15259_ (.A(_08332_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__xnor2_1 _15260_ (.A(_08288_),
    .B(_08334_),
    .Y(_08335_));
 sky130_fd_sc_hd__xnor2_1 _15261_ (.A(_08284_),
    .B(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__xnor2_1 _15262_ (.A(_08327_),
    .B(_08329_),
    .Y(_08337_));
 sky130_fd_sc_hd__nor2_1 _15263_ (.A(_08295_),
    .B(_08326_),
    .Y(_08338_));
 sky130_fd_sc_hd__and2_1 _15264_ (.A(_08328_),
    .B(_08338_),
    .X(_08339_));
 sky130_fd_sc_hd__a21boi_2 _15265_ (.A1(\rbzero.wall_tracer.stepDistX[-11] ),
    .A2(_06162_),
    .B1_N(_08138_),
    .Y(_08340_));
 sky130_fd_sc_hd__clkbuf_4 _15266_ (.A(_08340_),
    .X(_08341_));
 sky130_fd_sc_hd__o22a_1 _15267_ (.A1(_08296_),
    .A2(_08317_),
    .B1(_08326_),
    .B2(_08308_),
    .X(_08342_));
 sky130_fd_sc_hd__nor4_2 _15268_ (.A(_08321_),
    .B(_08339_),
    .C(_08341_),
    .D(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__nor2_1 _15269_ (.A(_08339_),
    .B(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__xnor2_1 _15270_ (.A(_08337_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__or3_2 _15271_ (.A(_08127_),
    .B(_08138_),
    .C(_08345_),
    .X(_08346_));
 sky130_fd_sc_hd__o21ai_1 _15272_ (.A1(_08337_),
    .A2(_08344_),
    .B1(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__or2b_1 _15273_ (.A(_08336_),
    .B_N(_08347_),
    .X(_08348_));
 sky130_fd_sc_hd__a21boi_1 _15274_ (.A1(_08284_),
    .A2(_08335_),
    .B1_N(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__or2_1 _15275_ (.A(_08150_),
    .B(_08349_),
    .X(_08350_));
 sky130_fd_sc_hd__buf_2 _15276_ (.A(_08156_),
    .X(_08351_));
 sky130_fd_sc_hd__clkbuf_4 _15277_ (.A(_08223_),
    .X(_08352_));
 sky130_fd_sc_hd__buf_2 _15278_ (.A(_08177_),
    .X(_08353_));
 sky130_fd_sc_hd__or2_1 _15279_ (.A(_08353_),
    .B(_08243_),
    .X(_08354_));
 sky130_fd_sc_hd__o21ai_1 _15280_ (.A1(_08351_),
    .A2(_08352_),
    .B1(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__nor2_1 _15281_ (.A(_08211_),
    .B(_08267_),
    .Y(_08356_));
 sky130_fd_sc_hd__or3_1 _15282_ (.A(_08351_),
    .B(_08223_),
    .C(_08354_),
    .X(_08357_));
 sky130_fd_sc_hd__a21bo_1 _15283_ (.A1(_08355_),
    .A2(_08356_),
    .B1_N(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__clkbuf_4 _15284_ (.A(_08204_),
    .X(_08359_));
 sky130_fd_sc_hd__buf_4 _15285_ (.A(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__clkinv_2 _15286_ (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_08361_));
 sky130_fd_sc_hd__or3b_2 _15287_ (.A(_07834_),
    .B(_07953_),
    .C_N(_07959_),
    .X(_08362_));
 sky130_fd_sc_hd__xnor2_2 _15288_ (.A(_07966_),
    .B(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__nand2_1 _15289_ (.A(_04510_),
    .B(_08160_),
    .Y(_08364_));
 sky130_fd_sc_hd__o211a_1 _15290_ (.A1(_04510_),
    .A2(_06070_),
    .B1(_08119_),
    .C1(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__a21oi_4 _15291_ (.A1(_08132_),
    .A2(_08363_),
    .B1(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__and3_1 _15292_ (.A(\rbzero.trace_state[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .C(_08142_),
    .X(_08367_));
 sky130_fd_sc_hd__a21oi_4 _15293_ (.A1(_08144_),
    .A2(_08366_),
    .B1(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__mux2_1 _15294_ (.A0(_08361_),
    .A1(_08368_),
    .S(_08130_),
    .X(_08369_));
 sky130_fd_sc_hd__nor2_2 _15295_ (.A(_08171_),
    .B(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__xor2_1 _15296_ (.A(_07953_),
    .B(_07960_),
    .X(_08371_));
 sky130_fd_sc_hd__nor2_1 _15297_ (.A(_04509_),
    .B(_06051_),
    .Y(_08372_));
 sky130_fd_sc_hd__a211o_1 _15298_ (.A1(_04510_),
    .A2(_06396_),
    .B1(_08132_),
    .C1(_08372_),
    .X(_08373_));
 sky130_fd_sc_hd__o21a_4 _15299_ (.A1(_08119_),
    .A2(_08371_),
    .B1(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__nand2_1 _15300_ (.A(\rbzero.wall_tracer.stepDistY[-1] ),
    .B(_08135_),
    .Y(_08375_));
 sky130_fd_sc_hd__nand2_1 _15301_ (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .B(_06161_),
    .Y(_08376_));
 sky130_fd_sc_hd__o211a_2 _15302_ (.A1(_08319_),
    .A2(_08374_),
    .B1(_08375_),
    .C1(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__buf_2 _15303_ (.A(_08377_),
    .X(_08378_));
 sky130_fd_sc_hd__nor2_1 _15304_ (.A(_08191_),
    .B(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__xnor2_2 _15305_ (.A(_08370_),
    .B(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__clkinv_2 _15306_ (.A(_06044_),
    .Y(_08381_));
 sky130_fd_sc_hd__mux2_1 _15307_ (.A0(_08381_),
    .A1(_06341_),
    .S(\rbzero.side_hot ),
    .X(_08382_));
 sky130_fd_sc_hd__mux2_1 _15308_ (.A0(_07953_),
    .A1(_08382_),
    .S(_08118_),
    .X(_08383_));
 sky130_fd_sc_hd__o2bb2a_2 _15309_ (.A1_N(\rbzero.wall_tracer.stepDistY[-2] ),
    .A2_N(_08135_),
    .B1(_08383_),
    .B2(_08142_),
    .X(_08384_));
 sky130_fd_sc_hd__clkbuf_4 _15310_ (.A(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__a21boi_2 _15311_ (.A1(\rbzero.wall_tracer.stepDistX[-2] ),
    .A2(_06161_),
    .B1_N(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__clkbuf_4 _15312_ (.A(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__nand2_1 _15313_ (.A(_08370_),
    .B(_08379_),
    .Y(_08388_));
 sky130_fd_sc_hd__o31ai_4 _15314_ (.A1(_08360_),
    .A2(_08380_),
    .A3(_08387_),
    .B1(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__nor2_1 _15315_ (.A(_08351_),
    .B(_08243_),
    .Y(_08390_));
 sky130_fd_sc_hd__nor2_1 _15316_ (.A(_08223_),
    .B(_08387_),
    .Y(_08391_));
 sky130_fd_sc_hd__xnor2_1 _15317_ (.A(_08390_),
    .B(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__or3_1 _15318_ (.A(_08353_),
    .B(_08267_),
    .C(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__clkbuf_4 _15319_ (.A(_08267_),
    .X(_08394_));
 sky130_fd_sc_hd__o21ai_1 _15320_ (.A1(_08353_),
    .A2(_08394_),
    .B1(_08392_),
    .Y(_08395_));
 sky130_fd_sc_hd__nand2_1 _15321_ (.A(_08393_),
    .B(_08395_),
    .Y(_08396_));
 sky130_fd_sc_hd__xor2_1 _15322_ (.A(_08389_),
    .B(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__xnor2_1 _15323_ (.A(_08358_),
    .B(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__clkbuf_4 _15324_ (.A(_08191_),
    .X(_08399_));
 sky130_fd_sc_hd__mux2_1 _15325_ (.A0(_06039_),
    .A1(_06331_),
    .S(_04510_),
    .X(_08400_));
 sky130_fd_sc_hd__nand2_2 _15326_ (.A(_08119_),
    .B(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__a21o_1 _15327_ (.A1(_07966_),
    .A2(_08362_),
    .B1(_07971_),
    .X(_08402_));
 sky130_fd_sc_hd__nand3_1 _15328_ (.A(_07966_),
    .B(_07971_),
    .C(_08362_),
    .Y(_08403_));
 sky130_fd_sc_hd__a21o_1 _15329_ (.A1(_08402_),
    .A2(_08403_),
    .B1(_08119_),
    .X(_08404_));
 sky130_fd_sc_hd__a21o_4 _15330_ (.A1(_08401_),
    .A2(_08404_),
    .B1(_08319_),
    .X(_08405_));
 sky130_fd_sc_hd__buf_6 _15331_ (.A(_08135_),
    .X(_08406_));
 sky130_fd_sc_hd__a22oi_2 _15332_ (.A1(\rbzero.wall_tracer.stepDistX[1] ),
    .A2(_06161_),
    .B1(_08406_),
    .B2(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_08407_));
 sky130_fd_sc_hd__and2_1 _15333_ (.A(_08405_),
    .B(_08407_),
    .X(_08408_));
 sky130_fd_sc_hd__clkbuf_4 _15334_ (.A(_08408_),
    .X(_08409_));
 sky130_fd_sc_hd__nor2_2 _15335_ (.A(_08399_),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__buf_2 _15336_ (.A(_08369_),
    .X(_08411_));
 sky130_fd_sc_hd__clkbuf_4 _15337_ (.A(_08171_),
    .X(_08412_));
 sky130_fd_sc_hd__o22ai_1 _15338_ (.A1(_08399_),
    .A2(_08411_),
    .B1(_08409_),
    .B2(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__a21bo_1 _15339_ (.A1(_08370_),
    .A2(_08410_),
    .B1_N(_08413_),
    .X(_08414_));
 sky130_fd_sc_hd__nor2_1 _15340_ (.A(_08359_),
    .B(_08378_),
    .Y(_08415_));
 sky130_fd_sc_hd__xnor2_2 _15341_ (.A(_08414_),
    .B(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__inv_2 _15342_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_08417_));
 sky130_fd_sc_hd__nor2_1 _15343_ (.A(_08417_),
    .B(_08143_),
    .Y(_08418_));
 sky130_fd_sc_hd__a221oi_4 _15344_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_06158_),
    .B1(_06160_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__clkbuf_4 _15345_ (.A(_08419_),
    .X(_08420_));
 sky130_fd_sc_hd__xor2_1 _15346_ (.A(_07976_),
    .B(_08402_),
    .X(_08421_));
 sky130_fd_sc_hd__nor2_1 _15347_ (.A(_04511_),
    .B(_06035_),
    .Y(_08422_));
 sky130_fd_sc_hd__a211o_1 _15348_ (.A1(_04511_),
    .A2(_06327_),
    .B1(_08132_),
    .C1(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__o21ai_4 _15349_ (.A1(_08119_),
    .A2(_08421_),
    .B1(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__a22o_1 _15350_ (.A1(\rbzero.wall_tracer.stepDistX[2] ),
    .A2(_06161_),
    .B1(_08406_),
    .B2(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_08425_));
 sky130_fd_sc_hd__a21oi_2 _15351_ (.A1(_08124_),
    .A2(_08424_),
    .B1(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__clkbuf_4 _15352_ (.A(_08426_),
    .X(_08427_));
 sky130_fd_sc_hd__nor2_1 _15353_ (.A(_08420_),
    .B(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__clkbuf_4 _15354_ (.A(_08132_),
    .X(_08429_));
 sky130_fd_sc_hd__a2111o_1 _15355_ (.A1(_07966_),
    .A2(_08362_),
    .B1(_07983_),
    .C1(_07976_),
    .D1(_07971_),
    .X(_08430_));
 sky130_fd_sc_hd__buf_2 _15356_ (.A(_08430_),
    .X(_08431_));
 sky130_fd_sc_hd__o21ai_1 _15357_ (.A1(_07976_),
    .A2(_08402_),
    .B1(_07983_),
    .Y(_08432_));
 sky130_fd_sc_hd__mux2_2 _15358_ (.A0(_06073_),
    .A1(_06413_),
    .S(_04510_),
    .X(_08433_));
 sky130_fd_sc_hd__a21o_1 _15359_ (.A1(_08119_),
    .A2(_08433_),
    .B1(_08135_),
    .X(_08434_));
 sky130_fd_sc_hd__a31o_1 _15360_ (.A1(_08429_),
    .A2(_08431_),
    .A3(_08432_),
    .B1(_08434_),
    .X(_08435_));
 sky130_fd_sc_hd__nand2_2 _15361_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08123_),
    .Y(_08436_));
 sky130_fd_sc_hd__buf_2 _15362_ (.A(_08436_),
    .X(_08437_));
 sky130_fd_sc_hd__nor2_1 _15363_ (.A(_08435_),
    .B(_08437_),
    .Y(_08438_));
 sky130_fd_sc_hd__nor2_2 _15364_ (.A(_08018_),
    .B(_08142_),
    .Y(_08439_));
 sky130_fd_sc_hd__nand2_1 _15365_ (.A(\rbzero.wall_tracer.stepDistY[4] ),
    .B(_08135_),
    .Y(_08440_));
 sky130_fd_sc_hd__nand2_1 _15366_ (.A(_07989_),
    .B(_08431_),
    .Y(_08441_));
 sky130_fd_sc_hd__or2_1 _15367_ (.A(_07989_),
    .B(_08431_),
    .X(_08442_));
 sky130_fd_sc_hd__a31o_1 _15368_ (.A1(_08132_),
    .A2(_08441_),
    .A3(_08442_),
    .B1(_08434_),
    .X(_08443_));
 sky130_fd_sc_hd__nand2_1 _15369_ (.A(_08440_),
    .B(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__nand2_1 _15370_ (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .B(_08319_),
    .Y(_08445_));
 sky130_fd_sc_hd__a21o_1 _15371_ (.A1(_08435_),
    .A2(_08445_),
    .B1(_06162_),
    .X(_08446_));
 sky130_fd_sc_hd__nand2_4 _15372_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_08144_),
    .Y(_08447_));
 sky130_fd_sc_hd__a21o_2 _15373_ (.A1(_08440_),
    .A2(_08443_),
    .B1(_06162_),
    .X(_08448_));
 sky130_fd_sc_hd__nand2_1 _15374_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08143_),
    .Y(_08449_));
 sky130_fd_sc_hd__clkbuf_4 _15375_ (.A(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__o22a_1 _15376_ (.A1(_08446_),
    .A2(_08447_),
    .B1(_08448_),
    .B2(_08450_),
    .X(_08451_));
 sky130_fd_sc_hd__a31oi_2 _15377_ (.A1(_08438_),
    .A2(_08439_),
    .A3(_08444_),
    .B1(_08451_),
    .Y(_08452_));
 sky130_fd_sc_hd__xnor2_2 _15378_ (.A(_08428_),
    .B(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__clkbuf_4 _15379_ (.A(_08446_),
    .X(_08454_));
 sky130_fd_sc_hd__nand2_1 _15380_ (.A(_08424_),
    .B(_08439_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand2_1 _15381_ (.A(_08405_),
    .B(_08407_),
    .Y(_08456_));
 sky130_fd_sc_hd__a221o_4 _15382_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08123_),
    .B1(_06161_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08418_),
    .X(_08457_));
 sky130_fd_sc_hd__nand2_1 _15383_ (.A(_08456_),
    .B(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__xnor2_1 _15384_ (.A(_08438_),
    .B(_08455_),
    .Y(_08459_));
 sky130_fd_sc_hd__or2b_1 _15385_ (.A(_08458_),
    .B_N(_08459_),
    .X(_08460_));
 sky130_fd_sc_hd__o31a_1 _15386_ (.A1(_08450_),
    .A2(_08454_),
    .A3(_08455_),
    .B1(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__xor2_2 _15387_ (.A(_08453_),
    .B(_08461_),
    .X(_08462_));
 sky130_fd_sc_hd__xnor2_2 _15388_ (.A(_08416_),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nor2_1 _15389_ (.A(_08359_),
    .B(_08387_),
    .Y(_08464_));
 sky130_fd_sc_hd__xnor2_2 _15390_ (.A(_08380_),
    .B(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__xor2_2 _15391_ (.A(_08458_),
    .B(_08459_),
    .X(_08466_));
 sky130_fd_sc_hd__or4b_1 _15392_ (.A(_08018_),
    .B(_08405_),
    .C(_08437_),
    .D_N(_08424_),
    .X(_08467_));
 sky130_fd_sc_hd__nor2_1 _15393_ (.A(_06160_),
    .B(_08450_),
    .Y(_08468_));
 sky130_fd_sc_hd__a2bb2o_1 _15394_ (.A1_N(_08018_),
    .A2_N(_08405_),
    .B1(_08424_),
    .B2(_08468_),
    .X(_08469_));
 sky130_fd_sc_hd__or4bb_1 _15395_ (.A(_08369_),
    .B(_08419_),
    .C_N(_08467_),
    .D_N(_08469_),
    .X(_08470_));
 sky130_fd_sc_hd__and2_1 _15396_ (.A(_08467_),
    .B(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__xor2_2 _15397_ (.A(_08466_),
    .B(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__nor2_1 _15398_ (.A(_08466_),
    .B(_08471_),
    .Y(_08473_));
 sky130_fd_sc_hd__a21o_1 _15399_ (.A1(_08465_),
    .A2(_08472_),
    .B1(_08473_),
    .X(_08474_));
 sky130_fd_sc_hd__xnor2_1 _15400_ (.A(_08463_),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__xnor2_1 _15401_ (.A(_08398_),
    .B(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__xnor2_2 _15402_ (.A(_08465_),
    .B(_08472_),
    .Y(_08477_));
 sky130_fd_sc_hd__a2bb2o_1 _15403_ (.A1_N(_08411_),
    .A2_N(_08420_),
    .B1(_08467_),
    .B2(_08469_),
    .X(_08478_));
 sky130_fd_sc_hd__and2_4 _15404_ (.A(_08401_),
    .B(_08404_),
    .X(_08479_));
 sky130_fd_sc_hd__nand2_4 _15405_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_06158_),
    .Y(_08480_));
 sky130_fd_sc_hd__o22ai_2 _15406_ (.A1(_08479_),
    .A2(_08437_),
    .B1(_08480_),
    .B2(_08368_),
    .Y(_08481_));
 sky130_fd_sc_hd__nor2_1 _15407_ (.A(_08377_),
    .B(_08419_),
    .Y(_08482_));
 sky130_fd_sc_hd__and3_1 _15408_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08123_),
    .C(_08366_),
    .X(_08483_));
 sky130_fd_sc_hd__or3b_1 _15409_ (.A(_08018_),
    .B(_08405_),
    .C_N(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__a21bo_1 _15410_ (.A1(_08481_),
    .A2(_08482_),
    .B1_N(_08484_),
    .X(_08485_));
 sky130_fd_sc_hd__nand3_1 _15411_ (.A(_08470_),
    .B(_08478_),
    .C(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__a21o_1 _15412_ (.A1(_08470_),
    .A2(_08478_),
    .B1(_08485_),
    .X(_08487_));
 sky130_fd_sc_hd__nor2_1 _15413_ (.A(_08171_),
    .B(_08387_),
    .Y(_08488_));
 sky130_fd_sc_hd__or3b_1 _15414_ (.A(_08191_),
    .B(_08377_),
    .C_N(_08488_),
    .X(_08489_));
 sky130_fd_sc_hd__o22ai_1 _15415_ (.A1(_08171_),
    .A2(_08377_),
    .B1(_08387_),
    .B2(_08399_),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_1 _15416_ (.A(_08489_),
    .B(_08490_),
    .Y(_08491_));
 sky130_fd_sc_hd__nor2_1 _15417_ (.A(_08351_),
    .B(_08204_),
    .Y(_08492_));
 sky130_fd_sc_hd__xnor2_1 _15418_ (.A(_08491_),
    .B(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__nand3_1 _15419_ (.A(_08486_),
    .B(_08487_),
    .C(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__and2_1 _15420_ (.A(_08486_),
    .B(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__xor2_1 _15421_ (.A(_08477_),
    .B(_08495_),
    .X(_08496_));
 sky130_fd_sc_hd__nor2_2 _15422_ (.A(_08205_),
    .B(_08209_),
    .Y(_08497_));
 sky130_fd_sc_hd__a2bb2o_1 _15423_ (.A1_N(_08353_),
    .A2_N(_08223_),
    .B1(_08247_),
    .B2(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__nor2_1 _15424_ (.A(_08230_),
    .B(_08267_),
    .Y(_08499_));
 sky130_fd_sc_hd__or3_1 _15425_ (.A(_08211_),
    .B(_08223_),
    .C(_08354_),
    .X(_08500_));
 sky130_fd_sc_hd__a21bo_1 _15426_ (.A1(_08498_),
    .A2(_08499_),
    .B1_N(_08500_),
    .X(_08501_));
 sky130_fd_sc_hd__a21bo_1 _15427_ (.A1(_08490_),
    .A2(_08492_),
    .B1_N(_08489_),
    .X(_08502_));
 sky130_fd_sc_hd__and2_1 _15428_ (.A(_08357_),
    .B(_08355_),
    .X(_08503_));
 sky130_fd_sc_hd__xnor2_1 _15429_ (.A(_08503_),
    .B(_08356_),
    .Y(_08504_));
 sky130_fd_sc_hd__xor2_1 _15430_ (.A(_08502_),
    .B(_08504_),
    .X(_08505_));
 sky130_fd_sc_hd__xnor2_1 _15431_ (.A(_08501_),
    .B(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__nor2_1 _15432_ (.A(_08477_),
    .B(_08495_),
    .Y(_08507_));
 sky130_fd_sc_hd__a21o_1 _15433_ (.A1(_08496_),
    .A2(_08506_),
    .B1(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__xnor2_1 _15434_ (.A(_08476_),
    .B(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__or4_1 _15435_ (.A(_08230_),
    .B(_08255_),
    .C(_08296_),
    .D(_08308_),
    .X(_08510_));
 sky130_fd_sc_hd__o21ai_2 _15436_ (.A1(\rbzero.wall_tracer.stepDistY[-7] ),
    .A2(_08318_),
    .B1(_08253_),
    .Y(_08511_));
 sky130_fd_sc_hd__inv_2 _15437_ (.A(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__clkinv_2 _15438_ (.A(_08308_),
    .Y(_08513_));
 sky130_fd_sc_hd__nor2_1 _15439_ (.A(_08230_),
    .B(_08296_),
    .Y(_08514_));
 sky130_fd_sc_hd__a31o_1 _15440_ (.A1(_08250_),
    .A2(_08512_),
    .A3(_08513_),
    .B1(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__nand2_1 _15441_ (.A(_08510_),
    .B(_08515_),
    .Y(_08516_));
 sky130_fd_sc_hd__or2_1 _15442_ (.A(_08280_),
    .B(_08321_),
    .X(_08517_));
 sky130_fd_sc_hd__xnor2_1 _15443_ (.A(_08516_),
    .B(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__o2bb2a_1 _15444_ (.A1_N(_08297_),
    .A2_N(_08309_),
    .B1(_08310_),
    .B2(_08322_),
    .X(_08519_));
 sky130_fd_sc_hd__a22o_4 _15445_ (.A1(_08311_),
    .A2(_08406_),
    .B1(_08314_),
    .B2(_08124_),
    .X(_08520_));
 sky130_fd_sc_hd__nor2_1 _15446_ (.A(_08125_),
    .B(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__xnor2_1 _15447_ (.A(_08149_),
    .B(_08521_),
    .Y(_08522_));
 sky130_fd_sc_hd__buf_4 _15448_ (.A(_08124_),
    .X(_08523_));
 sky130_fd_sc_hd__nand2_2 _15449_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08523_),
    .Y(_08524_));
 sky130_fd_sc_hd__nor2_1 _15450_ (.A(_08138_),
    .B(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__nand2_1 _15451_ (.A(_08522_),
    .B(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__or2_1 _15452_ (.A(_08522_),
    .B(_08525_),
    .X(_08527_));
 sky130_fd_sc_hd__and2_1 _15453_ (.A(_08526_),
    .B(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__xor2_1 _15454_ (.A(_08518_),
    .B(_08519_),
    .X(_08529_));
 sky130_fd_sc_hd__nand2_1 _15455_ (.A(_08528_),
    .B(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__o21ai_1 _15456_ (.A1(_08518_),
    .A2(_08519_),
    .B1(_08530_),
    .Y(_08531_));
 sky130_fd_sc_hd__or2b_1 _15457_ (.A(_08504_),
    .B_N(_08502_),
    .X(_08532_));
 sky130_fd_sc_hd__or2b_1 _15458_ (.A(_08505_),
    .B_N(_08501_),
    .X(_08533_));
 sky130_fd_sc_hd__clkbuf_4 _15459_ (.A(_08524_),
    .X(_08534_));
 sky130_fd_sc_hd__o22ai_1 _15460_ (.A1(_08125_),
    .A2(_08278_),
    .B1(_08520_),
    .B2(_08148_),
    .Y(_08535_));
 sky130_fd_sc_hd__or4_1 _15461_ (.A(_08125_),
    .B(_08148_),
    .C(_08278_),
    .D(_08520_),
    .X(_08536_));
 sky130_fd_sc_hd__nand2_1 _15462_ (.A(_08535_),
    .B(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__or3_1 _15463_ (.A(_08147_),
    .B(_08534_),
    .C(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__o21ai_1 _15464_ (.A1(_08285_),
    .A2(_08534_),
    .B1(_08537_),
    .Y(_08539_));
 sky130_fd_sc_hd__and2_1 _15465_ (.A(_08538_),
    .B(_08539_),
    .X(_08540_));
 sky130_fd_sc_hd__nor2_1 _15466_ (.A(_08211_),
    .B(_08325_),
    .Y(_08541_));
 sky130_fd_sc_hd__o22a_1 _15467_ (.A1(_08211_),
    .A2(_08296_),
    .B1(_08308_),
    .B2(_08230_),
    .X(_08542_));
 sky130_fd_sc_hd__a21o_1 _15468_ (.A1(_08514_),
    .A2(_08541_),
    .B1(_08542_),
    .X(_08543_));
 sky130_fd_sc_hd__or2_1 _15469_ (.A(_08255_),
    .B(_08321_),
    .X(_08544_));
 sky130_fd_sc_hd__xnor2_1 _15470_ (.A(_08543_),
    .B(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__buf_2 _15471_ (.A(_08321_),
    .X(_08546_));
 sky130_fd_sc_hd__o31a_1 _15472_ (.A1(_08280_),
    .A2(_08546_),
    .A3(_08516_),
    .B1(_08510_),
    .X(_08547_));
 sky130_fd_sc_hd__nor2_1 _15473_ (.A(_08545_),
    .B(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__and2_1 _15474_ (.A(_08545_),
    .B(_08547_),
    .X(_08549_));
 sky130_fd_sc_hd__nor2_1 _15475_ (.A(_08548_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__xnor2_1 _15476_ (.A(_08540_),
    .B(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__a21o_1 _15477_ (.A1(_08532_),
    .A2(_08533_),
    .B1(_08551_),
    .X(_08552_));
 sky130_fd_sc_hd__nand3_1 _15478_ (.A(_08532_),
    .B(_08533_),
    .C(_08551_),
    .Y(_08553_));
 sky130_fd_sc_hd__nand2_1 _15479_ (.A(_08552_),
    .B(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__xnor2_1 _15480_ (.A(_08531_),
    .B(_08554_),
    .Y(_08555_));
 sky130_fd_sc_hd__xnor2_1 _15481_ (.A(_08509_),
    .B(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__xnor2_1 _15482_ (.A(_08496_),
    .B(_08506_),
    .Y(_08557_));
 sky130_fd_sc_hd__a21o_1 _15483_ (.A1(_08486_),
    .A2(_08487_),
    .B1(_08493_),
    .X(_08558_));
 sky130_fd_sc_hd__nand3_1 _15484_ (.A(_08484_),
    .B(_08481_),
    .C(_08482_),
    .Y(_08559_));
 sky130_fd_sc_hd__a21o_1 _15485_ (.A1(_08484_),
    .A2(_08481_),
    .B1(_08482_),
    .X(_08560_));
 sky130_fd_sc_hd__nor2_1 _15486_ (.A(_08374_),
    .B(_08480_),
    .Y(_08561_));
 sky130_fd_sc_hd__xor2_1 _15487_ (.A(_08483_),
    .B(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__nor2_1 _15488_ (.A(_08386_),
    .B(_08419_),
    .Y(_08563_));
 sky130_fd_sc_hd__nand2_1 _15489_ (.A(_08483_),
    .B(_08561_),
    .Y(_08564_));
 sky130_fd_sc_hd__a21bo_1 _15490_ (.A1(_08562_),
    .A2(_08563_),
    .B1_N(_08564_),
    .X(_08565_));
 sky130_fd_sc_hd__a21o_1 _15491_ (.A1(_08559_),
    .A2(_08560_),
    .B1(_08565_),
    .X(_08566_));
 sky130_fd_sc_hd__nor2_1 _15492_ (.A(_08351_),
    .B(_08191_),
    .Y(_08567_));
 sky130_fd_sc_hd__xnor2_1 _15493_ (.A(_08567_),
    .B(_08488_),
    .Y(_08568_));
 sky130_fd_sc_hd__or3_1 _15494_ (.A(_08353_),
    .B(_08204_),
    .C(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__o21ai_1 _15495_ (.A1(_08353_),
    .A2(_08204_),
    .B1(_08568_),
    .Y(_08570_));
 sky130_fd_sc_hd__and2_1 _15496_ (.A(_08569_),
    .B(_08570_),
    .X(_08571_));
 sky130_fd_sc_hd__and3_1 _15497_ (.A(_08559_),
    .B(_08560_),
    .C(_08565_),
    .X(_08572_));
 sky130_fd_sc_hd__a21o_1 _15498_ (.A1(_08566_),
    .A2(_08571_),
    .B1(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__a21o_1 _15499_ (.A1(_08494_),
    .A2(_08558_),
    .B1(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__a21bo_1 _15500_ (.A1(_08248_),
    .A2(_08268_),
    .B1_N(_08244_),
    .X(_08575_));
 sky130_fd_sc_hd__a21bo_1 _15501_ (.A1(_08567_),
    .A2(_08488_),
    .B1_N(_08569_),
    .X(_08576_));
 sky130_fd_sc_hd__nand2_1 _15502_ (.A(_08500_),
    .B(_08498_),
    .Y(_08577_));
 sky130_fd_sc_hd__xor2_1 _15503_ (.A(_08577_),
    .B(_08499_),
    .X(_08578_));
 sky130_fd_sc_hd__xor2_1 _15504_ (.A(_08576_),
    .B(_08578_),
    .X(_08579_));
 sky130_fd_sc_hd__xnor2_1 _15505_ (.A(_08575_),
    .B(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__nand3_1 _15506_ (.A(_08494_),
    .B(_08558_),
    .C(_08573_),
    .Y(_08581_));
 sky130_fd_sc_hd__a21boi_1 _15507_ (.A1(_08574_),
    .A2(_08580_),
    .B1_N(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__nor2_1 _15508_ (.A(_08557_),
    .B(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__and2_1 _15509_ (.A(_08557_),
    .B(_08582_),
    .X(_08584_));
 sky130_fd_sc_hd__nor2_1 _15510_ (.A(_08583_),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__a31o_1 _15511_ (.A1(_08150_),
    .A2(_08287_),
    .A3(_08334_),
    .B1(_08332_),
    .X(_08586_));
 sky130_fd_sc_hd__or2b_1 _15512_ (.A(_08578_),
    .B_N(_08576_),
    .X(_08587_));
 sky130_fd_sc_hd__or2b_1 _15513_ (.A(_08579_),
    .B_N(_08575_),
    .X(_08588_));
 sky130_fd_sc_hd__or2_1 _15514_ (.A(_08528_),
    .B(_08529_),
    .X(_08589_));
 sky130_fd_sc_hd__nand2_1 _15515_ (.A(_08530_),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__a21o_1 _15516_ (.A1(_08587_),
    .A2(_08588_),
    .B1(_08590_),
    .X(_08591_));
 sky130_fd_sc_hd__nand3_1 _15517_ (.A(_08587_),
    .B(_08588_),
    .C(_08590_),
    .Y(_08592_));
 sky130_fd_sc_hd__nand2_1 _15518_ (.A(_08591_),
    .B(_08592_),
    .Y(_08593_));
 sky130_fd_sc_hd__xnor2_1 _15519_ (.A(_08586_),
    .B(_08593_),
    .Y(_08594_));
 sky130_fd_sc_hd__a21oi_1 _15520_ (.A1(_08585_),
    .A2(_08594_),
    .B1(_08583_),
    .Y(_08595_));
 sky130_fd_sc_hd__xor2_1 _15521_ (.A(_08556_),
    .B(_08595_),
    .X(_08596_));
 sky130_fd_sc_hd__or2b_1 _15522_ (.A(_08593_),
    .B_N(_08586_),
    .X(_08597_));
 sky130_fd_sc_hd__buf_4 _15523_ (.A(_08138_),
    .X(_08598_));
 sky130_fd_sc_hd__nand2_4 _15524_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08124_),
    .Y(_08599_));
 sky130_fd_sc_hd__clkbuf_4 _15525_ (.A(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__or2_1 _15526_ (.A(_08598_),
    .B(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__buf_2 _15527_ (.A(_08520_),
    .X(_08602_));
 sky130_fd_sc_hd__o31a_1 _15528_ (.A1(_08127_),
    .A2(_08149_),
    .A3(_08602_),
    .B1(_08526_),
    .X(_08603_));
 sky130_fd_sc_hd__nor2_1 _15529_ (.A(_08601_),
    .B(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__and2_1 _15530_ (.A(_08601_),
    .B(_08603_),
    .X(_08605_));
 sky130_fd_sc_hd__or2_1 _15531_ (.A(_08604_),
    .B(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__a21oi_2 _15532_ (.A1(_08591_),
    .A2(_08597_),
    .B1(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__and3_1 _15533_ (.A(_08591_),
    .B(_08597_),
    .C(_08606_),
    .X(_08608_));
 sky130_fd_sc_hd__nor2_1 _15534_ (.A(_08607_),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__xnor2_1 _15535_ (.A(_08596_),
    .B(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__xnor2_1 _15536_ (.A(_08585_),
    .B(_08594_),
    .Y(_08611_));
 sky130_fd_sc_hd__and3_1 _15537_ (.A(_08581_),
    .B(_08574_),
    .C(_08580_),
    .X(_08612_));
 sky130_fd_sc_hd__a21oi_1 _15538_ (.A1(_08581_),
    .A2(_08574_),
    .B1(_08580_),
    .Y(_08613_));
 sky130_fd_sc_hd__or2_1 _15539_ (.A(_08612_),
    .B(_08613_),
    .X(_08614_));
 sky130_fd_sc_hd__and2b_1 _15540_ (.A_N(_08572_),
    .B(_08566_),
    .X(_08615_));
 sky130_fd_sc_hd__xnor2_1 _15541_ (.A(_08615_),
    .B(_08571_),
    .Y(_08616_));
 sky130_fd_sc_hd__xnor2_1 _15542_ (.A(_08562_),
    .B(_08563_),
    .Y(_08617_));
 sky130_fd_sc_hd__inv_2 _15543_ (.A(_08449_),
    .Y(_08618_));
 sky130_fd_sc_hd__and4bb_1 _15544_ (.A_N(_08374_),
    .B_N(_08384_),
    .C(_08618_),
    .D(_08439_),
    .X(_08619_));
 sky130_fd_sc_hd__or2_1 _15545_ (.A(_08156_),
    .B(_08419_),
    .X(_08620_));
 sky130_fd_sc_hd__o22a_1 _15546_ (.A1(_08374_),
    .A2(_08436_),
    .B1(_08447_),
    .B2(_08384_),
    .X(_08621_));
 sky130_fd_sc_hd__or3_1 _15547_ (.A(_08619_),
    .B(_08620_),
    .C(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__and2b_1 _15548_ (.A_N(_08619_),
    .B(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__xor2_1 _15549_ (.A(_08617_),
    .B(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__nand2_1 _15550_ (.A(_08213_),
    .B(_08192_),
    .Y(_08625_));
 sky130_fd_sc_hd__xnor2_1 _15551_ (.A(_08625_),
    .B(_08212_),
    .Y(_08626_));
 sky130_fd_sc_hd__nor2_1 _15552_ (.A(_08617_),
    .B(_08623_),
    .Y(_08627_));
 sky130_fd_sc_hd__a21oi_1 _15553_ (.A1(_08624_),
    .A2(_08626_),
    .B1(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__xor2_1 _15554_ (.A(_08616_),
    .B(_08628_),
    .X(_08629_));
 sky130_fd_sc_hd__xnor2_1 _15555_ (.A(_08282_),
    .B(_08270_),
    .Y(_08630_));
 sky130_fd_sc_hd__nor2_1 _15556_ (.A(_08616_),
    .B(_08628_),
    .Y(_08631_));
 sky130_fd_sc_hd__a21oi_2 _15557_ (.A1(_08629_),
    .A2(_08630_),
    .B1(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__xor2_1 _15558_ (.A(_08614_),
    .B(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__xnor2_1 _15559_ (.A(_08347_),
    .B(_08336_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand2_1 _15560_ (.A(_08633_),
    .B(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__o21a_1 _15561_ (.A1(_08614_),
    .A2(_08632_),
    .B1(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__xor2_1 _15562_ (.A(_08611_),
    .B(_08636_),
    .X(_08637_));
 sky130_fd_sc_hd__nand2_1 _15563_ (.A(_08150_),
    .B(_08349_),
    .Y(_08638_));
 sky130_fd_sc_hd__and2_1 _15564_ (.A(_08350_),
    .B(_08638_),
    .X(_08639_));
 sky130_fd_sc_hd__o2bb2a_1 _15565_ (.A1_N(_08637_),
    .A2_N(_08639_),
    .B1(_08611_),
    .B2(_08636_),
    .X(_08640_));
 sky130_fd_sc_hd__xor2_1 _15566_ (.A(_08610_),
    .B(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__xnor2_2 _15567_ (.A(_08350_),
    .B(_08641_),
    .Y(_08642_));
 sky130_fd_sc_hd__or2_1 _15568_ (.A(_08633_),
    .B(_08634_),
    .X(_08643_));
 sky130_fd_sc_hd__nand2_1 _15569_ (.A(_08635_),
    .B(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__xnor2_1 _15570_ (.A(_08629_),
    .B(_08630_),
    .Y(_08645_));
 sky130_fd_sc_hd__xnor2_1 _15571_ (.A(_08624_),
    .B(_08626_),
    .Y(_08646_));
 sky130_fd_sc_hd__o21ai_1 _15572_ (.A1(_08619_),
    .A2(_08621_),
    .B1(_08620_),
    .Y(_08647_));
 sky130_fd_sc_hd__or4_1 _15573_ (.A(_08155_),
    .B(_08384_),
    .C(_08450_),
    .D(_08480_),
    .X(_08648_));
 sky130_fd_sc_hd__buf_4 _15574_ (.A(_08155_),
    .X(_08649_));
 sky130_fd_sc_hd__o22ai_1 _15575_ (.A1(_08385_),
    .A2(_08450_),
    .B1(_08480_),
    .B2(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__or4bb_1 _15576_ (.A(_08177_),
    .B(_08419_),
    .C_N(_08648_),
    .D_N(_08650_),
    .X(_08651_));
 sky130_fd_sc_hd__nand2_1 _15577_ (.A(_08648_),
    .B(_08651_),
    .Y(_08652_));
 sky130_fd_sc_hd__nand3_1 _15578_ (.A(_08622_),
    .B(_08647_),
    .C(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__or2_1 _15579_ (.A(_08204_),
    .B(_08230_),
    .X(_08654_));
 sky130_fd_sc_hd__or3_1 _15580_ (.A(_08170_),
    .B(_08205_),
    .C(_08209_),
    .X(_08655_));
 sky130_fd_sc_hd__or3_1 _15581_ (.A(_08191_),
    .B(_08177_),
    .C(_08655_),
    .X(_08656_));
 sky130_fd_sc_hd__inv_2 _15582_ (.A(_08190_),
    .Y(_08657_));
 sky130_fd_sc_hd__a2bb2o_1 _15583_ (.A1_N(_08170_),
    .A2_N(_08177_),
    .B1(_08497_),
    .B2(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__nand2_1 _15584_ (.A(_08656_),
    .B(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__xor2_1 _15585_ (.A(_08654_),
    .B(_08659_),
    .X(_08660_));
 sky130_fd_sc_hd__a21o_1 _15586_ (.A1(_08622_),
    .A2(_08647_),
    .B1(_08652_),
    .X(_08661_));
 sky130_fd_sc_hd__nand3_1 _15587_ (.A(_08653_),
    .B(_08660_),
    .C(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__and2_1 _15588_ (.A(_08653_),
    .B(_08662_),
    .X(_08663_));
 sky130_fd_sc_hd__xor2_1 _15589_ (.A(_08646_),
    .B(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__nor2_1 _15590_ (.A(_08266_),
    .B(_08317_),
    .Y(_08665_));
 sky130_fd_sc_hd__nor2_1 _15591_ (.A(_08222_),
    .B(_08254_),
    .Y(_08666_));
 sky130_fd_sc_hd__or2_1 _15592_ (.A(_08242_),
    .B(_08279_),
    .X(_08667_));
 sky130_fd_sc_hd__xnor2_1 _15593_ (.A(_08666_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__or3_1 _15594_ (.A(_08223_),
    .B(_08255_),
    .C(_08667_),
    .X(_08669_));
 sky130_fd_sc_hd__a21bo_1 _15595_ (.A1(_08665_),
    .A2(_08668_),
    .B1_N(_08669_),
    .X(_08670_));
 sky130_fd_sc_hd__o21ai_1 _15596_ (.A1(_08654_),
    .A2(_08659_),
    .B1(_08656_),
    .Y(_08671_));
 sky130_fd_sc_hd__o21ai_1 _15597_ (.A1(_08267_),
    .A2(_08280_),
    .B1(_08273_),
    .Y(_08672_));
 sky130_fd_sc_hd__nand2_1 _15598_ (.A(_08281_),
    .B(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__xor2_1 _15599_ (.A(_08671_),
    .B(_08673_),
    .X(_08674_));
 sky130_fd_sc_hd__xnor2_1 _15600_ (.A(_08670_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__nor2_1 _15601_ (.A(_08646_),
    .B(_08663_),
    .Y(_08676_));
 sky130_fd_sc_hd__a21oi_1 _15602_ (.A1(_08664_),
    .A2(_08675_),
    .B1(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__xor2_1 _15603_ (.A(_08645_),
    .B(_08677_),
    .X(_08678_));
 sky130_fd_sc_hd__nor2_1 _15604_ (.A(_08325_),
    .B(_08341_),
    .Y(_08679_));
 sky130_fd_sc_hd__nand2_1 _15605_ (.A(_08338_),
    .B(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__o22a_1 _15606_ (.A1(_08546_),
    .A2(_08341_),
    .B1(_08342_),
    .B2(_08339_),
    .X(_08681_));
 sky130_fd_sc_hd__or3_1 _15607_ (.A(_08343_),
    .B(_08680_),
    .C(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__or2b_1 _15608_ (.A(_08673_),
    .B_N(_08671_),
    .X(_08683_));
 sky130_fd_sc_hd__or2b_1 _15609_ (.A(_08674_),
    .B_N(_08670_),
    .X(_08684_));
 sky130_fd_sc_hd__nand2_2 _15610_ (.A(_08683_),
    .B(_08684_),
    .Y(_08685_));
 sky130_fd_sc_hd__o21ai_2 _15611_ (.A1(_08127_),
    .A2(_08598_),
    .B1(_08345_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand2_1 _15612_ (.A(_08346_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__xnor2_2 _15613_ (.A(_08685_),
    .B(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__xnor2_1 _15614_ (.A(_08682_),
    .B(_08688_),
    .Y(_08689_));
 sky130_fd_sc_hd__nor2_1 _15615_ (.A(_08645_),
    .B(_08677_),
    .Y(_08690_));
 sky130_fd_sc_hd__a21oi_1 _15616_ (.A1(_08678_),
    .A2(_08689_),
    .B1(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__xnor2_2 _15617_ (.A(_08644_),
    .B(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__nor2_1 _15618_ (.A(_08343_),
    .B(_08681_),
    .Y(_08693_));
 sky130_fd_sc_hd__and3_1 _15619_ (.A(_08338_),
    .B(_08679_),
    .C(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__a32oi_4 _15620_ (.A1(_08346_),
    .A2(_08685_),
    .A3(_08686_),
    .B1(_08688_),
    .B2(_08694_),
    .Y(_08695_));
 sky130_fd_sc_hd__xnor2_2 _15621_ (.A(_08692_),
    .B(_08695_),
    .Y(_08696_));
 sky130_fd_sc_hd__xnor2_1 _15622_ (.A(_08665_),
    .B(_08668_),
    .Y(_08697_));
 sky130_fd_sc_hd__or3_1 _15623_ (.A(_08190_),
    .B(_08224_),
    .C(_08228_),
    .X(_08698_));
 sky130_fd_sc_hd__xor2_1 _15624_ (.A(_08655_),
    .B(_08698_),
    .X(_08699_));
 sky130_fd_sc_hd__nor2_1 _15625_ (.A(_08204_),
    .B(_08255_),
    .Y(_08700_));
 sky130_fd_sc_hd__a2bb2o_1 _15626_ (.A1_N(_08655_),
    .A2_N(_08698_),
    .B1(_08699_),
    .B2(_08700_),
    .X(_08701_));
 sky130_fd_sc_hd__or2b_1 _15627_ (.A(_08697_),
    .B_N(_08701_),
    .X(_08702_));
 sky130_fd_sc_hd__xor2_1 _15628_ (.A(_08701_),
    .B(_08697_),
    .X(_08703_));
 sky130_fd_sc_hd__or3_1 _15629_ (.A(_08222_),
    .B(_08242_),
    .C(_08316_),
    .X(_08704_));
 sky130_fd_sc_hd__nor2_1 _15630_ (.A(_08266_),
    .B(_08326_),
    .Y(_08705_));
 sky130_fd_sc_hd__o32a_1 _15631_ (.A1(_08222_),
    .A2(_08274_),
    .A3(_08278_),
    .B1(_08316_),
    .B2(_08243_),
    .X(_08706_));
 sky130_fd_sc_hd__o21ba_1 _15632_ (.A1(_08279_),
    .A2(_08704_),
    .B1_N(_08706_),
    .X(_08707_));
 sky130_fd_sc_hd__nand2_1 _15633_ (.A(_08705_),
    .B(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__o21ai_1 _15634_ (.A1(_08280_),
    .A2(_08704_),
    .B1(_08708_),
    .Y(_08709_));
 sky130_fd_sc_hd__or2b_1 _15635_ (.A(_08703_),
    .B_N(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__o21ai_1 _15636_ (.A1(_08343_),
    .A2(_08681_),
    .B1(_08680_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_1 _15637_ (.A(_08682_),
    .B(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__a21oi_2 _15638_ (.A1(_08702_),
    .A2(_08710_),
    .B1(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__xnor2_1 _15639_ (.A(_08678_),
    .B(_08689_),
    .Y(_08714_));
 sky130_fd_sc_hd__xnor2_1 _15640_ (.A(_08664_),
    .B(_08675_),
    .Y(_08715_));
 sky130_fd_sc_hd__a21o_1 _15641_ (.A1(_08653_),
    .A2(_08661_),
    .B1(_08660_),
    .X(_08716_));
 sky130_fd_sc_hd__a2bb2o_1 _15642_ (.A1_N(_08177_),
    .A2_N(_08419_),
    .B1(_08648_),
    .B2(_08650_),
    .X(_08717_));
 sky130_fd_sc_hd__o22ai_2 _15643_ (.A1(_08649_),
    .A2(_08436_),
    .B1(_08480_),
    .B2(_08176_),
    .Y(_08718_));
 sky130_fd_sc_hd__and4bb_1 _15644_ (.A_N(_08649_),
    .B_N(_08176_),
    .C(_08468_),
    .D(_08439_),
    .X(_08719_));
 sky130_fd_sc_hd__a31o_1 _15645_ (.A1(_08497_),
    .A2(_08457_),
    .A3(_08718_),
    .B1(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__nand3_1 _15646_ (.A(_08651_),
    .B(_08717_),
    .C(_08720_),
    .Y(_08721_));
 sky130_fd_sc_hd__xor2_1 _15647_ (.A(_08700_),
    .B(_08699_),
    .X(_08722_));
 sky130_fd_sc_hd__a21o_1 _15648_ (.A1(_08651_),
    .A2(_08717_),
    .B1(_08720_),
    .X(_08723_));
 sky130_fd_sc_hd__nand3_1 _15649_ (.A(_08721_),
    .B(_08722_),
    .C(_08723_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand2_1 _15650_ (.A(_08721_),
    .B(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__nand3_1 _15651_ (.A(_08662_),
    .B(_08716_),
    .C(_08725_),
    .Y(_08726_));
 sky130_fd_sc_hd__xnor2_1 _15652_ (.A(_08709_),
    .B(_08703_),
    .Y(_08727_));
 sky130_fd_sc_hd__a21o_1 _15653_ (.A1(_08662_),
    .A2(_08716_),
    .B1(_08725_),
    .X(_08728_));
 sky130_fd_sc_hd__nand3_1 _15654_ (.A(_08726_),
    .B(_08727_),
    .C(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__and2_1 _15655_ (.A(_08726_),
    .B(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__xor2_1 _15656_ (.A(_08715_),
    .B(_08730_),
    .X(_08731_));
 sky130_fd_sc_hd__and3_1 _15657_ (.A(_08702_),
    .B(_08710_),
    .C(_08712_),
    .X(_08732_));
 sky130_fd_sc_hd__nor2_1 _15658_ (.A(_08713_),
    .B(_08732_),
    .Y(_08733_));
 sky130_fd_sc_hd__nor2_1 _15659_ (.A(_08715_),
    .B(_08730_),
    .Y(_08734_));
 sky130_fd_sc_hd__a21o_1 _15660_ (.A1(_08731_),
    .A2(_08733_),
    .B1(_08734_),
    .X(_08735_));
 sky130_fd_sc_hd__xnor2_1 _15661_ (.A(_08714_),
    .B(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__or2b_1 _15662_ (.A(_08714_),
    .B_N(_08735_),
    .X(_08737_));
 sky130_fd_sc_hd__a21boi_2 _15663_ (.A1(_08713_),
    .A2(_08736_),
    .B1_N(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__nor2_1 _15664_ (.A(_08696_),
    .B(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__inv_2 _15665_ (.A(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__xnor2_1 _15666_ (.A(_08637_),
    .B(_08639_),
    .Y(_08741_));
 sky130_fd_sc_hd__or2_1 _15667_ (.A(_08644_),
    .B(_08691_),
    .X(_08742_));
 sky130_fd_sc_hd__o21a_1 _15668_ (.A1(_08692_),
    .A2(_08695_),
    .B1(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__nor2_1 _15669_ (.A(_08741_),
    .B(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__and2_1 _15670_ (.A(_08741_),
    .B(_08743_),
    .X(_08745_));
 sky130_fd_sc_hd__or2_1 _15671_ (.A(_08744_),
    .B(_08745_),
    .X(_08746_));
 sky130_fd_sc_hd__nor2_1 _15672_ (.A(_08740_),
    .B(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__xnor2_1 _15673_ (.A(_08713_),
    .B(_08736_),
    .Y(_08748_));
 sky130_fd_sc_hd__nor2_1 _15674_ (.A(_08204_),
    .B(_08280_),
    .Y(_08749_));
 sky130_fd_sc_hd__or3_1 _15675_ (.A(_08170_),
    .B(_08224_),
    .C(_08245_),
    .X(_08750_));
 sky130_fd_sc_hd__o2111a_1 _15676_ (.A1(\rbzero.wall_tracer.stepDistY[-7] ),
    .A2(_08144_),
    .B1(_08657_),
    .C1(_08250_),
    .D1(_08253_),
    .X(_08751_));
 sky130_fd_sc_hd__xnor2_1 _15677_ (.A(_08750_),
    .B(_08751_),
    .Y(_08752_));
 sky130_fd_sc_hd__or3_1 _15678_ (.A(_08171_),
    .B(_08254_),
    .C(_08698_),
    .X(_08753_));
 sky130_fd_sc_hd__a21boi_1 _15679_ (.A1(_08749_),
    .A2(_08752_),
    .B1_N(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__xnor2_1 _15680_ (.A(_08705_),
    .B(_08707_),
    .Y(_08755_));
 sky130_fd_sc_hd__or2_1 _15681_ (.A(_08754_),
    .B(_08755_),
    .X(_08756_));
 sky130_fd_sc_hd__xnor2_1 _15682_ (.A(_08754_),
    .B(_08755_),
    .Y(_08757_));
 sky130_fd_sc_hd__o221ai_4 _15683_ (.A1(\rbzero.wall_tracer.stepDistX[-10] ),
    .A2(_08130_),
    .B1(_08145_),
    .B2(_08146_),
    .C1(_08247_),
    .Y(_08758_));
 sky130_fd_sc_hd__nor2_1 _15684_ (.A(_08223_),
    .B(_08316_),
    .Y(_08759_));
 sky130_fd_sc_hd__xnor2_1 _15685_ (.A(_08759_),
    .B(_08758_),
    .Y(_08760_));
 sky130_fd_sc_hd__or3b_1 _15686_ (.A(_08267_),
    .B(_08340_),
    .C_N(_08760_),
    .X(_08761_));
 sky130_fd_sc_hd__o31ai_2 _15687_ (.A1(_08352_),
    .A2(_08317_),
    .A3(_08758_),
    .B1(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__or2b_1 _15688_ (.A(_08757_),
    .B_N(_08762_),
    .X(_08763_));
 sky130_fd_sc_hd__or2_1 _15689_ (.A(_08338_),
    .B(_08679_),
    .X(_08764_));
 sky130_fd_sc_hd__nand2_1 _15690_ (.A(_08680_),
    .B(_08764_),
    .Y(_08765_));
 sky130_fd_sc_hd__a21oi_2 _15691_ (.A1(_08756_),
    .A2(_08763_),
    .B1(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__xnor2_1 _15692_ (.A(_08731_),
    .B(_08733_),
    .Y(_08767_));
 sky130_fd_sc_hd__a21o_1 _15693_ (.A1(_08726_),
    .A2(_08728_),
    .B1(_08727_),
    .X(_08768_));
 sky130_fd_sc_hd__a21o_1 _15694_ (.A1(_08721_),
    .A2(_08723_),
    .B1(_08722_),
    .X(_08769_));
 sky130_fd_sc_hd__xor2_1 _15695_ (.A(_08749_),
    .B(_08752_),
    .X(_08770_));
 sky130_fd_sc_hd__or4b_1 _15696_ (.A(_08211_),
    .B(_08419_),
    .C(_08719_),
    .D_N(_08718_),
    .X(_08771_));
 sky130_fd_sc_hd__or4_1 _15697_ (.A(_08649_),
    .B(_08176_),
    .C(_08436_),
    .D(_08480_),
    .X(_08772_));
 sky130_fd_sc_hd__a22o_1 _15698_ (.A1(_08497_),
    .A2(_08457_),
    .B1(_08772_),
    .B2(_08718_),
    .X(_08773_));
 sky130_fd_sc_hd__o22ai_1 _15699_ (.A1(_08176_),
    .A2(_08436_),
    .B1(_08480_),
    .B2(_08209_),
    .Y(_08774_));
 sky130_fd_sc_hd__and4bb_1 _15700_ (.A_N(_08176_),
    .B_N(_08209_),
    .C(_08468_),
    .D(_08439_),
    .X(_08775_));
 sky130_fd_sc_hd__a31o_1 _15701_ (.A1(_08246_),
    .A2(_08457_),
    .A3(_08774_),
    .B1(_08775_),
    .X(_08776_));
 sky130_fd_sc_hd__a21o_1 _15702_ (.A1(_08771_),
    .A2(_08773_),
    .B1(_08776_),
    .X(_08777_));
 sky130_fd_sc_hd__and3_1 _15703_ (.A(_08771_),
    .B(_08773_),
    .C(_08776_),
    .X(_08778_));
 sky130_fd_sc_hd__a21o_1 _15704_ (.A1(_08770_),
    .A2(_08777_),
    .B1(_08778_),
    .X(_08779_));
 sky130_fd_sc_hd__nand3_1 _15705_ (.A(_08724_),
    .B(_08769_),
    .C(_08779_),
    .Y(_08780_));
 sky130_fd_sc_hd__xnor2_1 _15706_ (.A(_08762_),
    .B(_08757_),
    .Y(_08781_));
 sky130_fd_sc_hd__a21o_1 _15707_ (.A1(_08724_),
    .A2(_08769_),
    .B1(_08779_),
    .X(_08782_));
 sky130_fd_sc_hd__nand3_1 _15708_ (.A(_08780_),
    .B(_08781_),
    .C(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__nand2_1 _15709_ (.A(_08780_),
    .B(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__a21o_1 _15710_ (.A1(_08729_),
    .A2(_08768_),
    .B1(_08784_),
    .X(_08785_));
 sky130_fd_sc_hd__and3_1 _15711_ (.A(_08756_),
    .B(_08763_),
    .C(_08765_),
    .X(_08786_));
 sky130_fd_sc_hd__nor2_1 _15712_ (.A(_08766_),
    .B(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__nand3_1 _15713_ (.A(_08729_),
    .B(_08768_),
    .C(_08784_),
    .Y(_08788_));
 sky130_fd_sc_hd__a21boi_1 _15714_ (.A1(_08785_),
    .A2(_08787_),
    .B1_N(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__xor2_1 _15715_ (.A(_08767_),
    .B(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__nor2_1 _15716_ (.A(_08767_),
    .B(_08789_),
    .Y(_08791_));
 sky130_fd_sc_hd__a21oi_1 _15717_ (.A1(_08766_),
    .A2(_08790_),
    .B1(_08791_),
    .Y(_08792_));
 sky130_fd_sc_hd__nor2_1 _15718_ (.A(_08748_),
    .B(_08792_),
    .Y(_08793_));
 sky130_fd_sc_hd__xor2_2 _15719_ (.A(_08696_),
    .B(_08738_),
    .X(_08794_));
 sky130_fd_sc_hd__nand2_1 _15720_ (.A(_08793_),
    .B(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__xnor2_1 _15721_ (.A(_08766_),
    .B(_08790_),
    .Y(_08796_));
 sky130_fd_sc_hd__clkbuf_4 _15722_ (.A(_08296_),
    .X(_08797_));
 sky130_fd_sc_hd__clkbuf_4 _15723_ (.A(_08797_),
    .X(_08798_));
 sky130_fd_sc_hd__or2_1 _15724_ (.A(_08798_),
    .B(_08341_),
    .X(_08799_));
 sky130_fd_sc_hd__nor2_1 _15725_ (.A(_08171_),
    .B(_08255_),
    .Y(_08800_));
 sky130_fd_sc_hd__nor2_1 _15726_ (.A(_08191_),
    .B(_08280_),
    .Y(_08801_));
 sky130_fd_sc_hd__xnor2_1 _15727_ (.A(_08800_),
    .B(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__or2_1 _15728_ (.A(_08204_),
    .B(_08317_),
    .X(_08803_));
 sky130_fd_sc_hd__o2bb2ai_1 _15729_ (.A1_N(_08800_),
    .A2_N(_08801_),
    .B1(_08802_),
    .B2(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__or2_1 _15730_ (.A(_08267_),
    .B(_08340_),
    .X(_08805_));
 sky130_fd_sc_hd__xnor2_1 _15731_ (.A(_08805_),
    .B(_08760_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand2_1 _15732_ (.A(_08804_),
    .B(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__or2_1 _15733_ (.A(_08804_),
    .B(_08806_),
    .X(_08808_));
 sky130_fd_sc_hd__nand2_1 _15734_ (.A(_08807_),
    .B(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__or2_1 _15735_ (.A(_08223_),
    .B(_08341_),
    .X(_08810_));
 sky130_fd_sc_hd__clkbuf_2 _15736_ (.A(_08810_),
    .X(_08811_));
 sky130_fd_sc_hd__o31a_1 _15737_ (.A1(_08758_),
    .A2(_08809_),
    .A3(_08811_),
    .B1(_08807_),
    .X(_08812_));
 sky130_fd_sc_hd__nor2_1 _15738_ (.A(_08799_),
    .B(_08812_),
    .Y(_08813_));
 sky130_fd_sc_hd__and3_1 _15739_ (.A(_08788_),
    .B(_08785_),
    .C(_08787_),
    .X(_08814_));
 sky130_fd_sc_hd__a21oi_1 _15740_ (.A1(_08788_),
    .A2(_08785_),
    .B1(_08787_),
    .Y(_08815_));
 sky130_fd_sc_hd__or2_1 _15741_ (.A(_08814_),
    .B(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__and2_1 _15742_ (.A(_08799_),
    .B(_08812_),
    .X(_08817_));
 sky130_fd_sc_hd__nor2_1 _15743_ (.A(_08813_),
    .B(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__a21o_1 _15744_ (.A1(_08780_),
    .A2(_08782_),
    .B1(_08781_),
    .X(_08819_));
 sky130_fd_sc_hd__nand2_1 _15745_ (.A(_08783_),
    .B(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__nor2_1 _15746_ (.A(_08758_),
    .B(_08811_),
    .Y(_08821_));
 sky130_fd_sc_hd__xnor2_1 _15747_ (.A(_08809_),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__and2b_1 _15748_ (.A_N(_08778_),
    .B(_08777_),
    .X(_08823_));
 sky130_fd_sc_hd__xnor2_1 _15749_ (.A(_08770_),
    .B(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__xor2_1 _15750_ (.A(_08803_),
    .B(_08802_),
    .X(_08825_));
 sky130_fd_sc_hd__nor2_1 _15751_ (.A(_08230_),
    .B(_08419_),
    .Y(_08826_));
 sky130_fd_sc_hd__and2b_1 _15752_ (.A_N(_08775_),
    .B(_08774_),
    .X(_08827_));
 sky130_fd_sc_hd__xnor2_1 _15753_ (.A(_08826_),
    .B(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__nor2_1 _15754_ (.A(_08209_),
    .B(_08437_),
    .Y(_08829_));
 sky130_fd_sc_hd__clkbuf_4 _15755_ (.A(_08480_),
    .X(_08830_));
 sky130_fd_sc_hd__nor2_1 _15756_ (.A(_08245_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__nor2_1 _15757_ (.A(_08829_),
    .B(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__or4_1 _15758_ (.A(_08209_),
    .B(_08245_),
    .C(_08437_),
    .D(_08480_),
    .X(_08833_));
 sky130_fd_sc_hd__o31a_1 _15759_ (.A1(_08255_),
    .A2(_08420_),
    .A3(_08832_),
    .B1(_08833_),
    .X(_08834_));
 sky130_fd_sc_hd__xor2_1 _15760_ (.A(_08828_),
    .B(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__nor2_1 _15761_ (.A(_08828_),
    .B(_08834_),
    .Y(_08836_));
 sky130_fd_sc_hd__a21oi_1 _15762_ (.A1(_08825_),
    .A2(_08835_),
    .B1(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__nor2_1 _15763_ (.A(_08824_),
    .B(_08837_),
    .Y(_08838_));
 sky130_fd_sc_hd__and2_1 _15764_ (.A(_08824_),
    .B(_08837_),
    .X(_08839_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(_08838_),
    .B(_08839_),
    .Y(_08840_));
 sky130_fd_sc_hd__a21o_1 _15766_ (.A1(_08822_),
    .A2(_08840_),
    .B1(_08838_),
    .X(_08841_));
 sky130_fd_sc_hd__xnor2_1 _15767_ (.A(_08820_),
    .B(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__and3_1 _15768_ (.A(_08783_),
    .B(_08819_),
    .C(_08841_),
    .X(_08843_));
 sky130_fd_sc_hd__a21oi_1 _15769_ (.A1(_08818_),
    .A2(_08842_),
    .B1(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__xor2_1 _15770_ (.A(_08816_),
    .B(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _15771_ (.A(_08816_),
    .B(_08844_),
    .Y(_08846_));
 sky130_fd_sc_hd__a21oi_1 _15772_ (.A1(_08813_),
    .A2(_08845_),
    .B1(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__nor2_1 _15773_ (.A(_08796_),
    .B(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__xor2_1 _15774_ (.A(_08748_),
    .B(_08792_),
    .X(_08849_));
 sky130_fd_sc_hd__and2_1 _15775_ (.A(_08848_),
    .B(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__xor2_1 _15776_ (.A(_08796_),
    .B(_08847_),
    .X(_08851_));
 sky130_fd_sc_hd__xnor2_1 _15777_ (.A(_08813_),
    .B(_08845_),
    .Y(_08852_));
 sky130_fd_sc_hd__xnor2_1 _15778_ (.A(_08822_),
    .B(_08840_),
    .Y(_08853_));
 sky130_fd_sc_hd__xnor2_1 _15779_ (.A(_08825_),
    .B(_08835_),
    .Y(_08854_));
 sky130_fd_sc_hd__nor2_1 _15780_ (.A(_08255_),
    .B(_08420_),
    .Y(_08855_));
 sky130_fd_sc_hd__o21a_1 _15781_ (.A1(_08829_),
    .A2(_08831_),
    .B1(_08833_),
    .X(_08856_));
 sky130_fd_sc_hd__xnor2_1 _15782_ (.A(_08855_),
    .B(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__or2_1 _15783_ (.A(_08280_),
    .B(_08420_),
    .X(_08858_));
 sky130_fd_sc_hd__o22a_1 _15784_ (.A1(_08245_),
    .A2(_08437_),
    .B1(_08830_),
    .B2(_08511_),
    .X(_08859_));
 sky130_fd_sc_hd__clkbuf_4 _15785_ (.A(_08511_),
    .X(_08860_));
 sky130_fd_sc_hd__or3b_1 _15786_ (.A(_08860_),
    .B(_08437_),
    .C_N(_08831_),
    .X(_08861_));
 sky130_fd_sc_hd__o21a_1 _15787_ (.A1(_08858_),
    .A2(_08859_),
    .B1(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__nor2_1 _15788_ (.A(_08857_),
    .B(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__and2_1 _15789_ (.A(_08857_),
    .B(_08862_),
    .X(_08864_));
 sky130_fd_sc_hd__nor2_1 _15790_ (.A(_08863_),
    .B(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__buf_2 _15791_ (.A(_08326_),
    .X(_08866_));
 sky130_fd_sc_hd__or2_1 _15792_ (.A(_08359_),
    .B(_08866_),
    .X(_08867_));
 sky130_fd_sc_hd__or2_1 _15793_ (.A(_08171_),
    .B(_08280_),
    .X(_08868_));
 sky130_fd_sc_hd__or2_2 _15794_ (.A(_08191_),
    .B(_08317_),
    .X(_08869_));
 sky130_fd_sc_hd__xnor2_1 _15795_ (.A(_08868_),
    .B(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__xor2_1 _15796_ (.A(_08867_),
    .B(_08870_),
    .X(_08871_));
 sky130_fd_sc_hd__a21oi_1 _15797_ (.A1(_08865_),
    .A2(_08871_),
    .B1(_08863_),
    .Y(_08872_));
 sky130_fd_sc_hd__nand2_1 _15798_ (.A(_08854_),
    .B(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__o22ai_2 _15799_ (.A1(_08868_),
    .A2(_08869_),
    .B1(_08870_),
    .B2(_08867_),
    .Y(_08874_));
 sky130_fd_sc_hd__clkbuf_4 _15800_ (.A(_08352_),
    .X(_08875_));
 sky130_fd_sc_hd__buf_4 _15801_ (.A(_08243_),
    .X(_08876_));
 sky130_fd_sc_hd__o22a_1 _15802_ (.A1(_08875_),
    .A2(_08866_),
    .B1(_08341_),
    .B2(_08876_),
    .X(_08877_));
 sky130_fd_sc_hd__or2_1 _15803_ (.A(_08821_),
    .B(_08877_),
    .X(_08878_));
 sky130_fd_sc_hd__xnor2_1 _15804_ (.A(_08874_),
    .B(_08878_),
    .Y(_08879_));
 sky130_fd_sc_hd__nor2_1 _15805_ (.A(_08854_),
    .B(_08872_),
    .Y(_08880_));
 sky130_fd_sc_hd__a21oi_1 _15806_ (.A1(_08873_),
    .A2(_08879_),
    .B1(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__or2_1 _15807_ (.A(_08853_),
    .B(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__and2b_1 _15808_ (.A_N(_08878_),
    .B(_08874_),
    .X(_08883_));
 sky130_fd_sc_hd__nand2_1 _15809_ (.A(_08853_),
    .B(_08881_),
    .Y(_08884_));
 sky130_fd_sc_hd__and2_1 _15810_ (.A(_08882_),
    .B(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__nand2_1 _15811_ (.A(_08883_),
    .B(_08885_),
    .Y(_08886_));
 sky130_fd_sc_hd__xnor2_1 _15812_ (.A(_08818_),
    .B(_08842_),
    .Y(_08887_));
 sky130_fd_sc_hd__a21o_1 _15813_ (.A1(_08882_),
    .A2(_08886_),
    .B1(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__nor2_1 _15814_ (.A(_08852_),
    .B(_08888_),
    .Y(_08889_));
 sky130_fd_sc_hd__and2_1 _15815_ (.A(_08851_),
    .B(_08889_),
    .X(_08890_));
 sky130_fd_sc_hd__xnor2_1 _15816_ (.A(_08851_),
    .B(_08889_),
    .Y(_08891_));
 sky130_fd_sc_hd__nand2_1 _15817_ (.A(_08887_),
    .B(_08882_),
    .Y(_08892_));
 sky130_fd_sc_hd__and2b_1 _15818_ (.A_N(_08880_),
    .B(_08873_),
    .X(_08893_));
 sky130_fd_sc_hd__xnor2_1 _15819_ (.A(_08893_),
    .B(_08879_),
    .Y(_08894_));
 sky130_fd_sc_hd__xnor2_1 _15820_ (.A(_08865_),
    .B(_08871_),
    .Y(_08895_));
 sky130_fd_sc_hd__or2_1 _15821_ (.A(_08359_),
    .B(_08341_),
    .X(_08896_));
 sky130_fd_sc_hd__o22ai_1 _15822_ (.A1(_08412_),
    .A2(_08317_),
    .B1(_08866_),
    .B2(_08399_),
    .Y(_08897_));
 sky130_fd_sc_hd__o31a_1 _15823_ (.A1(_08412_),
    .A2(_08866_),
    .A3(_08869_),
    .B1(_08897_),
    .X(_08898_));
 sky130_fd_sc_hd__xnor2_1 _15824_ (.A(_08896_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__a31o_1 _15825_ (.A1(_08512_),
    .A2(_08468_),
    .A3(_08831_),
    .B1(_08859_),
    .X(_08900_));
 sky130_fd_sc_hd__xnor2_1 _15826_ (.A(_08858_),
    .B(_08900_),
    .Y(_08901_));
 sky130_fd_sc_hd__o22a_1 _15827_ (.A1(_08860_),
    .A2(_08437_),
    .B1(_08830_),
    .B2(_08278_),
    .X(_08902_));
 sky130_fd_sc_hd__or2_1 _15828_ (.A(_08278_),
    .B(_08437_),
    .X(_08903_));
 sky130_fd_sc_hd__or3_1 _15829_ (.A(_08860_),
    .B(_08830_),
    .C(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__o31a_1 _15830_ (.A1(_08317_),
    .A2(_08420_),
    .A3(_08902_),
    .B1(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__nor2_1 _15831_ (.A(_08901_),
    .B(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__and2_1 _15832_ (.A(_08901_),
    .B(_08905_),
    .X(_08907_));
 sky130_fd_sc_hd__nor2_1 _15833_ (.A(_08906_),
    .B(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__a21oi_1 _15834_ (.A1(_08899_),
    .A2(_08908_),
    .B1(_08906_),
    .Y(_08909_));
 sky130_fd_sc_hd__xor2_1 _15835_ (.A(_08895_),
    .B(_08909_),
    .X(_08910_));
 sky130_fd_sc_hd__clkbuf_4 _15836_ (.A(_08412_),
    .X(_08911_));
 sky130_fd_sc_hd__or2b_1 _15837_ (.A(_08896_),
    .B_N(_08898_),
    .X(_08912_));
 sky130_fd_sc_hd__o31a_1 _15838_ (.A1(_08911_),
    .A2(_08866_),
    .A3(_08869_),
    .B1(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__xor2_1 _15839_ (.A(_08811_),
    .B(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__nand2_1 _15840_ (.A(_08910_),
    .B(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__o21a_1 _15841_ (.A1(_08895_),
    .A2(_08909_),
    .B1(_08915_),
    .X(_08916_));
 sky130_fd_sc_hd__or2_1 _15842_ (.A(_08894_),
    .B(_08916_),
    .X(_08917_));
 sky130_fd_sc_hd__xnor2_1 _15843_ (.A(_08894_),
    .B(_08916_),
    .Y(_08918_));
 sky130_fd_sc_hd__or3_1 _15844_ (.A(_08811_),
    .B(_08913_),
    .C(_08918_),
    .X(_08919_));
 sky130_fd_sc_hd__or2_1 _15845_ (.A(_08883_),
    .B(_08885_),
    .X(_08920_));
 sky130_fd_sc_hd__nand2_1 _15846_ (.A(_08886_),
    .B(_08920_),
    .Y(_08921_));
 sky130_fd_sc_hd__a211oi_1 _15847_ (.A1(_08917_),
    .A2(_08919_),
    .B1(_08852_),
    .C1(_08921_),
    .Y(_08922_));
 sky130_fd_sc_hd__and3_1 _15848_ (.A(_08888_),
    .B(_08892_),
    .C(_08922_),
    .X(_08923_));
 sky130_fd_sc_hd__xnor2_1 _15849_ (.A(_08891_),
    .B(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__or2_1 _15850_ (.A(_08910_),
    .B(_08914_),
    .X(_08925_));
 sky130_fd_sc_hd__nand2_1 _15851_ (.A(_08915_),
    .B(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__xnor2_1 _15852_ (.A(_08899_),
    .B(_08908_),
    .Y(_08927_));
 sky130_fd_sc_hd__clkbuf_4 _15853_ (.A(_08420_),
    .X(_08928_));
 sky130_fd_sc_hd__nor2_1 _15854_ (.A(_08317_),
    .B(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__inv_2 _15855_ (.A(_08904_),
    .Y(_08930_));
 sky130_fd_sc_hd__nor2_1 _15856_ (.A(_08930_),
    .B(_08902_),
    .Y(_08931_));
 sky130_fd_sc_hd__xnor2_1 _15857_ (.A(_08929_),
    .B(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__or2_1 _15858_ (.A(_08866_),
    .B(_08928_),
    .X(_08933_));
 sky130_fd_sc_hd__o21a_1 _15859_ (.A1(_08520_),
    .A2(_08830_),
    .B1(_08903_),
    .X(_08934_));
 sky130_fd_sc_hd__clkbuf_4 _15860_ (.A(_08278_),
    .X(_08935_));
 sky130_fd_sc_hd__nor2_1 _15861_ (.A(_08520_),
    .B(_08437_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand2_1 _15862_ (.A(_08439_),
    .B(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__or2_1 _15863_ (.A(_08935_),
    .B(_08937_),
    .X(_08938_));
 sky130_fd_sc_hd__o21a_1 _15864_ (.A1(_08933_),
    .A2(_08934_),
    .B1(_08938_),
    .X(_08939_));
 sky130_fd_sc_hd__nand2_1 _15865_ (.A(_08932_),
    .B(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__clkbuf_4 _15866_ (.A(_08399_),
    .X(_08941_));
 sky130_fd_sc_hd__or2_1 _15867_ (.A(_08911_),
    .B(_08341_),
    .X(_08942_));
 sky130_fd_sc_hd__o22ai_1 _15868_ (.A1(_08911_),
    .A2(_08866_),
    .B1(_08341_),
    .B2(_08941_),
    .Y(_08943_));
 sky130_fd_sc_hd__o31a_1 _15869_ (.A1(_08941_),
    .A2(_08866_),
    .A3(_08942_),
    .B1(_08943_),
    .X(_08944_));
 sky130_fd_sc_hd__nor2_1 _15870_ (.A(_08932_),
    .B(_08939_),
    .Y(_08945_));
 sky130_fd_sc_hd__a21oi_1 _15871_ (.A1(_08940_),
    .A2(_08944_),
    .B1(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__xnor2_1 _15872_ (.A(_08927_),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__or4_1 _15873_ (.A(_08941_),
    .B(_08866_),
    .C(_08942_),
    .D(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__o21a_1 _15874_ (.A1(_08927_),
    .A2(_08946_),
    .B1(_08948_),
    .X(_08949_));
 sky130_fd_sc_hd__and2b_1 _15875_ (.A_N(_08945_),
    .B(_08940_),
    .X(_08950_));
 sky130_fd_sc_hd__xnor2_1 _15876_ (.A(_08950_),
    .B(_08944_),
    .Y(_08951_));
 sky130_fd_sc_hd__nor2_1 _15877_ (.A(_08147_),
    .B(_08830_),
    .Y(_08952_));
 sky130_fd_sc_hd__nor2_1 _15878_ (.A(_08341_),
    .B(_08928_),
    .Y(_08953_));
 sky130_fd_sc_hd__xor2_1 _15879_ (.A(_08936_),
    .B(_08952_),
    .X(_08954_));
 sky130_fd_sc_hd__and2_1 _15880_ (.A(_08953_),
    .B(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__a21o_1 _15881_ (.A1(_08936_),
    .A2(_08952_),
    .B1(_08955_),
    .X(_08956_));
 sky130_fd_sc_hd__o21ba_1 _15882_ (.A1(_08935_),
    .A2(_08937_),
    .B1_N(_08934_),
    .X(_08957_));
 sky130_fd_sc_hd__xnor2_1 _15883_ (.A(_08933_),
    .B(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__xnor2_1 _15884_ (.A(_08956_),
    .B(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__nor2_1 _15885_ (.A(_08942_),
    .B(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__a21oi_1 _15886_ (.A1(_08956_),
    .A2(_08958_),
    .B1(_08960_),
    .Y(_08961_));
 sky130_fd_sc_hd__a2bb2o_1 _15887_ (.A1_N(_08953_),
    .A2_N(_08954_),
    .B1(_08959_),
    .B2(_08942_),
    .X(_08962_));
 sky130_fd_sc_hd__or4b_1 _15888_ (.A(_08598_),
    .B(_08450_),
    .C(_08955_),
    .D_N(_08952_),
    .X(_08963_));
 sky130_fd_sc_hd__a211o_1 _15889_ (.A1(_08951_),
    .A2(_08961_),
    .B1(_08962_),
    .C1(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__o22a_1 _15890_ (.A1(_08951_),
    .A2(_08961_),
    .B1(_08964_),
    .B2(_08960_),
    .X(_08965_));
 sky130_fd_sc_hd__o31ai_1 _15891_ (.A1(_08941_),
    .A2(_08866_),
    .A3(_08942_),
    .B1(_08947_),
    .Y(_08966_));
 sky130_fd_sc_hd__nand2_1 _15892_ (.A(_08948_),
    .B(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__a211o_1 _15893_ (.A1(_08926_),
    .A2(_08949_),
    .B1(_08965_),
    .C1(_08967_),
    .X(_08968_));
 sky130_fd_sc_hd__o21a_1 _15894_ (.A1(_08926_),
    .A2(_08949_),
    .B1(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__o21ai_1 _15895_ (.A1(_08811_),
    .A2(_08913_),
    .B1(_08918_),
    .Y(_08970_));
 sky130_fd_sc_hd__and4b_1 _15896_ (.A_N(_08969_),
    .B(_08970_),
    .C(_08919_),
    .D(_08888_),
    .X(_08971_));
 sky130_fd_sc_hd__or2b_1 _15897_ (.A(_08892_),
    .B_N(_08886_),
    .X(_08972_));
 sky130_fd_sc_hd__xor2_1 _15898_ (.A(_08921_),
    .B(_08917_),
    .X(_08973_));
 sky130_fd_sc_hd__and4b_1 _15899_ (.A_N(_08852_),
    .B(_08971_),
    .C(_08972_),
    .D(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__and2b_1 _15900_ (.A_N(_08891_),
    .B(_08923_),
    .X(_08975_));
 sky130_fd_sc_hd__a21o_1 _15901_ (.A1(_08924_),
    .A2(_08974_),
    .B1(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__nor2_1 _15902_ (.A(_08848_),
    .B(_08890_),
    .Y(_08977_));
 sky130_fd_sc_hd__xnor2_1 _15903_ (.A(_08849_),
    .B(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__a22o_2 _15904_ (.A1(_08849_),
    .A2(_08890_),
    .B1(_08976_),
    .B2(_08978_),
    .X(_08979_));
 sky130_fd_sc_hd__nor2_1 _15905_ (.A(_08793_),
    .B(_08850_),
    .Y(_08980_));
 sky130_fd_sc_hd__xnor2_2 _15906_ (.A(_08794_),
    .B(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__a22o_2 _15907_ (.A1(_08794_),
    .A2(_08850_),
    .B1(_08979_),
    .B2(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__nand2_1 _15908_ (.A(_08740_),
    .B(_08795_),
    .Y(_08983_));
 sky130_fd_sc_hd__xnor2_2 _15909_ (.A(_08746_),
    .B(_08983_),
    .Y(_08984_));
 sky130_fd_sc_hd__a2bb2o_2 _15910_ (.A1_N(_08746_),
    .A2_N(_08795_),
    .B1(_08982_),
    .B2(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__nor2_1 _15911_ (.A(_08744_),
    .B(_08747_),
    .Y(_08986_));
 sky130_fd_sc_hd__xnor2_2 _15912_ (.A(_08642_),
    .B(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__a22o_2 _15913_ (.A1(_08642_),
    .A2(_08747_),
    .B1(_08985_),
    .B2(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__a21o_1 _15914_ (.A1(_08540_),
    .A2(_08550_),
    .B1(_08548_),
    .X(_08989_));
 sky130_fd_sc_hd__or2b_1 _15915_ (.A(_08396_),
    .B_N(_08389_),
    .X(_08990_));
 sky130_fd_sc_hd__or2b_1 _15916_ (.A(_08397_),
    .B_N(_08358_),
    .X(_08991_));
 sky130_fd_sc_hd__or4_1 _15917_ (.A(_08125_),
    .B(_08148_),
    .C(_08860_),
    .D(_08278_),
    .X(_08992_));
 sky130_fd_sc_hd__o22ai_1 _15918_ (.A1(_08126_),
    .A2(_08860_),
    .B1(_08935_),
    .B2(_08148_),
    .Y(_08993_));
 sky130_fd_sc_hd__nand2_1 _15919_ (.A(_08992_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__or3_1 _15920_ (.A(_08602_),
    .B(_08534_),
    .C(_08994_),
    .X(_08995_));
 sky130_fd_sc_hd__o21ai_1 _15921_ (.A1(_08602_),
    .A2(_08534_),
    .B1(_08994_),
    .Y(_08996_));
 sky130_fd_sc_hd__and2_1 _15922_ (.A(_08995_),
    .B(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__nor2_1 _15923_ (.A(_08353_),
    .B(_08296_),
    .Y(_08998_));
 sky130_fd_sc_hd__xnor2_1 _15924_ (.A(_08541_),
    .B(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__or2_1 _15925_ (.A(_08230_),
    .B(_08546_),
    .X(_09000_));
 sky130_fd_sc_hd__xnor2_1 _15926_ (.A(_08999_),
    .B(_09000_),
    .Y(_09001_));
 sky130_fd_sc_hd__nand2_1 _15927_ (.A(_08514_),
    .B(_08541_),
    .Y(_09002_));
 sky130_fd_sc_hd__o31a_1 _15928_ (.A1(_08255_),
    .A2(_08546_),
    .A3(_08542_),
    .B1(_09002_),
    .X(_09003_));
 sky130_fd_sc_hd__nor2_1 _15929_ (.A(_09001_),
    .B(_09003_),
    .Y(_09004_));
 sky130_fd_sc_hd__and2_1 _15930_ (.A(_09001_),
    .B(_09003_),
    .X(_09005_));
 sky130_fd_sc_hd__nor2_1 _15931_ (.A(_09004_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__xnor2_1 _15932_ (.A(_08997_),
    .B(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__a21o_1 _15933_ (.A1(_08990_),
    .A2(_08991_),
    .B1(_09007_),
    .X(_09008_));
 sky130_fd_sc_hd__nand3_1 _15934_ (.A(_08990_),
    .B(_08991_),
    .C(_09007_),
    .Y(_09009_));
 sky130_fd_sc_hd__nand2_1 _15935_ (.A(_09008_),
    .B(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__xnor2_1 _15936_ (.A(_08989_),
    .B(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__a21bo_1 _15937_ (.A1(_08390_),
    .A2(_08391_),
    .B1_N(_08393_),
    .X(_09012_));
 sky130_fd_sc_hd__a22o_1 _15938_ (.A1(_08370_),
    .A2(_08410_),
    .B1(_08413_),
    .B2(_08415_),
    .X(_09013_));
 sky130_fd_sc_hd__nor2_1 _15939_ (.A(_08243_),
    .B(_08378_),
    .Y(_09014_));
 sky130_fd_sc_hd__o22ai_1 _15940_ (.A1(_08352_),
    .A2(_08378_),
    .B1(_08387_),
    .B2(_08243_),
    .Y(_09015_));
 sky130_fd_sc_hd__a21bo_1 _15941_ (.A1(_08391_),
    .A2(_09014_),
    .B1_N(_09015_),
    .X(_09016_));
 sky130_fd_sc_hd__nor2_1 _15942_ (.A(_08351_),
    .B(_08394_),
    .Y(_09017_));
 sky130_fd_sc_hd__xor2_2 _15943_ (.A(_09016_),
    .B(_09017_),
    .X(_09018_));
 sky130_fd_sc_hd__xnor2_2 _15944_ (.A(_09013_),
    .B(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__xor2_2 _15945_ (.A(_09012_),
    .B(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__nor2_2 _15946_ (.A(_08412_),
    .B(_08426_),
    .Y(_09021_));
 sky130_fd_sc_hd__xnor2_2 _15947_ (.A(_08410_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__nor2_1 _15948_ (.A(_08359_),
    .B(_08411_),
    .Y(_09023_));
 sky130_fd_sc_hd__xnor2_2 _15949_ (.A(_09022_),
    .B(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand2_4 _15950_ (.A(\rbzero.wall_tracer.stepDistX[3] ),
    .B(_06162_),
    .Y(_09025_));
 sky130_fd_sc_hd__nand2_1 _15951_ (.A(_08446_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__and2_1 _15952_ (.A(_08457_),
    .B(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__nand2_1 _15953_ (.A(_08439_),
    .B(_08444_),
    .Y(_09028_));
 sky130_fd_sc_hd__or3_1 _15954_ (.A(_07989_),
    .B(_07992_),
    .C(_08431_),
    .X(_09029_));
 sky130_fd_sc_hd__o21ai_1 _15955_ (.A1(_07989_),
    .A2(_08431_),
    .B1(_07992_),
    .Y(_09030_));
 sky130_fd_sc_hd__a31o_1 _15956_ (.A1(_08429_),
    .A2(_09029_),
    .A3(_09030_),
    .B1(_08434_),
    .X(_09031_));
 sky130_fd_sc_hd__nand2_1 _15957_ (.A(\rbzero.wall_tracer.stepDistY[5] ),
    .B(_08319_),
    .Y(_09032_));
 sky130_fd_sc_hd__a21oi_1 _15958_ (.A1(_09031_),
    .A2(_09032_),
    .B1(_06163_),
    .Y(_09033_));
 sky130_fd_sc_hd__nand2_1 _15959_ (.A(_08618_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__xor2_2 _15960_ (.A(_09028_),
    .B(_09034_),
    .X(_09035_));
 sky130_fd_sc_hd__xnor2_2 _15961_ (.A(_09027_),
    .B(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__or3_1 _15962_ (.A(_08450_),
    .B(_08446_),
    .C(_09028_),
    .X(_09037_));
 sky130_fd_sc_hd__o31a_1 _15963_ (.A1(_08928_),
    .A2(_08427_),
    .A3(_08451_),
    .B1(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__xor2_2 _15964_ (.A(_09036_),
    .B(_09038_),
    .X(_09039_));
 sky130_fd_sc_hd__xnor2_2 _15965_ (.A(_09024_),
    .B(_09039_),
    .Y(_09040_));
 sky130_fd_sc_hd__nor2_1 _15966_ (.A(_08453_),
    .B(_08461_),
    .Y(_09041_));
 sky130_fd_sc_hd__a21o_1 _15967_ (.A1(_08416_),
    .A2(_08462_),
    .B1(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__xnor2_1 _15968_ (.A(_09040_),
    .B(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__xnor2_2 _15969_ (.A(_09020_),
    .B(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__or2b_1 _15970_ (.A(_08463_),
    .B_N(_08474_),
    .X(_09045_));
 sky130_fd_sc_hd__a21boi_1 _15971_ (.A1(_08398_),
    .A2(_08475_),
    .B1_N(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__xor2_1 _15972_ (.A(_09044_),
    .B(_09046_),
    .X(_09047_));
 sky130_fd_sc_hd__xnor2_1 _15973_ (.A(_09011_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__and2b_1 _15974_ (.A_N(_08476_),
    .B(_08508_),
    .X(_09049_));
 sky130_fd_sc_hd__a21oi_1 _15975_ (.A1(_08509_),
    .A2(_08555_),
    .B1(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__nor2_1 _15976_ (.A(_09048_),
    .B(_09050_),
    .Y(_09051_));
 sky130_fd_sc_hd__nand2_1 _15977_ (.A(_09048_),
    .B(_09050_),
    .Y(_09052_));
 sky130_fd_sc_hd__and2b_1 _15978_ (.A_N(_09051_),
    .B(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__or2b_1 _15979_ (.A(_08554_),
    .B_N(_08531_),
    .X(_09054_));
 sky130_fd_sc_hd__nand2_4 _15980_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08124_),
    .Y(_09055_));
 sky130_fd_sc_hd__clkbuf_4 _15981_ (.A(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__or2_1 _15982_ (.A(_08147_),
    .B(_09056_),
    .X(_09057_));
 sky130_fd_sc_hd__nor2_1 _15983_ (.A(_08601_),
    .B(_09057_),
    .Y(_09058_));
 sky130_fd_sc_hd__o22a_1 _15984_ (.A1(_08285_),
    .A2(_08600_),
    .B1(_09056_),
    .B2(_08598_),
    .X(_09059_));
 sky130_fd_sc_hd__or2_1 _15985_ (.A(_09058_),
    .B(_09059_),
    .X(_09060_));
 sky130_fd_sc_hd__a21oi_1 _15986_ (.A1(_08536_),
    .A2(_08538_),
    .B1(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__and3_1 _15987_ (.A(_08536_),
    .B(_08538_),
    .C(_09060_),
    .X(_09062_));
 sky130_fd_sc_hd__nor2_1 _15988_ (.A(_09061_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_1 _15989_ (.A(_08604_),
    .B(_09063_),
    .Y(_09064_));
 sky130_fd_sc_hd__or2_1 _15990_ (.A(_08604_),
    .B(_09063_),
    .X(_09065_));
 sky130_fd_sc_hd__nand2_1 _15991_ (.A(_09064_),
    .B(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__a21oi_2 _15992_ (.A1(_08552_),
    .A2(_09054_),
    .B1(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__and3_1 _15993_ (.A(_08552_),
    .B(_09054_),
    .C(_09066_),
    .X(_09068_));
 sky130_fd_sc_hd__nor2_1 _15994_ (.A(_09067_),
    .B(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__xnor2_1 _15995_ (.A(_09053_),
    .B(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__nor2_1 _15996_ (.A(_08556_),
    .B(_08595_),
    .Y(_09071_));
 sky130_fd_sc_hd__a21oi_1 _15997_ (.A1(_08596_),
    .A2(_08609_),
    .B1(_09071_),
    .Y(_09072_));
 sky130_fd_sc_hd__xor2_1 _15998_ (.A(_09070_),
    .B(_09072_),
    .X(_09073_));
 sky130_fd_sc_hd__xnor2_1 _15999_ (.A(_08607_),
    .B(_09073_),
    .Y(_09074_));
 sky130_fd_sc_hd__or2b_1 _16000_ (.A(_08350_),
    .B_N(_08641_),
    .X(_09075_));
 sky130_fd_sc_hd__o21a_1 _16001_ (.A1(_08610_),
    .A2(_08640_),
    .B1(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__xor2_1 _16002_ (.A(_09074_),
    .B(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__and2_1 _16003_ (.A(_08642_),
    .B(_08744_),
    .X(_09078_));
 sky130_fd_sc_hd__nand2_1 _16004_ (.A(_09077_),
    .B(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__or2_1 _16005_ (.A(_09077_),
    .B(_09078_),
    .X(_09080_));
 sky130_fd_sc_hd__and2_2 _16006_ (.A(_09079_),
    .B(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__xor2_4 _16007_ (.A(_08988_),
    .B(_09081_),
    .X(_09082_));
 sky130_fd_sc_hd__and2b_1 _16008_ (.A_N(_08122_),
    .B(_09082_),
    .X(_09083_));
 sky130_fd_sc_hd__and2b_1 _16009_ (.A_N(_09082_),
    .B(_08122_),
    .X(_09084_));
 sky130_fd_sc_hd__nor2_1 _16010_ (.A(_09083_),
    .B(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__xor2_4 _16011_ (.A(_08985_),
    .B(_08987_),
    .X(_09086_));
 sky130_fd_sc_hd__mux2_1 _16012_ (.A0(\rbzero.debug_overlay.playerY[-7] ),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_04511_),
    .X(_09087_));
 sky130_fd_sc_hd__and2_1 _16013_ (.A(_09086_),
    .B(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__mux2_1 _16014_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_04511_),
    .X(_09089_));
 sky130_fd_sc_hd__xor2_4 _16015_ (.A(_08979_),
    .B(_08981_),
    .X(_09090_));
 sky130_fd_sc_hd__mux2_1 _16016_ (.A0(\rbzero.debug_overlay.playerY[-9] ),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_04511_),
    .X(_09091_));
 sky130_fd_sc_hd__and3_1 _16017_ (.A(_09089_),
    .B(_09090_),
    .C(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__xnor2_4 _16018_ (.A(_08982_),
    .B(_08984_),
    .Y(_09093_));
 sky130_fd_sc_hd__a21oi_1 _16019_ (.A1(_09090_),
    .A2(_09091_),
    .B1(_09089_),
    .Y(_09094_));
 sky130_fd_sc_hd__nor2_1 _16020_ (.A(_09093_),
    .B(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__or2_1 _16021_ (.A(_09086_),
    .B(_09087_),
    .X(_09096_));
 sky130_fd_sc_hd__o31a_1 _16022_ (.A1(_09088_),
    .A2(_09092_),
    .A3(_09095_),
    .B1(_09096_),
    .X(_09097_));
 sky130_fd_sc_hd__xnor2_1 _16023_ (.A(_09085_),
    .B(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__clkbuf_4 _16024_ (.A(_08178_),
    .X(_09099_));
 sky130_fd_sc_hd__clkbuf_4 _16025_ (.A(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__mux2_1 _16026_ (.A0(_09100_),
    .A1(_06076_),
    .S(_08115_),
    .X(_09101_));
 sky130_fd_sc_hd__buf_2 _16027_ (.A(_09101_),
    .X(_09102_));
 sky130_fd_sc_hd__nor2_1 _16028_ (.A(_09098_),
    .B(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__a211o_1 _16029_ (.A1(_09098_),
    .A2(_09102_),
    .B1(_09103_),
    .C1(_08429_),
    .X(_09104_));
 sky130_fd_sc_hd__o211a_1 _16030_ (.A1(\rbzero.texu_hot[0] ),
    .A2(_08120_),
    .B1(_09104_),
    .C1(_08059_),
    .X(_00466_));
 sky130_fd_sc_hd__a21bo_2 _16031_ (.A1(_08988_),
    .A2(_09081_),
    .B1_N(_09079_),
    .X(_09105_));
 sky130_fd_sc_hd__or2_2 _16032_ (.A(_09074_),
    .B(_09076_),
    .X(_09106_));
 sky130_fd_sc_hd__or2b_1 _16033_ (.A(_09010_),
    .B_N(_08989_),
    .X(_09107_));
 sky130_fd_sc_hd__nor2_1 _16034_ (.A(_08602_),
    .B(_08600_),
    .Y(_09108_));
 sky130_fd_sc_hd__xnor2_1 _16035_ (.A(_09057_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand2_4 _16036_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08523_),
    .Y(_09110_));
 sky130_fd_sc_hd__buf_4 _16037_ (.A(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__nor2_1 _16038_ (.A(_08598_),
    .B(_09111_),
    .Y(_09112_));
 sky130_fd_sc_hd__xnor2_1 _16039_ (.A(_09109_),
    .B(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__and3_1 _16040_ (.A(_08992_),
    .B(_08995_),
    .C(_09113_),
    .X(_09114_));
 sky130_fd_sc_hd__a21oi_1 _16041_ (.A1(_08992_),
    .A2(_08995_),
    .B1(_09113_),
    .Y(_09115_));
 sky130_fd_sc_hd__nor4_1 _16042_ (.A(_09058_),
    .B(_09061_),
    .C(_09114_),
    .D(_09115_),
    .Y(_09116_));
 sky130_fd_sc_hd__o22a_1 _16043_ (.A1(_09058_),
    .A2(_09061_),
    .B1(_09114_),
    .B2(_09115_),
    .X(_09117_));
 sky130_fd_sc_hd__nor2_1 _16044_ (.A(_09116_),
    .B(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__a21oi_1 _16045_ (.A1(_09008_),
    .A2(_09107_),
    .B1(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__and3_1 _16046_ (.A(_09008_),
    .B(_09107_),
    .C(_09118_),
    .X(_09120_));
 sky130_fd_sc_hd__nor2_1 _16047_ (.A(_09119_),
    .B(_09120_),
    .Y(_09121_));
 sky130_fd_sc_hd__xnor2_1 _16048_ (.A(_09064_),
    .B(_09121_),
    .Y(_09122_));
 sky130_fd_sc_hd__a21o_1 _16049_ (.A1(_08997_),
    .A2(_09006_),
    .B1(_09004_),
    .X(_09123_));
 sky130_fd_sc_hd__or2b_1 _16050_ (.A(_09018_),
    .B_N(_09013_),
    .X(_09124_));
 sky130_fd_sc_hd__nand2_1 _16051_ (.A(_09012_),
    .B(_09019_),
    .Y(_09125_));
 sky130_fd_sc_hd__or4_1 _16052_ (.A(_08125_),
    .B(_08148_),
    .C(_08245_),
    .D(_08860_),
    .X(_09126_));
 sky130_fd_sc_hd__clkbuf_4 _16053_ (.A(_08245_),
    .X(_09127_));
 sky130_fd_sc_hd__buf_2 _16054_ (.A(_08860_),
    .X(_09128_));
 sky130_fd_sc_hd__o22ai_1 _16055_ (.A1(_08126_),
    .A2(_09127_),
    .B1(_09128_),
    .B2(_08286_),
    .Y(_09129_));
 sky130_fd_sc_hd__nand2_1 _16056_ (.A(_09126_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__or3_1 _16057_ (.A(_08935_),
    .B(_08534_),
    .C(_09130_),
    .X(_09131_));
 sky130_fd_sc_hd__buf_4 _16058_ (.A(_08534_),
    .X(_09132_));
 sky130_fd_sc_hd__o21ai_1 _16059_ (.A1(_08935_),
    .A2(_09132_),
    .B1(_09130_),
    .Y(_09133_));
 sky130_fd_sc_hd__and2_1 _16060_ (.A(_09131_),
    .B(_09133_),
    .X(_09134_));
 sky130_fd_sc_hd__or2_1 _16061_ (.A(_08353_),
    .B(_08325_),
    .X(_09135_));
 sky130_fd_sc_hd__nor2_1 _16062_ (.A(_08351_),
    .B(_08296_),
    .Y(_09136_));
 sky130_fd_sc_hd__xnor2_1 _16063_ (.A(_09135_),
    .B(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__nor2_1 _16064_ (.A(_08211_),
    .B(_08546_),
    .Y(_09138_));
 sky130_fd_sc_hd__xnor2_1 _16065_ (.A(_09137_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__clkbuf_4 _16066_ (.A(_08546_),
    .X(_09140_));
 sky130_fd_sc_hd__nand2_1 _16067_ (.A(_08541_),
    .B(_08998_),
    .Y(_09141_));
 sky130_fd_sc_hd__o31a_1 _16068_ (.A1(_08230_),
    .A2(_09140_),
    .A3(_08999_),
    .B1(_09141_),
    .X(_09142_));
 sky130_fd_sc_hd__nor2_1 _16069_ (.A(_09139_),
    .B(_09142_),
    .Y(_09143_));
 sky130_fd_sc_hd__and2_1 _16070_ (.A(_09139_),
    .B(_09142_),
    .X(_09144_));
 sky130_fd_sc_hd__nor2_1 _16071_ (.A(_09143_),
    .B(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__xnor2_1 _16072_ (.A(_09134_),
    .B(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__a21o_1 _16073_ (.A1(_09124_),
    .A2(_09125_),
    .B1(_09146_),
    .X(_09147_));
 sky130_fd_sc_hd__nand3_1 _16074_ (.A(_09124_),
    .B(_09125_),
    .C(_09146_),
    .Y(_09148_));
 sky130_fd_sc_hd__nand2_1 _16075_ (.A(_09147_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__xnor2_1 _16076_ (.A(_09123_),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__a22o_1 _16077_ (.A1(_08391_),
    .A2(_09014_),
    .B1(_09015_),
    .B2(_09017_),
    .X(_09151_));
 sky130_fd_sc_hd__nand2_1 _16078_ (.A(_08410_),
    .B(_09021_),
    .Y(_09152_));
 sky130_fd_sc_hd__o31a_1 _16079_ (.A1(_08360_),
    .A2(_08411_),
    .A3(_09022_),
    .B1(_09152_),
    .X(_09153_));
 sky130_fd_sc_hd__nor2_1 _16080_ (.A(_08352_),
    .B(_08411_),
    .Y(_09154_));
 sky130_fd_sc_hd__xor2_1 _16081_ (.A(_09014_),
    .B(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__nor2_1 _16082_ (.A(_08394_),
    .B(_08387_),
    .Y(_09156_));
 sky130_fd_sc_hd__xnor2_1 _16083_ (.A(_09155_),
    .B(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__or2_1 _16084_ (.A(_09153_),
    .B(_09157_),
    .X(_09158_));
 sky130_fd_sc_hd__nand2_1 _16085_ (.A(_09153_),
    .B(_09157_),
    .Y(_09159_));
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(_09158_),
    .B(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__xnor2_1 _16087_ (.A(_09151_),
    .B(_09160_),
    .Y(_09161_));
 sky130_fd_sc_hd__nor2_1 _16088_ (.A(_08360_),
    .B(_08409_),
    .Y(_09162_));
 sky130_fd_sc_hd__a21oi_2 _16089_ (.A1(_08454_),
    .A2(_09025_),
    .B1(_08399_),
    .Y(_09163_));
 sky130_fd_sc_hd__a21o_1 _16090_ (.A1(_08454_),
    .A2(_09025_),
    .B1(_08412_),
    .X(_09164_));
 sky130_fd_sc_hd__o21a_1 _16091_ (.A1(_08941_),
    .A2(_08427_),
    .B1(_09164_),
    .X(_09165_));
 sky130_fd_sc_hd__a21oi_2 _16092_ (.A1(_09021_),
    .A2(_09163_),
    .B1(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__xor2_2 _16093_ (.A(_09162_),
    .B(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__nand2_4 _16094_ (.A(\rbzero.wall_tracer.stepDistX[4] ),
    .B(_06162_),
    .Y(_09168_));
 sky130_fd_sc_hd__and2_1 _16095_ (.A(_08448_),
    .B(_09168_),
    .X(_09169_));
 sky130_fd_sc_hd__buf_2 _16096_ (.A(_09169_),
    .X(_09170_));
 sky130_fd_sc_hd__nor2_1 _16097_ (.A(_08928_),
    .B(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__nand2_1 _16098_ (.A(\rbzero.wall_tracer.stepDistY[6] ),
    .B(_08406_),
    .Y(_09172_));
 sky130_fd_sc_hd__o31a_1 _16099_ (.A1(_07989_),
    .A2(_07992_),
    .A3(_08431_),
    .B1(_07994_),
    .X(_09173_));
 sky130_fd_sc_hd__or2_1 _16100_ (.A(_07992_),
    .B(_07994_),
    .X(_09174_));
 sky130_fd_sc_hd__nor3_1 _16101_ (.A(_07989_),
    .B(_08431_),
    .C(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__a21oi_2 _16102_ (.A1(_08120_),
    .A2(_08433_),
    .B1(_08135_),
    .Y(_09176_));
 sky130_fd_sc_hd__o31ai_2 _16103_ (.A1(_08120_),
    .A2(_09173_),
    .A3(_09175_),
    .B1(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__a21oi_1 _16104_ (.A1(_09172_),
    .A2(_09177_),
    .B1(_08830_),
    .Y(_09178_));
 sky130_fd_sc_hd__and3_1 _16105_ (.A(_08618_),
    .B(_09033_),
    .C(_09178_),
    .X(_09179_));
 sky130_fd_sc_hd__a21o_2 _16106_ (.A1(_09031_),
    .A2(_09032_),
    .B1(_06162_),
    .X(_09180_));
 sky130_fd_sc_hd__a21o_2 _16107_ (.A1(_09172_),
    .A2(_09177_),
    .B1(_06162_),
    .X(_09181_));
 sky130_fd_sc_hd__o22ai_1 _16108_ (.A1(_08447_),
    .A2(_09180_),
    .B1(_09181_),
    .B2(_08450_),
    .Y(_09182_));
 sky130_fd_sc_hd__or2b_1 _16109_ (.A(_09179_),
    .B_N(_09182_),
    .X(_09183_));
 sky130_fd_sc_hd__xnor2_2 _16110_ (.A(_09171_),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__nor2_1 _16111_ (.A(_09028_),
    .B(_09034_),
    .Y(_09185_));
 sky130_fd_sc_hd__a21oi_2 _16112_ (.A1(_09027_),
    .A2(_09035_),
    .B1(_09185_),
    .Y(_09186_));
 sky130_fd_sc_hd__xnor2_2 _16113_ (.A(_09184_),
    .B(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__xnor2_2 _16114_ (.A(_09167_),
    .B(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__nor2_1 _16115_ (.A(_09036_),
    .B(_09038_),
    .Y(_09189_));
 sky130_fd_sc_hd__a21o_1 _16116_ (.A1(_09024_),
    .A2(_09039_),
    .B1(_09189_),
    .X(_09190_));
 sky130_fd_sc_hd__xnor2_1 _16117_ (.A(_09188_),
    .B(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__xnor2_1 _16118_ (.A(_09161_),
    .B(_09191_),
    .Y(_09192_));
 sky130_fd_sc_hd__and2b_1 _16119_ (.A_N(_09040_),
    .B(_09042_),
    .X(_09193_));
 sky130_fd_sc_hd__a21oi_1 _16120_ (.A1(_09020_),
    .A2(_09043_),
    .B1(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__nor2_1 _16121_ (.A(_09192_),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__and2_1 _16122_ (.A(_09192_),
    .B(_09194_),
    .X(_09196_));
 sky130_fd_sc_hd__nor2_1 _16123_ (.A(_09195_),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__xnor2_1 _16124_ (.A(_09150_),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__nor2_1 _16125_ (.A(_09044_),
    .B(_09046_),
    .Y(_09199_));
 sky130_fd_sc_hd__a21oi_1 _16126_ (.A1(_09011_),
    .A2(_09047_),
    .B1(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__xor2_1 _16127_ (.A(_09198_),
    .B(_09200_),
    .X(_09201_));
 sky130_fd_sc_hd__xnor2_1 _16128_ (.A(_09122_),
    .B(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__a21oi_1 _16129_ (.A1(_09052_),
    .A2(_09069_),
    .B1(_09051_),
    .Y(_09203_));
 sky130_fd_sc_hd__nor2_1 _16130_ (.A(_09202_),
    .B(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__nand2_1 _16131_ (.A(_09202_),
    .B(_09203_),
    .Y(_09205_));
 sky130_fd_sc_hd__and2b_1 _16132_ (.A_N(_09204_),
    .B(_09205_),
    .X(_09206_));
 sky130_fd_sc_hd__xnor2_2 _16133_ (.A(_09067_),
    .B(_09206_),
    .Y(_09207_));
 sky130_fd_sc_hd__nor2_1 _16134_ (.A(_09070_),
    .B(_09072_),
    .Y(_09208_));
 sky130_fd_sc_hd__a21oi_2 _16135_ (.A1(_08607_),
    .A2(_09073_),
    .B1(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__xnor2_4 _16136_ (.A(_09207_),
    .B(_09209_),
    .Y(_09210_));
 sky130_fd_sc_hd__xor2_4 _16137_ (.A(_09106_),
    .B(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__xnor2_4 _16138_ (.A(_09105_),
    .B(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__and2b_1 _16139_ (.A_N(_04511_),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .X(_09213_));
 sky130_fd_sc_hd__a21oi_1 _16140_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_08115_),
    .B1(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__nor2_1 _16141_ (.A(_09212_),
    .B(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__and2_1 _16142_ (.A(_09212_),
    .B(_09214_),
    .X(_09216_));
 sky130_fd_sc_hd__or2_1 _16143_ (.A(_09215_),
    .B(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__a21oi_1 _16144_ (.A1(_09085_),
    .A2(_09097_),
    .B1(_09083_),
    .Y(_09218_));
 sky130_fd_sc_hd__xnor2_1 _16145_ (.A(_09217_),
    .B(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__nor2_1 _16146_ (.A(_09102_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__a211o_1 _16147_ (.A1(_09102_),
    .A2(_09219_),
    .B1(_09220_),
    .C1(_08429_),
    .X(_09221_));
 sky130_fd_sc_hd__o211a_1 _16148_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_08120_),
    .B1(_09221_),
    .C1(_08059_),
    .X(_00467_));
 sky130_fd_sc_hd__or2_2 _16149_ (.A(_09207_),
    .B(_09209_),
    .X(_09222_));
 sky130_fd_sc_hd__a31o_1 _16150_ (.A1(_08604_),
    .A2(_09063_),
    .A3(_09121_),
    .B1(_09119_),
    .X(_09223_));
 sky130_fd_sc_hd__or2b_1 _16151_ (.A(_09149_),
    .B_N(_09123_),
    .X(_09224_));
 sky130_fd_sc_hd__nand2_1 _16152_ (.A(_09147_),
    .B(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__nand2_2 _16153_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08523_),
    .Y(_09226_));
 sky130_fd_sc_hd__clkbuf_4 _16154_ (.A(_09226_),
    .X(_09227_));
 sky130_fd_sc_hd__buf_4 _16155_ (.A(_09227_),
    .X(_09228_));
 sky130_fd_sc_hd__nor2_1 _16156_ (.A(_08598_),
    .B(_09228_),
    .Y(_09229_));
 sky130_fd_sc_hd__or2_1 _16157_ (.A(_08520_),
    .B(_09055_),
    .X(_09230_));
 sky130_fd_sc_hd__or3_1 _16158_ (.A(_08285_),
    .B(_08600_),
    .C(_09230_),
    .X(_09231_));
 sky130_fd_sc_hd__a21bo_1 _16159_ (.A1(_09109_),
    .A2(_09112_),
    .B1_N(_09231_),
    .X(_09232_));
 sky130_fd_sc_hd__or2_1 _16160_ (.A(_08278_),
    .B(_08599_),
    .X(_09233_));
 sky130_fd_sc_hd__xnor2_1 _16161_ (.A(_09230_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__or3_1 _16162_ (.A(_08147_),
    .B(_09110_),
    .C(_09234_),
    .X(_09235_));
 sky130_fd_sc_hd__o21ai_1 _16163_ (.A1(_08285_),
    .A2(_09111_),
    .B1(_09234_),
    .Y(_09236_));
 sky130_fd_sc_hd__nand2_1 _16164_ (.A(_09235_),
    .B(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__a21o_1 _16165_ (.A1(_09126_),
    .A2(_09131_),
    .B1(_09237_),
    .X(_09238_));
 sky130_fd_sc_hd__nand3_1 _16166_ (.A(_09126_),
    .B(_09131_),
    .C(_09237_),
    .Y(_09239_));
 sky130_fd_sc_hd__nand2_1 _16167_ (.A(_09238_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__xnor2_1 _16168_ (.A(_09232_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__o21ba_1 _16169_ (.A1(_09058_),
    .A2(_09115_),
    .B1_N(_09114_),
    .X(_09242_));
 sky130_fd_sc_hd__xor2_1 _16170_ (.A(_09241_),
    .B(_09242_),
    .X(_09243_));
 sky130_fd_sc_hd__and2_1 _16171_ (.A(_09229_),
    .B(_09243_),
    .X(_09244_));
 sky130_fd_sc_hd__nor2_1 _16172_ (.A(_09229_),
    .B(_09243_),
    .Y(_09245_));
 sky130_fd_sc_hd__or2_1 _16173_ (.A(_09244_),
    .B(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__xor2_2 _16174_ (.A(_09225_),
    .B(_09246_),
    .X(_09247_));
 sky130_fd_sc_hd__or3b_2 _16175_ (.A(_09114_),
    .B(_09115_),
    .C_N(_09061_),
    .X(_09248_));
 sky130_fd_sc_hd__xor2_2 _16176_ (.A(_09247_),
    .B(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__a21o_1 _16177_ (.A1(_09134_),
    .A2(_09145_),
    .B1(_09143_),
    .X(_09250_));
 sky130_fd_sc_hd__or2b_1 _16178_ (.A(_09160_),
    .B_N(_09151_),
    .X(_09251_));
 sky130_fd_sc_hd__clkbuf_2 _16179_ (.A(_08209_),
    .X(_09252_));
 sky130_fd_sc_hd__or4_1 _16180_ (.A(_08126_),
    .B(_08286_),
    .C(_09252_),
    .D(_08245_),
    .X(_09253_));
 sky130_fd_sc_hd__o22ai_1 _16181_ (.A1(_08127_),
    .A2(_09252_),
    .B1(_09127_),
    .B2(_08286_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand2_1 _16182_ (.A(_09253_),
    .B(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__nor2_1 _16183_ (.A(_09128_),
    .B(_08534_),
    .Y(_09256_));
 sky130_fd_sc_hd__xnor2_1 _16184_ (.A(_09255_),
    .B(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_08325_),
    .B(_08387_),
    .Y(_09258_));
 sky130_fd_sc_hd__o22a_1 _16186_ (.A1(_08351_),
    .A2(_08325_),
    .B1(_08387_),
    .B2(_08797_),
    .X(_09259_));
 sky130_fd_sc_hd__a21o_1 _16187_ (.A1(_09136_),
    .A2(_09258_),
    .B1(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__or2_1 _16188_ (.A(_08353_),
    .B(_08546_),
    .X(_09261_));
 sky130_fd_sc_hd__xnor2_1 _16189_ (.A(_09260_),
    .B(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__and2b_1 _16190_ (.A_N(_09135_),
    .B(_09136_),
    .X(_09263_));
 sky130_fd_sc_hd__a21oi_1 _16191_ (.A1(_09137_),
    .A2(_09138_),
    .B1(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__nor2_1 _16192_ (.A(_09262_),
    .B(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__and2_1 _16193_ (.A(_09262_),
    .B(_09264_),
    .X(_09266_));
 sky130_fd_sc_hd__nor2_1 _16194_ (.A(_09265_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__xnor2_1 _16195_ (.A(_09257_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__a21o_1 _16196_ (.A1(_09158_),
    .A2(_09251_),
    .B1(_09268_),
    .X(_09269_));
 sky130_fd_sc_hd__nand3_1 _16197_ (.A(_09158_),
    .B(_09251_),
    .C(_09268_),
    .Y(_09270_));
 sky130_fd_sc_hd__nand2_1 _16198_ (.A(_09269_),
    .B(_09270_),
    .Y(_09271_));
 sky130_fd_sc_hd__xnor2_1 _16199_ (.A(_09250_),
    .B(_09271_),
    .Y(_09272_));
 sky130_fd_sc_hd__a22o_1 _16200_ (.A1(_09014_),
    .A2(_09154_),
    .B1(_09155_),
    .B2(_09156_),
    .X(_09273_));
 sky130_fd_sc_hd__a22o_1 _16201_ (.A1(_09021_),
    .A2(_09163_),
    .B1(_09166_),
    .B2(_09162_),
    .X(_09274_));
 sky130_fd_sc_hd__o22a_1 _16202_ (.A1(_08876_),
    .A2(_08411_),
    .B1(_08409_),
    .B2(_08352_),
    .X(_09275_));
 sky130_fd_sc_hd__a31o_1 _16203_ (.A1(_08247_),
    .A2(_08456_),
    .A3(_09154_),
    .B1(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__nor3_1 _16204_ (.A(_08394_),
    .B(_08378_),
    .C(_09276_),
    .Y(_09277_));
 sky130_fd_sc_hd__o21a_1 _16205_ (.A1(_08394_),
    .A2(_08378_),
    .B1(_09276_),
    .X(_09278_));
 sky130_fd_sc_hd__nor2_1 _16206_ (.A(_09277_),
    .B(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__xor2_1 _16207_ (.A(_09274_),
    .B(_09279_),
    .X(_09280_));
 sky130_fd_sc_hd__xor2_1 _16208_ (.A(_09273_),
    .B(_09280_),
    .X(_09281_));
 sky130_fd_sc_hd__nor2_1 _16209_ (.A(_08359_),
    .B(_08427_),
    .Y(_09282_));
 sky130_fd_sc_hd__a21oi_1 _16210_ (.A1(_08448_),
    .A2(_09168_),
    .B1(_08412_),
    .Y(_09283_));
 sky130_fd_sc_hd__xor2_1 _16211_ (.A(_09163_),
    .B(_09283_),
    .X(_09284_));
 sky130_fd_sc_hd__xor2_1 _16212_ (.A(_09282_),
    .B(_09284_),
    .X(_09285_));
 sky130_fd_sc_hd__clkbuf_4 _16213_ (.A(_09180_),
    .X(_09286_));
 sky130_fd_sc_hd__nand2_2 _16214_ (.A(\rbzero.wall_tracer.stepDistX[5] ),
    .B(_06163_),
    .Y(_09287_));
 sky130_fd_sc_hd__a21oi_1 _16215_ (.A1(_09286_),
    .A2(_09287_),
    .B1(_08420_),
    .Y(_09288_));
 sky130_fd_sc_hd__nor4_1 _16216_ (.A(_07989_),
    .B(_07999_),
    .C(_08431_),
    .D(_09174_),
    .Y(_09289_));
 sky130_fd_sc_hd__o31a_1 _16217_ (.A1(_07989_),
    .A2(_08431_),
    .A3(_09174_),
    .B1(_07999_),
    .X(_09290_));
 sky130_fd_sc_hd__o31a_2 _16218_ (.A1(_08120_),
    .A2(_09289_),
    .A3(_09290_),
    .B1(_09176_),
    .X(_09291_));
 sky130_fd_sc_hd__and3_1 _16219_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08124_),
    .C(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__xor2_1 _16220_ (.A(_09178_),
    .B(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__xor2_1 _16221_ (.A(_09288_),
    .B(_09293_),
    .X(_09294_));
 sky130_fd_sc_hd__clkbuf_4 _16222_ (.A(_08448_),
    .X(_09295_));
 sky130_fd_sc_hd__nand2_1 _16223_ (.A(_09295_),
    .B(_09168_),
    .Y(_09296_));
 sky130_fd_sc_hd__a31o_1 _16224_ (.A1(_08457_),
    .A2(_09296_),
    .A3(_09182_),
    .B1(_09179_),
    .X(_09297_));
 sky130_fd_sc_hd__xor2_1 _16225_ (.A(_09294_),
    .B(_09297_),
    .X(_09298_));
 sky130_fd_sc_hd__xnor2_1 _16226_ (.A(_09285_),
    .B(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__or2b_1 _16227_ (.A(_09186_),
    .B_N(_09184_),
    .X(_09300_));
 sky130_fd_sc_hd__a21boi_1 _16228_ (.A1(_09167_),
    .A2(_09187_),
    .B1_N(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__xor2_1 _16229_ (.A(_09299_),
    .B(_09301_),
    .X(_09302_));
 sky130_fd_sc_hd__xnor2_1 _16230_ (.A(_09281_),
    .B(_09302_),
    .Y(_09303_));
 sky130_fd_sc_hd__and2b_1 _16231_ (.A_N(_09188_),
    .B(_09190_),
    .X(_09304_));
 sky130_fd_sc_hd__a21oi_1 _16232_ (.A1(_09161_),
    .A2(_09191_),
    .B1(_09304_),
    .Y(_09305_));
 sky130_fd_sc_hd__nor2_1 _16233_ (.A(_09303_),
    .B(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand2_1 _16234_ (.A(_09303_),
    .B(_09305_),
    .Y(_09307_));
 sky130_fd_sc_hd__and2b_1 _16235_ (.A_N(_09306_),
    .B(_09307_),
    .X(_09308_));
 sky130_fd_sc_hd__xnor2_1 _16236_ (.A(_09272_),
    .B(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__a21oi_1 _16237_ (.A1(_09150_),
    .A2(_09197_),
    .B1(_09195_),
    .Y(_09310_));
 sky130_fd_sc_hd__nor2_1 _16238_ (.A(_09309_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__and2_1 _16239_ (.A(_09309_),
    .B(_09310_),
    .X(_09312_));
 sky130_fd_sc_hd__nor2_1 _16240_ (.A(_09311_),
    .B(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__xnor2_2 _16241_ (.A(_09249_),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(_09198_),
    .B(_09200_),
    .Y(_09315_));
 sky130_fd_sc_hd__a21oi_2 _16243_ (.A1(_09122_),
    .A2(_09201_),
    .B1(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__xor2_2 _16244_ (.A(_09314_),
    .B(_09316_),
    .X(_09317_));
 sky130_fd_sc_hd__xnor2_2 _16245_ (.A(_09223_),
    .B(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__a21oi_1 _16246_ (.A1(_09067_),
    .A2(_09205_),
    .B1(_09204_),
    .Y(_09319_));
 sky130_fd_sc_hd__xor2_2 _16247_ (.A(_09318_),
    .B(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__xnor2_4 _16248_ (.A(_09222_),
    .B(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__a21oi_1 _16249_ (.A1(_09106_),
    .A2(_09079_),
    .B1(_09210_),
    .Y(_09322_));
 sky130_fd_sc_hd__a31o_2 _16250_ (.A1(_08988_),
    .A2(_09081_),
    .A3(_09211_),
    .B1(_09322_),
    .X(_09323_));
 sky130_fd_sc_hd__xnor2_4 _16251_ (.A(_09321_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__and2b_1 _16252_ (.A_N(_08115_),
    .B(\rbzero.debug_overlay.playerY[-4] ),
    .X(_09325_));
 sky130_fd_sc_hd__a21oi_1 _16253_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_08115_),
    .B1(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__nor2_1 _16254_ (.A(_09324_),
    .B(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__and2_1 _16255_ (.A(_09324_),
    .B(_09326_),
    .X(_09328_));
 sky130_fd_sc_hd__or2_1 _16256_ (.A(_09327_),
    .B(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__o21ba_1 _16257_ (.A1(_09217_),
    .A2(_09218_),
    .B1_N(_09215_),
    .X(_09330_));
 sky130_fd_sc_hd__xnor2_1 _16258_ (.A(_09329_),
    .B(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__xnor2_1 _16259_ (.A(_09102_),
    .B(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__or2_1 _16260_ (.A(\rbzero.texu_hot[2] ),
    .B(_08120_),
    .X(_09333_));
 sky130_fd_sc_hd__o211a_1 _16261_ (.A1(_08429_),
    .A2(_09332_),
    .B1(_09333_),
    .C1(_08059_),
    .X(_00468_));
 sky130_fd_sc_hd__or2b_1 _16262_ (.A(_09222_),
    .B_N(_09320_),
    .X(_09334_));
 sky130_fd_sc_hd__a21boi_2 _16263_ (.A1(_09321_),
    .A2(_09323_),
    .B1_N(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__or2_1 _16264_ (.A(_09318_),
    .B(_09319_),
    .X(_09336_));
 sky130_fd_sc_hd__a21o_1 _16265_ (.A1(_09147_),
    .A2(_09224_),
    .B1(_09246_),
    .X(_09337_));
 sky130_fd_sc_hd__o21ai_1 _16266_ (.A1(_09247_),
    .A2(_09248_),
    .B1(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__a21o_1 _16267_ (.A1(_09241_),
    .A2(_09242_),
    .B1(_09244_),
    .X(_09339_));
 sky130_fd_sc_hd__or2b_1 _16268_ (.A(_09271_),
    .B_N(_09250_),
    .X(_09340_));
 sky130_fd_sc_hd__nand2_4 _16269_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08523_),
    .Y(_09341_));
 sky130_fd_sc_hd__buf_4 _16270_ (.A(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__nor2_1 _16271_ (.A(_08285_),
    .B(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__o22a_1 _16272_ (.A1(_08285_),
    .A2(_09228_),
    .B1(_09342_),
    .B2(_08598_),
    .X(_09344_));
 sky130_fd_sc_hd__a21oi_1 _16273_ (.A1(_09229_),
    .A2(_09343_),
    .B1(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__o21ai_1 _16274_ (.A1(_09230_),
    .A2(_09233_),
    .B1(_09235_),
    .Y(_09346_));
 sky130_fd_sc_hd__a21bo_1 _16275_ (.A1(_09254_),
    .A2(_09256_),
    .B1_N(_09253_),
    .X(_09347_));
 sky130_fd_sc_hd__nor2_1 _16276_ (.A(_08278_),
    .B(_09055_),
    .Y(_09348_));
 sky130_fd_sc_hd__nor2_1 _16277_ (.A(_08860_),
    .B(_08599_),
    .Y(_09349_));
 sky130_fd_sc_hd__xnor2_1 _16278_ (.A(_09348_),
    .B(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__or3_1 _16279_ (.A(_08520_),
    .B(_09110_),
    .C(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__o21ai_1 _16280_ (.A1(_08602_),
    .A2(_09110_),
    .B1(_09350_),
    .Y(_09352_));
 sky130_fd_sc_hd__and2_1 _16281_ (.A(_09351_),
    .B(_09352_),
    .X(_09353_));
 sky130_fd_sc_hd__and2_1 _16282_ (.A(_09347_),
    .B(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__or2_1 _16283_ (.A(_09347_),
    .B(_09353_),
    .X(_09355_));
 sky130_fd_sc_hd__and2b_1 _16284_ (.A_N(_09354_),
    .B(_09355_),
    .X(_09356_));
 sky130_fd_sc_hd__xnor2_1 _16285_ (.A(_09346_),
    .B(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__inv_2 _16286_ (.A(_09232_),
    .Y(_09358_));
 sky130_fd_sc_hd__o21a_1 _16287_ (.A1(_09358_),
    .A2(_09240_),
    .B1(_09238_),
    .X(_09359_));
 sky130_fd_sc_hd__xor2_1 _16288_ (.A(_09357_),
    .B(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__xnor2_1 _16289_ (.A(_09345_),
    .B(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__a21o_1 _16290_ (.A1(_09269_),
    .A2(_09340_),
    .B1(_09361_),
    .X(_09362_));
 sky130_fd_sc_hd__nand3_1 _16291_ (.A(_09269_),
    .B(_09340_),
    .C(_09361_),
    .Y(_09363_));
 sky130_fd_sc_hd__nand2_1 _16292_ (.A(_09362_),
    .B(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__xnor2_1 _16293_ (.A(_09339_),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__a21o_1 _16294_ (.A1(_09257_),
    .A2(_09267_),
    .B1(_09265_),
    .X(_09366_));
 sky130_fd_sc_hd__nand2_1 _16295_ (.A(_09274_),
    .B(_09279_),
    .Y(_09367_));
 sky130_fd_sc_hd__a21bo_1 _16296_ (.A1(_09273_),
    .A2(_09280_),
    .B1_N(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__buf_2 _16297_ (.A(_08176_),
    .X(_09369_));
 sky130_fd_sc_hd__o22ai_1 _16298_ (.A1(_08127_),
    .A2(_09369_),
    .B1(_09252_),
    .B2(_08286_),
    .Y(_09370_));
 sky130_fd_sc_hd__or4_1 _16299_ (.A(_08126_),
    .B(_08286_),
    .C(_09369_),
    .D(_09252_),
    .X(_09371_));
 sky130_fd_sc_hd__nand2_1 _16300_ (.A(_09370_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__nor2_1 _16301_ (.A(_09127_),
    .B(_08534_),
    .Y(_09373_));
 sky130_fd_sc_hd__xnor2_2 _16302_ (.A(_09372_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__nor2_1 _16303_ (.A(_08797_),
    .B(_08378_),
    .Y(_09375_));
 sky130_fd_sc_hd__xnor2_1 _16304_ (.A(_09258_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__or2_1 _16305_ (.A(_08351_),
    .B(_08546_),
    .X(_09377_));
 sky130_fd_sc_hd__xnor2_1 _16306_ (.A(_09376_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__nand2_1 _16307_ (.A(_09136_),
    .B(_09258_),
    .Y(_09379_));
 sky130_fd_sc_hd__o31a_1 _16308_ (.A1(_08353_),
    .A2(_09140_),
    .A3(_09259_),
    .B1(_09379_),
    .X(_09380_));
 sky130_fd_sc_hd__nor2_1 _16309_ (.A(_09378_),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__and2_1 _16310_ (.A(_09378_),
    .B(_09380_),
    .X(_09382_));
 sky130_fd_sc_hd__nor2_1 _16311_ (.A(_09381_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__xor2_2 _16312_ (.A(_09374_),
    .B(_09383_),
    .X(_09384_));
 sky130_fd_sc_hd__xnor2_1 _16313_ (.A(_09368_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__xnor2_1 _16314_ (.A(_09366_),
    .B(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__a31o_1 _16315_ (.A1(_08247_),
    .A2(_08456_),
    .A3(_09154_),
    .B1(_09277_),
    .X(_09387_));
 sky130_fd_sc_hd__a22o_1 _16316_ (.A1(_09163_),
    .A2(_09283_),
    .B1(_09284_),
    .B2(_09282_),
    .X(_09388_));
 sky130_fd_sc_hd__or4_1 _16317_ (.A(_08352_),
    .B(_08243_),
    .C(_08408_),
    .D(_08426_),
    .X(_09389_));
 sky130_fd_sc_hd__a2bb2o_1 _16318_ (.A1_N(_08352_),
    .A2_N(_08427_),
    .B1(_08247_),
    .B2(_08456_),
    .X(_09390_));
 sky130_fd_sc_hd__nor2_1 _16319_ (.A(_08267_),
    .B(_08411_),
    .Y(_09391_));
 sky130_fd_sc_hd__and3_1 _16320_ (.A(_09389_),
    .B(_09390_),
    .C(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__a21oi_1 _16321_ (.A1(_09389_),
    .A2(_09390_),
    .B1(_09391_),
    .Y(_09393_));
 sky130_fd_sc_hd__nor2_1 _16322_ (.A(_09392_),
    .B(_09393_),
    .Y(_09394_));
 sky130_fd_sc_hd__xnor2_1 _16323_ (.A(_09388_),
    .B(_09394_),
    .Y(_09395_));
 sky130_fd_sc_hd__xnor2_1 _16324_ (.A(_09387_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__a21oi_1 _16325_ (.A1(_08454_),
    .A2(_09025_),
    .B1(_08359_),
    .Y(_09397_));
 sky130_fd_sc_hd__a21o_1 _16326_ (.A1(_08448_),
    .A2(_09168_),
    .B1(_08399_),
    .X(_09398_));
 sky130_fd_sc_hd__a21oi_1 _16327_ (.A1(_09180_),
    .A2(_09287_),
    .B1(_08412_),
    .Y(_09399_));
 sky130_fd_sc_hd__xnor2_1 _16328_ (.A(_09398_),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__xor2_1 _16329_ (.A(_09397_),
    .B(_09400_),
    .X(_09401_));
 sky130_fd_sc_hd__nand2_1 _16330_ (.A(\rbzero.wall_tracer.stepDistX[6] ),
    .B(_06163_),
    .Y(_09402_));
 sky130_fd_sc_hd__and2_1 _16331_ (.A(_09181_),
    .B(_09402_),
    .X(_09403_));
 sky130_fd_sc_hd__o41a_1 _16332_ (.A1(_07988_),
    .A2(_07999_),
    .A3(_08431_),
    .A4(_09174_),
    .B1(_08003_),
    .X(_09404_));
 sky130_fd_sc_hd__a211o_1 _16333_ (.A1(_08002_),
    .A2(_09289_),
    .B1(_09404_),
    .C1(_08120_),
    .X(_09405_));
 sky130_fd_sc_hd__a22oi_4 _16334_ (.A1(\rbzero.wall_tracer.stepDistY[8] ),
    .A2(_08406_),
    .B1(_09176_),
    .B2(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__and3_1 _16335_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_08124_),
    .C(_09291_),
    .X(_09407_));
 sky130_fd_sc_hd__or4b_1 _16336_ (.A(_06163_),
    .B(_08450_),
    .C(_09406_),
    .D_N(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__a21oi_4 _16337_ (.A1(\rbzero.wall_tracer.stepDistY[7] ),
    .A2(_08406_),
    .B1(_09291_),
    .Y(_09409_));
 sky130_fd_sc_hd__o32ai_1 _16338_ (.A1(_06163_),
    .A2(_08450_),
    .A3(_09406_),
    .B1(_09409_),
    .B2(_08830_),
    .Y(_09410_));
 sky130_fd_sc_hd__or4bb_1 _16339_ (.A(_08928_),
    .B(_09403_),
    .C_N(_09408_),
    .D_N(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__a2bb2o_1 _16340_ (.A1_N(_08928_),
    .A2_N(_09403_),
    .B1(_09408_),
    .B2(_09410_),
    .X(_09412_));
 sky130_fd_sc_hd__nand2_1 _16341_ (.A(_09178_),
    .B(_09292_),
    .Y(_09413_));
 sky130_fd_sc_hd__a21bo_1 _16342_ (.A1(_09288_),
    .A2(_09293_),
    .B1_N(_09413_),
    .X(_09414_));
 sky130_fd_sc_hd__nand3_1 _16343_ (.A(_09411_),
    .B(_09412_),
    .C(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__a21o_1 _16344_ (.A1(_09411_),
    .A2(_09412_),
    .B1(_09414_),
    .X(_09416_));
 sky130_fd_sc_hd__nand3_1 _16345_ (.A(_09401_),
    .B(_09415_),
    .C(_09416_),
    .Y(_09417_));
 sky130_fd_sc_hd__a21o_1 _16346_ (.A1(_09415_),
    .A2(_09416_),
    .B1(_09401_),
    .X(_09418_));
 sky130_fd_sc_hd__and2_1 _16347_ (.A(_09294_),
    .B(_09297_),
    .X(_09419_));
 sky130_fd_sc_hd__a21o_1 _16348_ (.A1(_09285_),
    .A2(_09298_),
    .B1(_09419_),
    .X(_09420_));
 sky130_fd_sc_hd__nand3_1 _16349_ (.A(_09417_),
    .B(_09418_),
    .C(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__a21o_1 _16350_ (.A1(_09417_),
    .A2(_09418_),
    .B1(_09420_),
    .X(_09422_));
 sky130_fd_sc_hd__and3_1 _16351_ (.A(_09396_),
    .B(_09421_),
    .C(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__a21oi_1 _16352_ (.A1(_09421_),
    .A2(_09422_),
    .B1(_09396_),
    .Y(_09424_));
 sky130_fd_sc_hd__or2_1 _16353_ (.A(_09423_),
    .B(_09424_),
    .X(_09425_));
 sky130_fd_sc_hd__nor2_1 _16354_ (.A(_09299_),
    .B(_09301_),
    .Y(_09426_));
 sky130_fd_sc_hd__a21oi_1 _16355_ (.A1(_09281_),
    .A2(_09302_),
    .B1(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__xor2_1 _16356_ (.A(_09425_),
    .B(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__nand2_1 _16357_ (.A(_09386_),
    .B(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__or2_1 _16358_ (.A(_09386_),
    .B(_09428_),
    .X(_09430_));
 sky130_fd_sc_hd__nand2_1 _16359_ (.A(_09429_),
    .B(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__a21oi_1 _16360_ (.A1(_09272_),
    .A2(_09307_),
    .B1(_09306_),
    .Y(_09432_));
 sky130_fd_sc_hd__nor2_1 _16361_ (.A(_09431_),
    .B(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__and2_1 _16362_ (.A(_09431_),
    .B(_09432_),
    .X(_09434_));
 sky130_fd_sc_hd__nor2_1 _16363_ (.A(_09433_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__xnor2_1 _16364_ (.A(_09365_),
    .B(_09435_),
    .Y(_09436_));
 sky130_fd_sc_hd__a21oi_1 _16365_ (.A1(_09249_),
    .A2(_09313_),
    .B1(_09311_),
    .Y(_09437_));
 sky130_fd_sc_hd__xnor2_1 _16366_ (.A(_09436_),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__xor2_1 _16367_ (.A(_09338_),
    .B(_09438_),
    .X(_09439_));
 sky130_fd_sc_hd__nor2_1 _16368_ (.A(_09314_),
    .B(_09316_),
    .Y(_09440_));
 sky130_fd_sc_hd__a21oi_1 _16369_ (.A1(_09223_),
    .A2(_09317_),
    .B1(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__nor2_2 _16370_ (.A(_09439_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__and2_1 _16371_ (.A(_09439_),
    .B(_09441_),
    .X(_09443_));
 sky130_fd_sc_hd__or2_1 _16372_ (.A(_09442_),
    .B(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__xor2_2 _16373_ (.A(_09336_),
    .B(_09444_),
    .X(_09445_));
 sky130_fd_sc_hd__xor2_4 _16374_ (.A(_09335_),
    .B(_09445_),
    .X(_09446_));
 sky130_fd_sc_hd__mux2_1 _16375_ (.A0(_05056_),
    .A1(_05059_),
    .S(_08115_),
    .X(_09447_));
 sky130_fd_sc_hd__nor2_1 _16376_ (.A(_09446_),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__and2_1 _16377_ (.A(_09446_),
    .B(_09447_),
    .X(_09449_));
 sky130_fd_sc_hd__or2_1 _16378_ (.A(_09448_),
    .B(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__o21ba_1 _16379_ (.A1(_09329_),
    .A2(_09330_),
    .B1_N(_09327_),
    .X(_09451_));
 sky130_fd_sc_hd__xnor2_1 _16380_ (.A(_09450_),
    .B(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__nor2_1 _16381_ (.A(_09102_),
    .B(_09452_),
    .Y(_09453_));
 sky130_fd_sc_hd__a211o_1 _16382_ (.A1(_09102_),
    .A2(_09452_),
    .B1(_09453_),
    .C1(_08429_),
    .X(_09454_));
 sky130_fd_sc_hd__o211a_1 _16383_ (.A1(\rbzero.texu_hot[3] ),
    .A2(_08120_),
    .B1(_09454_),
    .C1(_08059_),
    .X(_00469_));
 sky130_fd_sc_hd__o21ba_1 _16384_ (.A1(_09450_),
    .A2(_09451_),
    .B1_N(_09448_),
    .X(_09455_));
 sky130_fd_sc_hd__a21oi_1 _16385_ (.A1(_09336_),
    .A2(_09334_),
    .B1(_09444_),
    .Y(_09456_));
 sky130_fd_sc_hd__a31o_2 _16386_ (.A1(_09321_),
    .A2(_09323_),
    .A3(_09445_),
    .B1(_09456_),
    .X(_09457_));
 sky130_fd_sc_hd__or2b_1 _16387_ (.A(_09438_),
    .B_N(_09338_),
    .X(_09458_));
 sky130_fd_sc_hd__o21ai_2 _16388_ (.A1(_09436_),
    .A2(_09437_),
    .B1(_09458_),
    .Y(_09459_));
 sky130_fd_sc_hd__or2b_1 _16389_ (.A(_09364_),
    .B_N(_09339_),
    .X(_09460_));
 sky130_fd_sc_hd__nand2_1 _16390_ (.A(_09362_),
    .B(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__a2bb2o_1 _16391_ (.A1_N(_09357_),
    .A2_N(_09359_),
    .B1(_09360_),
    .B2(_09345_),
    .X(_09462_));
 sky130_fd_sc_hd__nand2_1 _16392_ (.A(_09368_),
    .B(_09384_),
    .Y(_09463_));
 sky130_fd_sc_hd__or2b_1 _16393_ (.A(_09385_),
    .B_N(_09366_),
    .X(_09464_));
 sky130_fd_sc_hd__nand2_1 _16394_ (.A(_09229_),
    .B(_09343_),
    .Y(_09465_));
 sky130_fd_sc_hd__nor2_1 _16395_ (.A(_08602_),
    .B(_09227_),
    .Y(_09466_));
 sky130_fd_sc_hd__xnor2_1 _16396_ (.A(_09343_),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__nand2_1 _16397_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_08523_),
    .Y(_09468_));
 sky130_fd_sc_hd__clkbuf_4 _16398_ (.A(_09468_),
    .X(_09469_));
 sky130_fd_sc_hd__nor2_1 _16399_ (.A(_08598_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__xnor2_1 _16400_ (.A(_09467_),
    .B(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__xnor2_1 _16401_ (.A(_09465_),
    .B(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__a21bo_1 _16402_ (.A1(_09348_),
    .A2(_09349_),
    .B1_N(_09351_),
    .X(_09473_));
 sky130_fd_sc_hd__or2_1 _16403_ (.A(_08935_),
    .B(_09110_),
    .X(_09474_));
 sky130_fd_sc_hd__o22a_1 _16404_ (.A1(_08245_),
    .A2(_08599_),
    .B1(_09055_),
    .B2(_08860_),
    .X(_09475_));
 sky130_fd_sc_hd__or2_1 _16405_ (.A(_08245_),
    .B(_09055_),
    .X(_09476_));
 sky130_fd_sc_hd__or3_1 _16406_ (.A(_08860_),
    .B(_08599_),
    .C(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__and2b_1 _16407_ (.A_N(_09475_),
    .B(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__xor2_1 _16408_ (.A(_09474_),
    .B(_09478_),
    .X(_09479_));
 sky130_fd_sc_hd__a21bo_1 _16409_ (.A1(_09370_),
    .A2(_09373_),
    .B1_N(_09371_),
    .X(_09480_));
 sky130_fd_sc_hd__and2b_1 _16410_ (.A_N(_09479_),
    .B(_09480_),
    .X(_09481_));
 sky130_fd_sc_hd__and2b_1 _16411_ (.A_N(_09480_),
    .B(_09479_),
    .X(_09482_));
 sky130_fd_sc_hd__nor2_1 _16412_ (.A(_09481_),
    .B(_09482_),
    .Y(_09483_));
 sky130_fd_sc_hd__xnor2_1 _16413_ (.A(_09473_),
    .B(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__a21oi_1 _16414_ (.A1(_09346_),
    .A2(_09356_),
    .B1(_09354_),
    .Y(_09485_));
 sky130_fd_sc_hd__nor2_1 _16415_ (.A(_09484_),
    .B(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__and2_1 _16416_ (.A(_09484_),
    .B(_09485_),
    .X(_09487_));
 sky130_fd_sc_hd__nor2_1 _16417_ (.A(_09486_),
    .B(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__xnor2_1 _16418_ (.A(_09472_),
    .B(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__a21o_1 _16419_ (.A1(_09463_),
    .A2(_09464_),
    .B1(_09489_),
    .X(_09490_));
 sky130_fd_sc_hd__nand3_1 _16420_ (.A(_09463_),
    .B(_09464_),
    .C(_09489_),
    .Y(_09491_));
 sky130_fd_sc_hd__nand2_1 _16421_ (.A(_09490_),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__xnor2_1 _16422_ (.A(_09462_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__or2_1 _16423_ (.A(_09425_),
    .B(_09427_),
    .X(_09494_));
 sky130_fd_sc_hd__a21o_1 _16424_ (.A1(_09374_),
    .A2(_09383_),
    .B1(_09381_),
    .X(_09495_));
 sky130_fd_sc_hd__or2_1 _16425_ (.A(_09388_),
    .B(_09394_),
    .X(_09496_));
 sky130_fd_sc_hd__and2_1 _16426_ (.A(_09388_),
    .B(_09394_),
    .X(_09497_));
 sky130_fd_sc_hd__a21o_1 _16427_ (.A1(_09387_),
    .A2(_09496_),
    .B1(_09497_),
    .X(_09498_));
 sky130_fd_sc_hd__nor2_1 _16428_ (.A(_08125_),
    .B(_08649_),
    .Y(_09499_));
 sky130_fd_sc_hd__nor2_1 _16429_ (.A(_08148_),
    .B(_09369_),
    .Y(_09500_));
 sky130_fd_sc_hd__xnor2_1 _16430_ (.A(_09499_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__or3_1 _16431_ (.A(_09252_),
    .B(_08524_),
    .C(_09501_),
    .X(_09502_));
 sky130_fd_sc_hd__buf_2 _16432_ (.A(_09252_),
    .X(_09503_));
 sky130_fd_sc_hd__o21ai_1 _16433_ (.A1(_09503_),
    .A2(_09132_),
    .B1(_09501_),
    .Y(_09504_));
 sky130_fd_sc_hd__and2_1 _16434_ (.A(_09502_),
    .B(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__clkbuf_4 _16435_ (.A(_08325_),
    .X(_09506_));
 sky130_fd_sc_hd__nor2_1 _16436_ (.A(_09506_),
    .B(_08411_),
    .Y(_09507_));
 sky130_fd_sc_hd__o22a_1 _16437_ (.A1(_08797_),
    .A2(_08411_),
    .B1(_08378_),
    .B2(_09506_),
    .X(_09508_));
 sky130_fd_sc_hd__a21oi_1 _16438_ (.A1(_09375_),
    .A2(_09507_),
    .B1(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__nor2_1 _16439_ (.A(_09140_),
    .B(_08387_),
    .Y(_09510_));
 sky130_fd_sc_hd__xnor2_1 _16440_ (.A(_09509_),
    .B(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__clkbuf_4 _16441_ (.A(_09140_),
    .X(_09512_));
 sky130_fd_sc_hd__nand2_1 _16442_ (.A(_09258_),
    .B(_09375_),
    .Y(_09513_));
 sky130_fd_sc_hd__o31a_1 _16443_ (.A1(_08351_),
    .A2(_09512_),
    .A3(_09376_),
    .B1(_09513_),
    .X(_09514_));
 sky130_fd_sc_hd__nor2_1 _16444_ (.A(_09511_),
    .B(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand2_1 _16445_ (.A(_09511_),
    .B(_09514_),
    .Y(_09516_));
 sky130_fd_sc_hd__and2b_1 _16446_ (.A_N(_09515_),
    .B(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__xnor2_1 _16447_ (.A(_09505_),
    .B(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__xor2_1 _16448_ (.A(_09498_),
    .B(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__xnor2_1 _16449_ (.A(_09495_),
    .B(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__a21bo_1 _16450_ (.A1(_09390_),
    .A2(_09391_),
    .B1_N(_09389_),
    .X(_09521_));
 sky130_fd_sc_hd__nor2_1 _16451_ (.A(_08941_),
    .B(_09170_),
    .Y(_09522_));
 sky130_fd_sc_hd__a22o_1 _16452_ (.A1(_09522_),
    .A2(_09399_),
    .B1(_09400_),
    .B2(_09397_),
    .X(_09523_));
 sky130_fd_sc_hd__nor2_1 _16453_ (.A(_08876_),
    .B(_08427_),
    .Y(_09524_));
 sky130_fd_sc_hd__a21oi_1 _16454_ (.A1(_08454_),
    .A2(_09025_),
    .B1(_08875_),
    .Y(_09525_));
 sky130_fd_sc_hd__xnor2_1 _16455_ (.A(_09524_),
    .B(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__nor2_1 _16456_ (.A(_08394_),
    .B(_08409_),
    .Y(_09527_));
 sky130_fd_sc_hd__xnor2_1 _16457_ (.A(_09526_),
    .B(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__xor2_1 _16458_ (.A(_09523_),
    .B(_09528_),
    .X(_09529_));
 sky130_fd_sc_hd__xor2_1 _16459_ (.A(_09521_),
    .B(_09529_),
    .X(_09530_));
 sky130_fd_sc_hd__or3b_1 _16460_ (.A(_08941_),
    .B(_09403_),
    .C_N(_09399_),
    .X(_09531_));
 sky130_fd_sc_hd__and2_1 _16461_ (.A(_09180_),
    .B(_09287_),
    .X(_09532_));
 sky130_fd_sc_hd__buf_2 _16462_ (.A(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__clkbuf_4 _16463_ (.A(_09403_),
    .X(_09534_));
 sky130_fd_sc_hd__o22ai_2 _16464_ (.A1(_08941_),
    .A2(_09533_),
    .B1(_09534_),
    .B2(_08911_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand2_1 _16465_ (.A(_09531_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__nor2_1 _16466_ (.A(_08360_),
    .B(_09170_),
    .Y(_09537_));
 sky130_fd_sc_hd__xnor2_1 _16467_ (.A(_09536_),
    .B(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__inv_2 _16468_ (.A(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_09539_));
 sky130_fd_sc_hd__mux2_2 _16469_ (.A0(_09539_),
    .A1(_09409_),
    .S(_08130_),
    .X(_09540_));
 sky130_fd_sc_hd__nor2_1 _16470_ (.A(_08928_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__or4_1 _16471_ (.A(_07988_),
    .B(_07999_),
    .C(_08430_),
    .D(_09174_),
    .X(_09542_));
 sky130_fd_sc_hd__or3_1 _16472_ (.A(_08003_),
    .B(_08005_),
    .C(_09542_),
    .X(_09543_));
 sky130_fd_sc_hd__o21ai_1 _16473_ (.A1(_08003_),
    .A2(_09542_),
    .B1(_08005_),
    .Y(_09544_));
 sky130_fd_sc_hd__a31o_1 _16474_ (.A1(_08429_),
    .A2(_09543_),
    .A3(_09544_),
    .B1(_08434_),
    .X(_09545_));
 sky130_fd_sc_hd__or3b_1 _16475_ (.A(_08319_),
    .B(_09545_),
    .C_N(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_09546_));
 sky130_fd_sc_hd__nor2_1 _16476_ (.A(_08830_),
    .B(_09406_),
    .Y(_09547_));
 sky130_fd_sc_hd__xnor2_1 _16477_ (.A(_09546_),
    .B(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__xnor2_1 _16478_ (.A(_09541_),
    .B(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand2_1 _16479_ (.A(_09408_),
    .B(_09411_),
    .Y(_09550_));
 sky130_fd_sc_hd__xnor2_1 _16480_ (.A(_09549_),
    .B(_09550_),
    .Y(_09551_));
 sky130_fd_sc_hd__xnor2_1 _16481_ (.A(_09538_),
    .B(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__and2_1 _16482_ (.A(_09415_),
    .B(_09417_),
    .X(_09553_));
 sky130_fd_sc_hd__xor2_1 _16483_ (.A(_09552_),
    .B(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__xnor2_1 _16484_ (.A(_09530_),
    .B(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__a21boi_1 _16485_ (.A1(_09396_),
    .A2(_09422_),
    .B1_N(_09421_),
    .Y(_09556_));
 sky130_fd_sc_hd__xor2_1 _16486_ (.A(_09555_),
    .B(_09556_),
    .X(_09557_));
 sky130_fd_sc_hd__xnor2_1 _16487_ (.A(_09520_),
    .B(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__a21oi_1 _16488_ (.A1(_09494_),
    .A2(_09429_),
    .B1(_09558_),
    .Y(_09559_));
 sky130_fd_sc_hd__and3_1 _16489_ (.A(_09494_),
    .B(_09429_),
    .C(_09558_),
    .X(_09560_));
 sky130_fd_sc_hd__nor2_1 _16490_ (.A(_09559_),
    .B(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__xnor2_1 _16491_ (.A(_09493_),
    .B(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__a21oi_1 _16492_ (.A1(_09365_),
    .A2(_09435_),
    .B1(_09433_),
    .Y(_09563_));
 sky130_fd_sc_hd__or2_1 _16493_ (.A(_09562_),
    .B(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__nand2_1 _16494_ (.A(_09562_),
    .B(_09563_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand2_1 _16495_ (.A(_09564_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__xor2_1 _16496_ (.A(_09461_),
    .B(_09566_),
    .X(_09567_));
 sky130_fd_sc_hd__xnor2_2 _16497_ (.A(_09459_),
    .B(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__xnor2_4 _16498_ (.A(_09442_),
    .B(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__xnor2_4 _16499_ (.A(_09457_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__mux2_1 _16500_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_08115_),
    .X(_09571_));
 sky130_fd_sc_hd__nor2_1 _16501_ (.A(_09570_),
    .B(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__and2_1 _16502_ (.A(_09570_),
    .B(_09571_),
    .X(_09573_));
 sky130_fd_sc_hd__nor2_1 _16503_ (.A(_09572_),
    .B(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__xor2_1 _16504_ (.A(_09102_),
    .B(_09574_),
    .X(_09575_));
 sky130_fd_sc_hd__xnor2_1 _16505_ (.A(_09455_),
    .B(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__or2_1 _16506_ (.A(\rbzero.texu_hot[4] ),
    .B(_08120_),
    .X(_09577_));
 sky130_fd_sc_hd__o211a_1 _16507_ (.A1(_08429_),
    .A2(_09576_),
    .B1(_09577_),
    .C1(_04478_),
    .X(_00470_));
 sky130_fd_sc_hd__o21ba_1 _16508_ (.A1(_09455_),
    .A2(_09572_),
    .B1_N(_09573_),
    .X(_09578_));
 sky130_fd_sc_hd__inv_2 _16509_ (.A(_09569_),
    .Y(_09579_));
 sky130_fd_sc_hd__nand2_1 _16510_ (.A(_09442_),
    .B(_09568_),
    .Y(_09580_));
 sky130_fd_sc_hd__a21bo_1 _16511_ (.A1(_09457_),
    .A2(_09579_),
    .B1_N(_09580_),
    .X(_09581_));
 sky130_fd_sc_hd__or2b_2 _16512_ (.A(_09567_),
    .B_N(_09459_),
    .X(_09582_));
 sky130_fd_sc_hd__or2b_1 _16513_ (.A(_09566_),
    .B_N(_09461_),
    .X(_09583_));
 sky130_fd_sc_hd__or2b_1 _16514_ (.A(_09492_),
    .B_N(_09462_),
    .X(_09584_));
 sky130_fd_sc_hd__or2b_1 _16515_ (.A(_09465_),
    .B_N(_09471_),
    .X(_09585_));
 sky130_fd_sc_hd__a21oi_1 _16516_ (.A1(_09490_),
    .A2(_09584_),
    .B1(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__and3_1 _16517_ (.A(_09585_),
    .B(_09490_),
    .C(_09584_),
    .X(_09587_));
 sky130_fd_sc_hd__nor2_1 _16518_ (.A(_09586_),
    .B(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__nand2_4 _16519_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_08523_),
    .Y(_09589_));
 sky130_fd_sc_hd__or2_1 _16520_ (.A(_08137_),
    .B(_09589_),
    .X(_09590_));
 sky130_fd_sc_hd__xnor2_1 _16521_ (.A(_09588_),
    .B(_09590_),
    .Y(_09591_));
 sky130_fd_sc_hd__a21o_1 _16522_ (.A1(_09472_),
    .A2(_09488_),
    .B1(_09486_),
    .X(_09592_));
 sky130_fd_sc_hd__or2b_1 _16523_ (.A(_09518_),
    .B_N(_09498_),
    .X(_09593_));
 sky130_fd_sc_hd__or2b_1 _16524_ (.A(_09519_),
    .B_N(_09495_),
    .X(_09594_));
 sky130_fd_sc_hd__nor2_1 _16525_ (.A(_08602_),
    .B(_09342_),
    .Y(_09595_));
 sky130_fd_sc_hd__o22ai_1 _16526_ (.A1(_09128_),
    .A2(_09110_),
    .B1(_09226_),
    .B2(_08935_),
    .Y(_09596_));
 sky130_fd_sc_hd__o31a_1 _16527_ (.A1(_09128_),
    .A2(_09226_),
    .A3(_09474_),
    .B1(_09596_),
    .X(_09597_));
 sky130_fd_sc_hd__nand2_1 _16528_ (.A(_09595_),
    .B(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__or2_1 _16529_ (.A(_09595_),
    .B(_09597_),
    .X(_09599_));
 sky130_fd_sc_hd__nand2_1 _16530_ (.A(_09598_),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__nor2_1 _16531_ (.A(_08285_),
    .B(_09228_),
    .Y(_09601_));
 sky130_fd_sc_hd__nand2_1 _16532_ (.A(_09601_),
    .B(_09595_),
    .Y(_09602_));
 sky130_fd_sc_hd__o31a_1 _16533_ (.A1(_08598_),
    .A2(_09467_),
    .A3(_09469_),
    .B1(_09602_),
    .X(_09603_));
 sky130_fd_sc_hd__xor2_1 _16534_ (.A(_09600_),
    .B(_09603_),
    .X(_09604_));
 sky130_fd_sc_hd__buf_4 _16535_ (.A(_09469_),
    .X(_09605_));
 sky130_fd_sc_hd__nor2_1 _16536_ (.A(_08285_),
    .B(_09605_),
    .Y(_09606_));
 sky130_fd_sc_hd__xor2_1 _16537_ (.A(_09604_),
    .B(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__o21ai_1 _16538_ (.A1(_09474_),
    .A2(_09475_),
    .B1(_09477_),
    .Y(_09608_));
 sky130_fd_sc_hd__a21bo_1 _16539_ (.A1(_09499_),
    .A2(_09500_),
    .B1_N(_09502_),
    .X(_09609_));
 sky130_fd_sc_hd__o22a_1 _16540_ (.A1(_09369_),
    .A2(_08524_),
    .B1(_08599_),
    .B2(_09252_),
    .X(_09610_));
 sky130_fd_sc_hd__or2_1 _16541_ (.A(_08176_),
    .B(_08599_),
    .X(_09611_));
 sky130_fd_sc_hd__or3_1 _16542_ (.A(_09252_),
    .B(_08524_),
    .C(_09611_),
    .X(_09612_));
 sky130_fd_sc_hd__and2b_1 _16543_ (.A_N(_09610_),
    .B(_09612_),
    .X(_09613_));
 sky130_fd_sc_hd__xnor2_1 _16544_ (.A(_09476_),
    .B(_09613_),
    .Y(_09614_));
 sky130_fd_sc_hd__and2_1 _16545_ (.A(_09609_),
    .B(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__or2_1 _16546_ (.A(_09609_),
    .B(_09614_),
    .X(_09616_));
 sky130_fd_sc_hd__and2b_1 _16547_ (.A_N(_09615_),
    .B(_09616_),
    .X(_09617_));
 sky130_fd_sc_hd__xnor2_1 _16548_ (.A(_09608_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__a21oi_1 _16549_ (.A1(_09473_),
    .A2(_09483_),
    .B1(_09481_),
    .Y(_09619_));
 sky130_fd_sc_hd__nor2_1 _16550_ (.A(_09618_),
    .B(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__and2_1 _16551_ (.A(_09618_),
    .B(_09619_),
    .X(_09621_));
 sky130_fd_sc_hd__nor2_1 _16552_ (.A(_09620_),
    .B(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__xnor2_1 _16553_ (.A(_09607_),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__a21o_1 _16554_ (.A1(_09593_),
    .A2(_09594_),
    .B1(_09623_),
    .X(_09624_));
 sky130_fd_sc_hd__nand3_1 _16555_ (.A(_09593_),
    .B(_09594_),
    .C(_09623_),
    .Y(_09625_));
 sky130_fd_sc_hd__nand2_1 _16556_ (.A(_09624_),
    .B(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__xnor2_1 _16557_ (.A(_09592_),
    .B(_09626_),
    .Y(_09627_));
 sky130_fd_sc_hd__a21o_1 _16558_ (.A1(_09505_),
    .A2(_09516_),
    .B1(_09515_),
    .X(_09628_));
 sky130_fd_sc_hd__nand2_1 _16559_ (.A(_09523_),
    .B(_09528_),
    .Y(_09629_));
 sky130_fd_sc_hd__a21bo_1 _16560_ (.A1(_09521_),
    .A2(_09529_),
    .B1_N(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__or2_1 _16561_ (.A(_08286_),
    .B(_08649_),
    .X(_09631_));
 sky130_fd_sc_hd__or4_1 _16562_ (.A(_08126_),
    .B(_08546_),
    .C(_08378_),
    .D(_08385_),
    .X(_09632_));
 sky130_fd_sc_hd__o22ai_1 _16563_ (.A1(_09140_),
    .A2(_08378_),
    .B1(_08385_),
    .B2(_08127_),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2_1 _16564_ (.A(_09632_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__xor2_1 _16565_ (.A(_09631_),
    .B(_09634_),
    .X(_09635_));
 sky130_fd_sc_hd__nor2_2 _16566_ (.A(_08296_),
    .B(_08427_),
    .Y(_09636_));
 sky130_fd_sc_hd__o22ai_1 _16567_ (.A1(_08797_),
    .A2(_08409_),
    .B1(_08427_),
    .B2(_08394_),
    .Y(_09637_));
 sky130_fd_sc_hd__a21boi_1 _16568_ (.A1(_09527_),
    .A2(_09636_),
    .B1_N(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__xnor2_1 _16569_ (.A(_09507_),
    .B(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__a22oi_1 _16570_ (.A1(_09375_),
    .A2(_09507_),
    .B1(_09509_),
    .B2(_09510_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2_1 _16571_ (.A(_09639_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__nand2_1 _16572_ (.A(_09639_),
    .B(_09640_),
    .Y(_09642_));
 sky130_fd_sc_hd__and2b_1 _16573_ (.A_N(_09641_),
    .B(_09642_),
    .X(_09643_));
 sky130_fd_sc_hd__xnor2_1 _16574_ (.A(_09635_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__xor2_1 _16575_ (.A(_09630_),
    .B(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__xnor2_1 _16576_ (.A(_09628_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__buf_2 _16577_ (.A(_08394_),
    .X(_09647_));
 sky130_fd_sc_hd__or3_1 _16578_ (.A(_09647_),
    .B(_08409_),
    .C(_09526_),
    .X(_09648_));
 sky130_fd_sc_hd__a21bo_1 _16579_ (.A1(_09524_),
    .A2(_09525_),
    .B1_N(_09648_),
    .X(_09649_));
 sky130_fd_sc_hd__a21bo_1 _16580_ (.A1(_09535_),
    .A2(_09537_),
    .B1_N(_09531_),
    .X(_09650_));
 sky130_fd_sc_hd__and2_1 _16581_ (.A(_08247_),
    .B(_09026_),
    .X(_09651_));
 sky130_fd_sc_hd__a21o_1 _16582_ (.A1(_09286_),
    .A2(_09287_),
    .B1(_08359_),
    .X(_09652_));
 sky130_fd_sc_hd__a21oi_1 _16583_ (.A1(_09295_),
    .A2(_09168_),
    .B1(_08352_),
    .Y(_09653_));
 sky130_fd_sc_hd__xnor2_1 _16584_ (.A(_09652_),
    .B(_09653_),
    .Y(_09654_));
 sky130_fd_sc_hd__xor2_1 _16585_ (.A(_09651_),
    .B(_09654_),
    .X(_09655_));
 sky130_fd_sc_hd__and2_1 _16586_ (.A(_09650_),
    .B(_09655_),
    .X(_09656_));
 sky130_fd_sc_hd__nor2_1 _16587_ (.A(_09650_),
    .B(_09655_),
    .Y(_09657_));
 sky130_fd_sc_hd__nor2_1 _16588_ (.A(_09656_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__xor2_2 _16589_ (.A(_09649_),
    .B(_09658_),
    .X(_09659_));
 sky130_fd_sc_hd__or2_1 _16590_ (.A(_08399_),
    .B(_09403_),
    .X(_09660_));
 sky130_fd_sc_hd__clkinv_2 _16591_ (.A(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_09661_));
 sky130_fd_sc_hd__mux2_2 _16592_ (.A0(_09661_),
    .A1(_09406_),
    .S(_08130_),
    .X(_09662_));
 sky130_fd_sc_hd__clkbuf_4 _16593_ (.A(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__nor4_1 _16594_ (.A(_08911_),
    .B(_08928_),
    .C(_09540_),
    .D(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__o22a_1 _16595_ (.A1(_08412_),
    .A2(_09540_),
    .B1(_09662_),
    .B2(_08420_),
    .X(_09665_));
 sky130_fd_sc_hd__or3_1 _16596_ (.A(_09660_),
    .B(_09664_),
    .C(_09665_),
    .X(_09666_));
 sky130_fd_sc_hd__o21ai_1 _16597_ (.A1(_09664_),
    .A2(_09665_),
    .B1(_09660_),
    .Y(_09667_));
 sky130_fd_sc_hd__and2_1 _16598_ (.A(_09666_),
    .B(_09667_),
    .X(_09668_));
 sky130_fd_sc_hd__nor2_2 _16599_ (.A(_06135_),
    .B(_08319_),
    .Y(_09669_));
 sky130_fd_sc_hd__or4_1 _16600_ (.A(_08003_),
    .B(_08005_),
    .C(_08008_),
    .D(_09542_),
    .X(_09670_));
 sky130_fd_sc_hd__a21o_1 _16601_ (.A1(_08429_),
    .A2(_09670_),
    .B1(_08434_),
    .X(_09671_));
 sky130_fd_sc_hd__or3b_4 _16602_ (.A(_08319_),
    .B(_09671_),
    .C_N(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_09672_));
 sky130_fd_sc_hd__mux2_1 _16603_ (.A0(_06135_),
    .A1(_09669_),
    .S(_09672_),
    .X(_09673_));
 sky130_fd_sc_hd__nand2_1 _16604_ (.A(\rbzero.wall_tracer.stepDistY[9] ),
    .B(_08406_),
    .Y(_09674_));
 sky130_fd_sc_hd__a21oi_1 _16605_ (.A1(_09674_),
    .A2(_09545_),
    .B1(_08830_),
    .Y(_09675_));
 sky130_fd_sc_hd__xnor2_2 _16606_ (.A(_09673_),
    .B(_09675_),
    .Y(_09676_));
 sky130_fd_sc_hd__and2b_1 _16607_ (.A_N(_09546_),
    .B(_09547_),
    .X(_09677_));
 sky130_fd_sc_hd__a21o_1 _16608_ (.A1(_09541_),
    .A2(_09548_),
    .B1(_09677_),
    .X(_09678_));
 sky130_fd_sc_hd__xnor2_2 _16609_ (.A(_09676_),
    .B(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__xnor2_2 _16610_ (.A(_09668_),
    .B(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__and2b_1 _16611_ (.A_N(_09549_),
    .B(_09550_),
    .X(_09681_));
 sky130_fd_sc_hd__a21o_1 _16612_ (.A1(_09538_),
    .A2(_09551_),
    .B1(_09681_),
    .X(_09682_));
 sky130_fd_sc_hd__xnor2_2 _16613_ (.A(_09680_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__xnor2_2 _16614_ (.A(_09659_),
    .B(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__nor2_1 _16615_ (.A(_09552_),
    .B(_09553_),
    .Y(_09685_));
 sky130_fd_sc_hd__a21o_1 _16616_ (.A1(_09530_),
    .A2(_09554_),
    .B1(_09685_),
    .X(_09686_));
 sky130_fd_sc_hd__xnor2_1 _16617_ (.A(_09684_),
    .B(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__xnor2_2 _16618_ (.A(_09646_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__nor2_1 _16619_ (.A(_09555_),
    .B(_09556_),
    .Y(_09689_));
 sky130_fd_sc_hd__a21oi_1 _16620_ (.A1(_09520_),
    .A2(_09557_),
    .B1(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__nor2_1 _16621_ (.A(_09688_),
    .B(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__nand2_1 _16622_ (.A(_09688_),
    .B(_09690_),
    .Y(_09692_));
 sky130_fd_sc_hd__and2b_1 _16623_ (.A_N(_09691_),
    .B(_09692_),
    .X(_09693_));
 sky130_fd_sc_hd__xnor2_1 _16624_ (.A(_09627_),
    .B(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__a21oi_1 _16625_ (.A1(_09493_),
    .A2(_09561_),
    .B1(_09559_),
    .Y(_09695_));
 sky130_fd_sc_hd__xor2_1 _16626_ (.A(_09694_),
    .B(_09695_),
    .X(_09696_));
 sky130_fd_sc_hd__xnor2_1 _16627_ (.A(_09591_),
    .B(_09696_),
    .Y(_09697_));
 sky130_fd_sc_hd__a21oi_1 _16628_ (.A1(_09564_),
    .A2(_09583_),
    .B1(_09697_),
    .Y(_09698_));
 sky130_fd_sc_hd__and3_1 _16629_ (.A(_09564_),
    .B(_09583_),
    .C(_09697_),
    .X(_09699_));
 sky130_fd_sc_hd__or2_2 _16630_ (.A(_09698_),
    .B(_09699_),
    .X(_09700_));
 sky130_fd_sc_hd__xor2_4 _16631_ (.A(_09582_),
    .B(_09700_),
    .X(_09701_));
 sky130_fd_sc_hd__xnor2_4 _16632_ (.A(_09581_),
    .B(_09701_),
    .Y(_09702_));
 sky130_fd_sc_hd__mux2_1 _16633_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_08115_),
    .X(_09703_));
 sky130_fd_sc_hd__xor2_1 _16634_ (.A(_09102_),
    .B(_09703_),
    .X(_09704_));
 sky130_fd_sc_hd__xnor2_1 _16635_ (.A(_09702_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__xnor2_1 _16636_ (.A(_09578_),
    .B(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__or2_1 _16637_ (.A(\rbzero.texu_hot[5] ),
    .B(_08120_),
    .X(_09707_));
 sky130_fd_sc_hd__o211a_1 _16638_ (.A1(_08429_),
    .A2(_09706_),
    .B1(_09707_),
    .C1(_04478_),
    .X(_00471_));
 sky130_fd_sc_hd__and4_1 _16639_ (.A(_04484_),
    .B(_04666_),
    .C(_05077_),
    .D(_04692_),
    .X(_09708_));
 sky130_fd_sc_hd__buf_4 _16640_ (.A(_09708_),
    .X(_09709_));
 sky130_fd_sc_hd__or2_1 _16641_ (.A(_04094_),
    .B(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__buf_2 _16642_ (.A(_09710_),
    .X(_09711_));
 sky130_fd_sc_hd__nor2_1 _16643_ (.A(_04012_),
    .B(_09711_),
    .Y(_00472_));
 sky130_fd_sc_hd__clkbuf_4 _16644_ (.A(_08091_),
    .X(_09712_));
 sky130_fd_sc_hd__and3_1 _16645_ (.A(_09712_),
    .B(_04616_),
    .C(_04617_),
    .X(_09713_));
 sky130_fd_sc_hd__clkbuf_1 _16646_ (.A(_09713_),
    .X(_00473_));
 sky130_fd_sc_hd__a21o_1 _16647_ (.A1(_04585_),
    .A2(_04012_),
    .B1(_04587_),
    .X(_09714_));
 sky130_fd_sc_hd__and3b_1 _16648_ (.A_N(_04665_),
    .B(_09714_),
    .C(_08092_),
    .X(_09715_));
 sky130_fd_sc_hd__clkbuf_1 _16649_ (.A(_09715_),
    .X(_00474_));
 sky130_fd_sc_hd__nor2_1 _16650_ (.A(net65),
    .B(_05200_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _16651_ (.A(_05221_),
    .B(_09711_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _16652_ (.A(_05225_),
    .B(_09711_),
    .Y(_00477_));
 sky130_fd_sc_hd__nor2_1 _16653_ (.A(_05204_),
    .B(_09711_),
    .Y(_00478_));
 sky130_fd_sc_hd__nor2_4 _16654_ (.A(_04094_),
    .B(_09709_),
    .Y(_09716_));
 sky130_fd_sc_hd__and2_1 _16655_ (.A(_05229_),
    .B(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__clkbuf_1 _16656_ (.A(_09717_),
    .X(_00479_));
 sky130_fd_sc_hd__and3_1 _16657_ (.A(_04017_),
    .B(_04665_),
    .C(_05173_),
    .X(_09718_));
 sky130_fd_sc_hd__a21o_1 _16658_ (.A1(_04665_),
    .A2(_05173_),
    .B1(_04017_),
    .X(_09719_));
 sky130_fd_sc_hd__and3b_1 _16659_ (.A_N(_09718_),
    .B(_09719_),
    .C(_09716_),
    .X(_09720_));
 sky130_fd_sc_hd__clkbuf_1 _16660_ (.A(_09720_),
    .X(_00480_));
 sky130_fd_sc_hd__a21oi_1 _16661_ (.A1(_04018_),
    .A2(_09718_),
    .B1(_09711_),
    .Y(_09721_));
 sky130_fd_sc_hd__o21a_1 _16662_ (.A1(_04018_),
    .A2(_09718_),
    .B1(_09721_),
    .X(_00481_));
 sky130_fd_sc_hd__and3_1 _16663_ (.A(_04471_),
    .B(_04687_),
    .C(_09709_),
    .X(_09722_));
 sky130_fd_sc_hd__nor2_1 _16664_ (.A(_08111_),
    .B(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__clkbuf_8 _16665_ (.A(_09723_),
    .X(_09724_));
 sky130_fd_sc_hd__buf_4 _16666_ (.A(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__nand3_1 _16667_ (.A(_04471_),
    .B(_04687_),
    .C(_09709_),
    .Y(_09726_));
 sky130_fd_sc_hd__nor2_2 _16668_ (.A(_08111_),
    .B(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__clkbuf_8 _16669_ (.A(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__clkbuf_4 _16670_ (.A(_09728_),
    .X(_09729_));
 sky130_fd_sc_hd__a22o_1 _16671_ (.A1(_04702_),
    .A2(_09725_),
    .B1(_09729_),
    .B2(_08115_),
    .X(_00482_));
 sky130_fd_sc_hd__a22o_1 _16672_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_09725_),
    .B1(_09729_),
    .B2(_07897_),
    .X(_00483_));
 sky130_fd_sc_hd__or2_4 _16673_ (.A(_08111_),
    .B(_09726_),
    .X(_09730_));
 sky130_fd_sc_hd__buf_6 _16674_ (.A(_09730_),
    .X(_09731_));
 sky130_fd_sc_hd__a2bb2o_1 _16675_ (.A1_N(_07911_),
    .A2_N(_09731_),
    .B1(_09725_),
    .B2(\rbzero.row_render.size[1] ),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _16676_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_09725_),
    .B1(_09729_),
    .B2(_07920_),
    .X(_00485_));
 sky130_fd_sc_hd__a2bb2o_1 _16677_ (.A1_N(_07931_),
    .A2_N(_09731_),
    .B1(_09725_),
    .B2(\rbzero.row_render.size[3] ),
    .X(_00486_));
 sky130_fd_sc_hd__clkbuf_4 _16678_ (.A(_09724_),
    .X(_09732_));
 sky130_fd_sc_hd__a22o_1 _16679_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_09732_),
    .B1(_09729_),
    .B2(_07940_),
    .X(_00487_));
 sky130_fd_sc_hd__a22o_1 _16680_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_09732_),
    .B1(_09729_),
    .B2(_07948_),
    .X(_00488_));
 sky130_fd_sc_hd__a22o_1 _16681_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_09732_),
    .B1(_09729_),
    .B2(_07953_),
    .X(_00489_));
 sky130_fd_sc_hd__a22o_1 _16682_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_09732_),
    .B1(_09729_),
    .B2(_07960_),
    .X(_00490_));
 sky130_fd_sc_hd__a22o_1 _16683_ (.A1(\rbzero.row_render.size[8] ),
    .A2(_09732_),
    .B1(_09729_),
    .B2(_07966_),
    .X(_00491_));
 sky130_fd_sc_hd__a22o_1 _16684_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_09732_),
    .B1(_09729_),
    .B2(_07971_),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _16685_ (.A1(\rbzero.row_render.size[10] ),
    .A2(_09732_),
    .B1(_09729_),
    .B2(_07976_),
    .X(_00493_));
 sky130_fd_sc_hd__clkbuf_4 _16686_ (.A(_09728_),
    .X(_09733_));
 sky130_fd_sc_hd__a22o_1 _16687_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_09732_),
    .B1(_09733_),
    .B2(\rbzero.texu_hot[0] ),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _16688_ (.A1(\rbzero.row_render.texu[1] ),
    .A2(_09732_),
    .B1(_09733_),
    .B2(\rbzero.texu_hot[1] ),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _16689_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_09732_),
    .B1(_09733_),
    .B2(\rbzero.texu_hot[2] ),
    .X(_00496_));
 sky130_fd_sc_hd__clkbuf_4 _16690_ (.A(_09724_),
    .X(_09734_));
 sky130_fd_sc_hd__a22o_1 _16691_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(_09734_),
    .B1(_09733_),
    .B2(\rbzero.texu_hot[3] ),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _16692_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_09734_),
    .B1(_09733_),
    .B2(\rbzero.texu_hot[4] ),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_1 _16693_ (.A1(\rbzero.traced_texa[-11] ),
    .A2(_09734_),
    .B1(_09733_),
    .B2(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _16694_ (.A1(\rbzero.traced_texa[-10] ),
    .A2(_09734_),
    .B1(_09733_),
    .B2(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _16695_ (.A1(\rbzero.traced_texa[-9] ),
    .A2(_09734_),
    .B1(_09733_),
    .B2(net515),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_1 _16696_ (.A1(\rbzero.traced_texa[-8] ),
    .A2(_09734_),
    .B1(_09733_),
    .B2(net516),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _16697_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(_09734_),
    .B1(_09733_),
    .B2(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(_00503_));
 sky130_fd_sc_hd__clkbuf_4 _16698_ (.A(_09728_),
    .X(_09735_));
 sky130_fd_sc_hd__a22o_1 _16699_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(_09734_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _16700_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(_09734_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _16701_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(_09734_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(_00506_));
 sky130_fd_sc_hd__buf_2 _16702_ (.A(_09724_),
    .X(_09736_));
 sky130_fd_sc_hd__a22o_1 _16703_ (.A1(\rbzero.traced_texa[-3] ),
    .A2(_09736_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _16704_ (.A1(\rbzero.traced_texa[-2] ),
    .A2(_09736_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _16705_ (.A1(\rbzero.traced_texa[-1] ),
    .A2(_09736_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_00509_));
 sky130_fd_sc_hd__a22o_1 _16706_ (.A1(\rbzero.traced_texa[0] ),
    .A2(_09736_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_00510_));
 sky130_fd_sc_hd__a22o_1 _16707_ (.A1(\rbzero.traced_texa[1] ),
    .A2(_09736_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_00511_));
 sky130_fd_sc_hd__a22o_1 _16708_ (.A1(\rbzero.traced_texa[2] ),
    .A2(_09736_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _16709_ (.A1(\rbzero.traced_texa[3] ),
    .A2(_09736_),
    .B1(_09735_),
    .B2(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(_00513_));
 sky130_fd_sc_hd__buf_2 _16710_ (.A(_09728_),
    .X(_09737_));
 sky130_fd_sc_hd__a22o_1 _16711_ (.A1(\rbzero.traced_texa[4] ),
    .A2(_09736_),
    .B1(_09737_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_1 _16712_ (.A1(\rbzero.traced_texa[5] ),
    .A2(_09736_),
    .B1(_09737_),
    .B2(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _16713_ (.A1(\rbzero.traced_texa[6] ),
    .A2(_09736_),
    .B1(_09737_),
    .B2(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_00516_));
 sky130_fd_sc_hd__buf_6 _16714_ (.A(_09724_),
    .X(_09738_));
 sky130_fd_sc_hd__a22o_1 _16715_ (.A1(\rbzero.traced_texa[7] ),
    .A2(_09738_),
    .B1(_09737_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _16716_ (.A1(\rbzero.traced_texa[8] ),
    .A2(_09738_),
    .B1(_09737_),
    .B2(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_00518_));
 sky130_fd_sc_hd__a22o_1 _16717_ (.A1(\rbzero.traced_texa[9] ),
    .A2(_09738_),
    .B1(_09737_),
    .B2(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_00519_));
 sky130_fd_sc_hd__a22o_1 _16718_ (.A1(\rbzero.traced_texa[10] ),
    .A2(_09738_),
    .B1(_09737_),
    .B2(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _16719_ (.A0(\rbzero.wall_hot[0] ),
    .A1(\rbzero.row_render.wall[0] ),
    .S(_09730_),
    .X(_09739_));
 sky130_fd_sc_hd__clkbuf_1 _16720_ (.A(_09739_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _16721_ (.A0(\rbzero.wall_hot[1] ),
    .A1(\rbzero.row_render.wall[1] ),
    .S(_09730_),
    .X(_09740_));
 sky130_fd_sc_hd__clkbuf_1 _16722_ (.A(_09740_),
    .X(_00522_));
 sky130_fd_sc_hd__o21a_1 _16723_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(\rbzero.wall_tracer.mapX[5] ),
    .B1(_09100_),
    .X(_09741_));
 sky130_fd_sc_hd__xor2_1 _16724_ (.A(\rbzero.wall_tracer.mapX[5] ),
    .B(_09099_),
    .X(_09742_));
 sky130_fd_sc_hd__xnor2_1 _16725_ (.A(_06116_),
    .B(_09099_),
    .Y(_09743_));
 sky130_fd_sc_hd__and2_1 _16726_ (.A(_06105_),
    .B(_09099_),
    .X(_09744_));
 sky130_fd_sc_hd__xnor2_1 _16727_ (.A(_06122_),
    .B(_08178_),
    .Y(_09745_));
 sky130_fd_sc_hd__and2_1 _16728_ (.A(_06108_),
    .B(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__a21o_1 _16729_ (.A1(_06126_),
    .A2(_09099_),
    .B1(_09746_),
    .X(_09747_));
 sky130_fd_sc_hd__and2_1 _16730_ (.A(_06117_),
    .B(_08178_),
    .X(_09748_));
 sky130_fd_sc_hd__nor2_1 _16731_ (.A(_06117_),
    .B(_09099_),
    .Y(_09749_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_09748_),
    .B(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__a21o_1 _16733_ (.A1(_09747_),
    .A2(_09750_),
    .B1(_09748_),
    .X(_09751_));
 sky130_fd_sc_hd__nor2_1 _16734_ (.A(_06105_),
    .B(_09099_),
    .Y(_09752_));
 sky130_fd_sc_hd__o21ba_1 _16735_ (.A1(_09744_),
    .A2(_09751_),
    .B1_N(_09752_),
    .X(_09753_));
 sky130_fd_sc_hd__and3_1 _16736_ (.A(_09742_),
    .B(_09743_),
    .C(_09753_),
    .X(_09754_));
 sky130_fd_sc_hd__nand2_1 _16737_ (.A(\rbzero.wall_tracer.mapX[6] ),
    .B(_09099_),
    .Y(_09755_));
 sky130_fd_sc_hd__or2_1 _16738_ (.A(\rbzero.wall_tracer.mapX[6] ),
    .B(_09099_),
    .X(_09756_));
 sky130_fd_sc_hd__and2_1 _16739_ (.A(_09755_),
    .B(_09756_),
    .X(_09757_));
 sky130_fd_sc_hd__o21ai_1 _16740_ (.A1(_09741_),
    .A2(_09754_),
    .B1(_09757_),
    .Y(_09758_));
 sky130_fd_sc_hd__or3_1 _16741_ (.A(_09757_),
    .B(_09741_),
    .C(_09754_),
    .X(_09759_));
 sky130_fd_sc_hd__buf_6 _16742_ (.A(_06102_),
    .X(_09760_));
 sky130_fd_sc_hd__a21o_4 _16743_ (.A1(_08130_),
    .A2(_06252_),
    .B1(_08111_),
    .X(_09761_));
 sky130_fd_sc_hd__nor2_2 _16744_ (.A(_09760_),
    .B(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__buf_4 _16745_ (.A(_09761_),
    .X(_09763_));
 sky130_fd_sc_hd__a32o_1 _16746_ (.A1(_09758_),
    .A2(_09759_),
    .A3(_09762_),
    .B1(_09763_),
    .B2(\rbzero.wall_tracer.mapX[6] ),
    .X(_00523_));
 sky130_fd_sc_hd__xnor2_1 _16747_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(_09099_),
    .Y(_09764_));
 sky130_fd_sc_hd__a21o_1 _16748_ (.A1(_09755_),
    .A2(_09758_),
    .B1(_09764_),
    .X(_09765_));
 sky130_fd_sc_hd__nand3_1 _16749_ (.A(_09755_),
    .B(_09758_),
    .C(_09764_),
    .Y(_09766_));
 sky130_fd_sc_hd__a32o_1 _16750_ (.A1(_09762_),
    .A2(_09765_),
    .A3(_09766_),
    .B1(_09763_),
    .B2(\rbzero.wall_tracer.mapX[7] ),
    .X(_00524_));
 sky130_fd_sc_hd__clkbuf_4 _16751_ (.A(_09761_),
    .X(_09767_));
 sky130_fd_sc_hd__xor2_1 _16752_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(_09100_),
    .X(_09768_));
 sky130_fd_sc_hd__clkinv_2 _16753_ (.A(_09764_),
    .Y(_09769_));
 sky130_fd_sc_hd__and3_1 _16754_ (.A(_09757_),
    .B(_09754_),
    .C(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__o21a_1 _16755_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(\rbzero.wall_tracer.mapX[6] ),
    .B1(_09100_),
    .X(_09771_));
 sky130_fd_sc_hd__or3_1 _16756_ (.A(_09741_),
    .B(_09770_),
    .C(_09771_),
    .X(_09772_));
 sky130_fd_sc_hd__xor2_1 _16757_ (.A(_09768_),
    .B(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__a22o_1 _16758_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09767_),
    .B1(_09762_),
    .B2(_09773_),
    .X(_00525_));
 sky130_fd_sc_hd__a22o_1 _16759_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09100_),
    .B1(_09768_),
    .B2(_09772_),
    .X(_09774_));
 sky130_fd_sc_hd__xnor2_1 _16760_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(_09100_),
    .Y(_09775_));
 sky130_fd_sc_hd__xnor2_1 _16761_ (.A(_09774_),
    .B(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__a22o_1 _16762_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09767_),
    .B1(_09762_),
    .B2(_09776_),
    .X(_00526_));
 sky130_fd_sc_hd__o21a_1 _16763_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09100_),
    .B1(_09774_),
    .X(_09777_));
 sky130_fd_sc_hd__a21o_1 _16764_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09100_),
    .B1(_09777_),
    .X(_09778_));
 sky130_fd_sc_hd__xor2_1 _16765_ (.A(\rbzero.wall_tracer.mapX[10] ),
    .B(_09100_),
    .X(_09779_));
 sky130_fd_sc_hd__nand2_1 _16766_ (.A(_09778_),
    .B(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__o21a_1 _16767_ (.A1(_09778_),
    .A2(_09779_),
    .B1(_09762_),
    .X(_09781_));
 sky130_fd_sc_hd__a22o_1 _16768_ (.A1(\rbzero.wall_tracer.mapX[10] ),
    .A2(_09767_),
    .B1(_09780_),
    .B2(_09781_),
    .X(_00527_));
 sky130_fd_sc_hd__a21oi_4 _16769_ (.A1(_08130_),
    .A2(_06252_),
    .B1(_08111_),
    .Y(_09782_));
 sky130_fd_sc_hd__nor2_1 _16770_ (.A(_08924_),
    .B(_08974_),
    .Y(_09783_));
 sky130_fd_sc_hd__buf_6 _16771_ (.A(_08099_),
    .X(_09784_));
 sky130_fd_sc_hd__a211o_1 _16772_ (.A1(_08924_),
    .A2(_08974_),
    .B1(_09783_),
    .C1(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__o21ai_1 _16773_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09784_),
    .Y(_09786_));
 sky130_fd_sc_hd__a21o_1 _16774_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__and3_1 _16775_ (.A(_09782_),
    .B(_09785_),
    .C(_09787_),
    .X(_09788_));
 sky130_fd_sc_hd__a21oi_1 _16776_ (.A1(_06230_),
    .A2(_09767_),
    .B1(_09788_),
    .Y(_00528_));
 sky130_fd_sc_hd__clkbuf_8 _16777_ (.A(_06102_),
    .X(_09789_));
 sky130_fd_sc_hd__nand2_1 _16778_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_09790_));
 sky130_fd_sc_hd__or2_1 _16779_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_09791_));
 sky130_fd_sc_hd__and4_1 _16780_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .C(_09790_),
    .D(_09791_),
    .X(_09792_));
 sky130_fd_sc_hd__a22oi_1 _16781_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09790_),
    .B2(_09791_),
    .Y(_09793_));
 sky130_fd_sc_hd__clkbuf_4 _16782_ (.A(_09782_),
    .X(_09794_));
 sky130_fd_sc_hd__a21oi_1 _16783_ (.A1(_08976_),
    .A2(_08978_),
    .B1(_08100_),
    .Y(_09795_));
 sky130_fd_sc_hd__o21ai_1 _16784_ (.A1(_08976_),
    .A2(_08978_),
    .B1(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__o311a_1 _16785_ (.A1(_09789_),
    .A2(_09792_),
    .A3(_09793_),
    .B1(_09794_),
    .C1(_09796_),
    .X(_09797_));
 sky130_fd_sc_hd__a21oi_1 _16786_ (.A1(_06229_),
    .A2(_09767_),
    .B1(_09797_),
    .Y(_00529_));
 sky130_fd_sc_hd__a21o_1 _16787_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(\rbzero.wall_tracer.stepDistX[-10] ),
    .B1(_09792_),
    .X(_09798_));
 sky130_fd_sc_hd__or2_1 _16788_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_09799_));
 sky130_fd_sc_hd__nand2_1 _16789_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .Y(_09800_));
 sky130_fd_sc_hd__and3_1 _16790_ (.A(_09798_),
    .B(_09799_),
    .C(_09800_),
    .X(_09801_));
 sky130_fd_sc_hd__a21oi_1 _16791_ (.A1(_09799_),
    .A2(_09800_),
    .B1(_09798_),
    .Y(_09802_));
 sky130_fd_sc_hd__nand2_1 _16792_ (.A(_09760_),
    .B(_09090_),
    .Y(_09803_));
 sky130_fd_sc_hd__o311a_1 _16793_ (.A1(_09789_),
    .A2(_09801_),
    .A3(_09802_),
    .B1(_09794_),
    .C1(_09803_),
    .X(_09804_));
 sky130_fd_sc_hd__a21oi_1 _16794_ (.A1(_06228_),
    .A2(_09767_),
    .B1(_09804_),
    .Y(_00530_));
 sky130_fd_sc_hd__clkbuf_4 _16795_ (.A(_09782_),
    .X(_09805_));
 sky130_fd_sc_hd__or2_1 _16796_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_09806_));
 sky130_fd_sc_hd__nand2_1 _16797_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_09807_));
 sky130_fd_sc_hd__a21bo_1 _16798_ (.A1(_09798_),
    .A2(_09799_),
    .B1_N(_09800_),
    .X(_09808_));
 sky130_fd_sc_hd__nand3_1 _16799_ (.A(_09806_),
    .B(_09807_),
    .C(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__a21o_1 _16800_ (.A1(_09806_),
    .A2(_09807_),
    .B1(_09808_),
    .X(_09810_));
 sky130_fd_sc_hd__nor2_1 _16801_ (.A(_08100_),
    .B(_09093_),
    .Y(_09811_));
 sky130_fd_sc_hd__a311o_1 _16802_ (.A1(_08101_),
    .A2(_09809_),
    .A3(_09810_),
    .B1(_09761_),
    .C1(_09811_),
    .X(_09812_));
 sky130_fd_sc_hd__o21a_1 _16803_ (.A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .A2(_09805_),
    .B1(_09812_),
    .X(_00531_));
 sky130_fd_sc_hd__nor2_1 _16804_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09813_));
 sky130_fd_sc_hd__nand2_1 _16805_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09814_));
 sky130_fd_sc_hd__or2b_1 _16806_ (.A(_09813_),
    .B_N(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__a21boi_1 _16807_ (.A1(_09806_),
    .A2(_09808_),
    .B1_N(_09807_),
    .Y(_09816_));
 sky130_fd_sc_hd__xnor2_1 _16808_ (.A(_09815_),
    .B(_09816_),
    .Y(_09817_));
 sky130_fd_sc_hd__nand2_1 _16809_ (.A(_09760_),
    .B(_09086_),
    .Y(_09818_));
 sky130_fd_sc_hd__o211a_1 _16810_ (.A1(_09789_),
    .A2(_09817_),
    .B1(_09818_),
    .C1(_09794_),
    .X(_09819_));
 sky130_fd_sc_hd__a21oi_1 _16811_ (.A1(_06226_),
    .A2(_09767_),
    .B1(_09819_),
    .Y(_00532_));
 sky130_fd_sc_hd__or2_1 _16812_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_09820_));
 sky130_fd_sc_hd__nand2_1 _16813_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_09821_));
 sky130_fd_sc_hd__o21ai_1 _16814_ (.A1(_09813_),
    .A2(_09816_),
    .B1(_09814_),
    .Y(_09822_));
 sky130_fd_sc_hd__a21oi_1 _16815_ (.A1(_09820_),
    .A2(_09821_),
    .B1(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__buf_4 _16816_ (.A(_06101_),
    .X(_09824_));
 sky130_fd_sc_hd__a31o_1 _16817_ (.A1(_09820_),
    .A2(_09821_),
    .A3(_09822_),
    .B1(_09824_),
    .X(_09825_));
 sky130_fd_sc_hd__buf_6 _16818_ (.A(_09782_),
    .X(_09826_));
 sky130_fd_sc_hd__nand2_1 _16819_ (.A(_09760_),
    .B(_09082_),
    .Y(_09827_));
 sky130_fd_sc_hd__o211a_1 _16820_ (.A1(_09823_),
    .A2(_09825_),
    .B1(_09826_),
    .C1(_09827_),
    .X(_09828_));
 sky130_fd_sc_hd__a21oi_1 _16821_ (.A1(_06225_),
    .A2(_09767_),
    .B1(_09828_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_1 _16822_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09829_));
 sky130_fd_sc_hd__nand2_1 _16823_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09830_));
 sky130_fd_sc_hd__or2b_1 _16824_ (.A(_09829_),
    .B_N(_09830_),
    .X(_09831_));
 sky130_fd_sc_hd__a21boi_1 _16825_ (.A1(_09820_),
    .A2(_09822_),
    .B1_N(_09821_),
    .Y(_09832_));
 sky130_fd_sc_hd__xnor2_1 _16826_ (.A(_09831_),
    .B(_09832_),
    .Y(_09833_));
 sky130_fd_sc_hd__xor2_2 _16827_ (.A(_09105_),
    .B(_09211_),
    .X(_09834_));
 sky130_fd_sc_hd__nand2_1 _16828_ (.A(_09824_),
    .B(_09834_),
    .Y(_09835_));
 sky130_fd_sc_hd__o211a_1 _16829_ (.A1(_09789_),
    .A2(_09833_),
    .B1(_09835_),
    .C1(_09794_),
    .X(_09836_));
 sky130_fd_sc_hd__a21oi_1 _16830_ (.A1(_06224_),
    .A2(_09767_),
    .B1(_09836_),
    .Y(_00534_));
 sky130_fd_sc_hd__or2_1 _16831_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(_09837_));
 sky130_fd_sc_hd__nand2_1 _16832_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09838_));
 sky130_fd_sc_hd__o21ai_1 _16833_ (.A1(_09829_),
    .A2(_09832_),
    .B1(_09830_),
    .Y(_09839_));
 sky130_fd_sc_hd__a21oi_1 _16834_ (.A1(_09837_),
    .A2(_09838_),
    .B1(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__a31o_1 _16835_ (.A1(_09837_),
    .A2(_09838_),
    .A3(_09839_),
    .B1(_09824_),
    .X(_09841_));
 sky130_fd_sc_hd__or2_1 _16836_ (.A(_08100_),
    .B(_09324_),
    .X(_09842_));
 sky130_fd_sc_hd__o211a_1 _16837_ (.A1(_09840_),
    .A2(_09841_),
    .B1(_09826_),
    .C1(_09842_),
    .X(_09843_));
 sky130_fd_sc_hd__a21oi_1 _16838_ (.A1(_06223_),
    .A2(_09767_),
    .B1(_09843_),
    .Y(_00535_));
 sky130_fd_sc_hd__nor2_1 _16839_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09844_));
 sky130_fd_sc_hd__nand2_1 _16840_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09845_));
 sky130_fd_sc_hd__or2b_1 _16841_ (.A(_09844_),
    .B_N(_09845_),
    .X(_09846_));
 sky130_fd_sc_hd__a21boi_1 _16842_ (.A1(_09837_),
    .A2(_09839_),
    .B1_N(_09838_),
    .Y(_09847_));
 sky130_fd_sc_hd__xnor2_1 _16843_ (.A(_09846_),
    .B(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__or2_1 _16844_ (.A(_09784_),
    .B(_09446_),
    .X(_09849_));
 sky130_fd_sc_hd__o211a_1 _16845_ (.A1(_09789_),
    .A2(_09848_),
    .B1(_09849_),
    .C1(_09794_),
    .X(_09850_));
 sky130_fd_sc_hd__a21oi_1 _16846_ (.A1(_06222_),
    .A2(_09763_),
    .B1(_09850_),
    .Y(_00536_));
 sky130_fd_sc_hd__or2_1 _16847_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_09851_));
 sky130_fd_sc_hd__nand2_1 _16848_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_09852_));
 sky130_fd_sc_hd__o21ai_1 _16849_ (.A1(_09844_),
    .A2(_09847_),
    .B1(_09845_),
    .Y(_09853_));
 sky130_fd_sc_hd__a21oi_1 _16850_ (.A1(_09851_),
    .A2(_09852_),
    .B1(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__a31o_1 _16851_ (.A1(_09851_),
    .A2(_09852_),
    .A3(_09853_),
    .B1(_09824_),
    .X(_09855_));
 sky130_fd_sc_hd__nand2_1 _16852_ (.A(_09760_),
    .B(_09570_),
    .Y(_09856_));
 sky130_fd_sc_hd__o211a_1 _16853_ (.A1(_09854_),
    .A2(_09855_),
    .B1(_09826_),
    .C1(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__a21oi_1 _16854_ (.A1(_06220_),
    .A2(_09763_),
    .B1(_09857_),
    .Y(_00537_));
 sky130_fd_sc_hd__nor2_1 _16855_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_09858_));
 sky130_fd_sc_hd__and2_1 _16856_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(_09859_));
 sky130_fd_sc_hd__a21boi_1 _16857_ (.A1(_09851_),
    .A2(_09853_),
    .B1_N(_09852_),
    .Y(_09860_));
 sky130_fd_sc_hd__o21a_1 _16858_ (.A1(_09858_),
    .A2(_09859_),
    .B1(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__nor3_1 _16859_ (.A(_09858_),
    .B(_09859_),
    .C(_09860_),
    .Y(_09862_));
 sky130_fd_sc_hd__or2_1 _16860_ (.A(_09784_),
    .B(_09702_),
    .X(_09863_));
 sky130_fd_sc_hd__o311a_1 _16861_ (.A1(_09789_),
    .A2(_09861_),
    .A3(_09862_),
    .B1(_09794_),
    .C1(_09863_),
    .X(_09864_));
 sky130_fd_sc_hd__a21oi_1 _16862_ (.A1(_06216_),
    .A2(_09763_),
    .B1(_09864_),
    .Y(_00538_));
 sky130_fd_sc_hd__or2_1 _16863_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .X(_09865_));
 sky130_fd_sc_hd__nand2_1 _16864_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_09866_));
 sky130_fd_sc_hd__a211oi_1 _16865_ (.A1(_09865_),
    .A2(_09866_),
    .B1(_09859_),
    .C1(_09862_),
    .Y(_09867_));
 sky130_fd_sc_hd__o211a_1 _16866_ (.A1(_09859_),
    .A2(_09862_),
    .B1(_09865_),
    .C1(_09866_),
    .X(_09868_));
 sky130_fd_sc_hd__buf_4 _16867_ (.A(_09669_),
    .X(_09869_));
 sky130_fd_sc_hd__a31o_1 _16868_ (.A1(_08598_),
    .A2(_09588_),
    .A3(_09869_),
    .B1(_09586_),
    .X(_09870_));
 sky130_fd_sc_hd__or2b_1 _16869_ (.A(_09626_),
    .B_N(_09592_),
    .X(_09871_));
 sky130_fd_sc_hd__o2bb2a_1 _16870_ (.A1_N(_09604_),
    .A2_N(_09606_),
    .B1(_09600_),
    .B2(_09603_),
    .X(_09872_));
 sky130_fd_sc_hd__a21oi_1 _16871_ (.A1(_09624_),
    .A2(_09871_),
    .B1(_09872_),
    .Y(_09873_));
 sky130_fd_sc_hd__and3_1 _16872_ (.A(_09624_),
    .B(_09871_),
    .C(_09872_),
    .X(_09874_));
 sky130_fd_sc_hd__nor2_1 _16873_ (.A(_09873_),
    .B(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__a21o_1 _16874_ (.A1(_09607_),
    .A2(_09622_),
    .B1(_09620_),
    .X(_09876_));
 sky130_fd_sc_hd__or2b_1 _16875_ (.A(_09644_),
    .B_N(_09630_),
    .X(_09877_));
 sky130_fd_sc_hd__or2b_1 _16876_ (.A(_09645_),
    .B_N(_09628_),
    .X(_09878_));
 sky130_fd_sc_hd__nor2_1 _16877_ (.A(_09128_),
    .B(_09226_),
    .Y(_09879_));
 sky130_fd_sc_hd__nor2_1 _16878_ (.A(_08935_),
    .B(_09341_),
    .Y(_09880_));
 sky130_fd_sc_hd__xnor2_1 _16879_ (.A(_09879_),
    .B(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__nor2_1 _16880_ (.A(_08602_),
    .B(_09468_),
    .Y(_09882_));
 sky130_fd_sc_hd__xor2_1 _16881_ (.A(_09881_),
    .B(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__o31a_1 _16882_ (.A1(_09128_),
    .A2(_09227_),
    .A3(_09474_),
    .B1(_09598_),
    .X(_09884_));
 sky130_fd_sc_hd__nor2_1 _16883_ (.A(_09883_),
    .B(_09884_),
    .Y(_09885_));
 sky130_fd_sc_hd__nand2_1 _16884_ (.A(_09883_),
    .B(_09884_),
    .Y(_09886_));
 sky130_fd_sc_hd__and2b_1 _16885_ (.A_N(_09885_),
    .B(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__or2_1 _16886_ (.A(_08145_),
    .B(_09589_),
    .X(_09888_));
 sky130_fd_sc_hd__xnor2_1 _16887_ (.A(_09887_),
    .B(_09888_),
    .Y(_09889_));
 sky130_fd_sc_hd__o21ai_1 _16888_ (.A1(_09476_),
    .A2(_09610_),
    .B1(_09612_),
    .Y(_09890_));
 sky130_fd_sc_hd__o21ai_1 _16889_ (.A1(_09631_),
    .A2(_09634_),
    .B1(_09632_),
    .Y(_09891_));
 sky130_fd_sc_hd__o21a_1 _16890_ (.A1(_09252_),
    .A2(_09056_),
    .B1(_09611_),
    .X(_09892_));
 sky130_fd_sc_hd__or3_1 _16891_ (.A(_09252_),
    .B(_09056_),
    .C(_09611_),
    .X(_09893_));
 sky130_fd_sc_hd__or2b_1 _16892_ (.A(_09892_),
    .B_N(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__nor2_1 _16893_ (.A(_09127_),
    .B(_09111_),
    .Y(_09895_));
 sky130_fd_sc_hd__xnor2_1 _16894_ (.A(_09894_),
    .B(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__xor2_1 _16895_ (.A(_09891_),
    .B(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__xnor2_1 _16896_ (.A(_09890_),
    .B(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__a21oi_1 _16897_ (.A1(_09608_),
    .A2(_09616_),
    .B1(_09615_),
    .Y(_09899_));
 sky130_fd_sc_hd__nor2_1 _16898_ (.A(_09898_),
    .B(_09899_),
    .Y(_09900_));
 sky130_fd_sc_hd__and2_1 _16899_ (.A(_09898_),
    .B(_09899_),
    .X(_09901_));
 sky130_fd_sc_hd__nor2_1 _16900_ (.A(_09900_),
    .B(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__xnor2_1 _16901_ (.A(_09889_),
    .B(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__a21o_1 _16902_ (.A1(_09877_),
    .A2(_09878_),
    .B1(_09903_),
    .X(_09904_));
 sky130_fd_sc_hd__nand3_1 _16903_ (.A(_09877_),
    .B(_09878_),
    .C(_09903_),
    .Y(_09905_));
 sky130_fd_sc_hd__nand2_1 _16904_ (.A(_09904_),
    .B(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__xnor2_1 _16905_ (.A(_09876_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__a21o_1 _16906_ (.A1(_09635_),
    .A2(_09642_),
    .B1(_09641_),
    .X(_09908_));
 sky130_fd_sc_hd__a21o_1 _16907_ (.A1(_09649_),
    .A2(_09658_),
    .B1(_09656_),
    .X(_09909_));
 sky130_fd_sc_hd__o21a_2 _16908_ (.A1(_08319_),
    .A2(_08374_),
    .B1(_08375_),
    .X(_09910_));
 sky130_fd_sc_hd__clkbuf_4 _16909_ (.A(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__o22a_1 _16910_ (.A1(_08127_),
    .A2(_09911_),
    .B1(_08385_),
    .B2(_08286_),
    .X(_09912_));
 sky130_fd_sc_hd__or4_1 _16911_ (.A(_08126_),
    .B(_08286_),
    .C(_09910_),
    .D(_08385_),
    .X(_09913_));
 sky130_fd_sc_hd__or2b_1 _16912_ (.A(_09912_),
    .B_N(_09913_),
    .X(_09914_));
 sky130_fd_sc_hd__buf_2 _16913_ (.A(_08649_),
    .X(_09915_));
 sky130_fd_sc_hd__nor2_1 _16914_ (.A(_09915_),
    .B(_09132_),
    .Y(_09916_));
 sky130_fd_sc_hd__xnor2_1 _16915_ (.A(_09914_),
    .B(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__nor2_1 _16916_ (.A(_08325_),
    .B(_08409_),
    .Y(_09918_));
 sky130_fd_sc_hd__xnor2_1 _16917_ (.A(_09636_),
    .B(_09918_),
    .Y(_09919_));
 sky130_fd_sc_hd__or2_1 _16918_ (.A(_08546_),
    .B(_08411_),
    .X(_09920_));
 sky130_fd_sc_hd__xnor2_1 _16919_ (.A(_09919_),
    .B(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__a22oi_1 _16920_ (.A1(_09527_),
    .A2(_09636_),
    .B1(_09637_),
    .B2(_09507_),
    .Y(_09922_));
 sky130_fd_sc_hd__nor2_1 _16921_ (.A(_09921_),
    .B(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_1 _16922_ (.A(_09921_),
    .B(_09922_),
    .Y(_09924_));
 sky130_fd_sc_hd__and2b_1 _16923_ (.A_N(_09923_),
    .B(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__xnor2_1 _16924_ (.A(_09917_),
    .B(_09925_),
    .Y(_09926_));
 sky130_fd_sc_hd__xor2_1 _16925_ (.A(_09909_),
    .B(_09926_),
    .X(_09927_));
 sky130_fd_sc_hd__xnor2_1 _16926_ (.A(_09908_),
    .B(_09927_),
    .Y(_09928_));
 sky130_fd_sc_hd__a21oi_1 _16927_ (.A1(_09180_),
    .A2(_09287_),
    .B1(_08352_),
    .Y(_09929_));
 sky130_fd_sc_hd__a22o_1 _16928_ (.A1(_09537_),
    .A2(_09929_),
    .B1(_09654_),
    .B2(_09651_),
    .X(_09930_));
 sky130_fd_sc_hd__o21bai_1 _16929_ (.A1(_09660_),
    .A2(_09665_),
    .B1_N(_09664_),
    .Y(_09931_));
 sky130_fd_sc_hd__a21oi_1 _16930_ (.A1(_08448_),
    .A2(_09168_),
    .B1(_08243_),
    .Y(_09932_));
 sky130_fd_sc_hd__xnor2_1 _16931_ (.A(_09929_),
    .B(_09932_),
    .Y(_09933_));
 sky130_fd_sc_hd__a21o_1 _16932_ (.A1(_08454_),
    .A2(_09025_),
    .B1(_08267_),
    .X(_09934_));
 sky130_fd_sc_hd__xor2_1 _16933_ (.A(_09933_),
    .B(_09934_),
    .X(_09935_));
 sky130_fd_sc_hd__and2_1 _16934_ (.A(_09931_),
    .B(_09935_),
    .X(_09936_));
 sky130_fd_sc_hd__or2_1 _16935_ (.A(_09931_),
    .B(_09935_),
    .X(_09937_));
 sky130_fd_sc_hd__or2b_1 _16936_ (.A(_09936_),
    .B_N(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__xnor2_2 _16937_ (.A(_09930_),
    .B(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__or2_1 _16938_ (.A(_08359_),
    .B(_09534_),
    .X(_09940_));
 sky130_fd_sc_hd__nor2_1 _16939_ (.A(_08911_),
    .B(_09540_),
    .Y(_09941_));
 sky130_fd_sc_hd__nor2_1 _16940_ (.A(_08941_),
    .B(_09663_),
    .Y(_09942_));
 sky130_fd_sc_hd__o22a_1 _16941_ (.A1(_08399_),
    .A2(_09540_),
    .B1(_09663_),
    .B2(_08911_),
    .X(_09943_));
 sky130_fd_sc_hd__a21o_1 _16942_ (.A1(_09941_),
    .A2(_09942_),
    .B1(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__xor2_1 _16943_ (.A(_09940_),
    .B(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__a2bb2o_1 _16944_ (.A1_N(_06135_),
    .A2_N(_09672_),
    .B1(_09673_),
    .B2(_09675_),
    .X(_09946_));
 sky130_fd_sc_hd__nand2_2 _16945_ (.A(\rbzero.wall_tracer.stepDistX[10] ),
    .B(_06162_),
    .Y(_09947_));
 sky130_fd_sc_hd__nand2_1 _16946_ (.A(\rbzero.wall_tracer.stepDistY[10] ),
    .B(_08135_),
    .Y(_09948_));
 sky130_fd_sc_hd__a21o_1 _16947_ (.A1(_09671_),
    .A2(_09948_),
    .B1(_06162_),
    .X(_09949_));
 sky130_fd_sc_hd__a21o_2 _16948_ (.A1(_09947_),
    .A2(_09949_),
    .B1(_08420_),
    .X(_09950_));
 sky130_fd_sc_hd__a21o_1 _16949_ (.A1(_09674_),
    .A2(_09545_),
    .B1(_06163_),
    .X(_09951_));
 sky130_fd_sc_hd__nand2_2 _16950_ (.A(\rbzero.wall_tracer.stepDistX[9] ),
    .B(_06163_),
    .Y(_09952_));
 sky130_fd_sc_hd__a21oi_1 _16951_ (.A1(_09951_),
    .A2(_09952_),
    .B1(_08928_),
    .Y(_09953_));
 sky130_fd_sc_hd__nor2_1 _16952_ (.A(_08018_),
    .B(_08406_),
    .Y(_09954_));
 sky130_fd_sc_hd__or3_1 _16953_ (.A(_08018_),
    .B(_08319_),
    .C(_09671_),
    .X(_09955_));
 sky130_fd_sc_hd__mux2_1 _16954_ (.A0(_09954_),
    .A1(_09955_),
    .S(_09672_),
    .X(_09956_));
 sky130_fd_sc_hd__mux2_1 _16955_ (.A0(_09950_),
    .A1(_09953_),
    .S(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__xor2_1 _16956_ (.A(_09946_),
    .B(_09957_),
    .X(_09958_));
 sky130_fd_sc_hd__xnor2_1 _16957_ (.A(_09945_),
    .B(_09958_),
    .Y(_09959_));
 sky130_fd_sc_hd__or2b_1 _16958_ (.A(_09676_),
    .B_N(_09678_),
    .X(_09960_));
 sky130_fd_sc_hd__a21bo_1 _16959_ (.A1(_09668_),
    .A2(_09679_),
    .B1_N(_09960_),
    .X(_09961_));
 sky130_fd_sc_hd__xnor2_1 _16960_ (.A(_09959_),
    .B(_09961_),
    .Y(_09962_));
 sky130_fd_sc_hd__xnor2_2 _16961_ (.A(_09939_),
    .B(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__or2b_1 _16962_ (.A(_09680_),
    .B_N(_09682_),
    .X(_09964_));
 sky130_fd_sc_hd__a21bo_1 _16963_ (.A1(_09659_),
    .A2(_09683_),
    .B1_N(_09964_),
    .X(_09965_));
 sky130_fd_sc_hd__xnor2_1 _16964_ (.A(_09963_),
    .B(_09965_),
    .Y(_09966_));
 sky130_fd_sc_hd__xnor2_1 _16965_ (.A(_09928_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__and2b_1 _16966_ (.A_N(_09684_),
    .B(_09686_),
    .X(_09968_));
 sky130_fd_sc_hd__a21oi_1 _16967_ (.A1(_09646_),
    .A2(_09687_),
    .B1(_09968_),
    .Y(_09969_));
 sky130_fd_sc_hd__or2_1 _16968_ (.A(_09967_),
    .B(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__nand2_1 _16969_ (.A(_09967_),
    .B(_09969_),
    .Y(_09971_));
 sky130_fd_sc_hd__and2_1 _16970_ (.A(_09970_),
    .B(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__xnor2_1 _16971_ (.A(_09907_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__a21oi_1 _16972_ (.A1(_09627_),
    .A2(_09693_),
    .B1(_09691_),
    .Y(_09974_));
 sky130_fd_sc_hd__xor2_1 _16973_ (.A(_09973_),
    .B(_09974_),
    .X(_09975_));
 sky130_fd_sc_hd__nand2_1 _16974_ (.A(_09875_),
    .B(_09975_),
    .Y(_09976_));
 sky130_fd_sc_hd__or2_1 _16975_ (.A(_09875_),
    .B(_09975_),
    .X(_09977_));
 sky130_fd_sc_hd__nand2_1 _16976_ (.A(_09976_),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__o2bb2a_1 _16977_ (.A1_N(_09591_),
    .A2_N(_09696_),
    .B1(_09695_),
    .B2(_09694_),
    .X(_09979_));
 sky130_fd_sc_hd__xor2_1 _16978_ (.A(_09978_),
    .B(_09979_),
    .X(_09980_));
 sky130_fd_sc_hd__nand2_1 _16979_ (.A(_09870_),
    .B(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__or2_1 _16980_ (.A(_09870_),
    .B(_09980_),
    .X(_09982_));
 sky130_fd_sc_hd__and2_1 _16981_ (.A(_09981_),
    .B(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__nand2_1 _16982_ (.A(_09698_),
    .B(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__or2_1 _16983_ (.A(_09698_),
    .B(_09983_),
    .X(_09985_));
 sky130_fd_sc_hd__nand2_2 _16984_ (.A(_09984_),
    .B(_09985_),
    .Y(_09986_));
 sky130_fd_sc_hd__a21oi_1 _16985_ (.A1(_09582_),
    .A2(_09580_),
    .B1(_09700_),
    .Y(_09987_));
 sky130_fd_sc_hd__a31oi_4 _16986_ (.A1(_09457_),
    .A2(_09579_),
    .A3(_09701_),
    .B1(_09987_),
    .Y(_09988_));
 sky130_fd_sc_hd__xor2_4 _16987_ (.A(_09986_),
    .B(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__nand2_1 _16988_ (.A(_09760_),
    .B(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__o311a_1 _16989_ (.A1(_09789_),
    .A2(_09867_),
    .A3(_09868_),
    .B1(_09794_),
    .C1(_09990_),
    .X(_09991_));
 sky130_fd_sc_hd__a21oi_1 _16990_ (.A1(_06219_),
    .A2(_09763_),
    .B1(_09991_),
    .Y(_00539_));
 sky130_fd_sc_hd__or2_1 _16991_ (.A(_09978_),
    .B(_09979_),
    .X(_09992_));
 sky130_fd_sc_hd__or2b_1 _16992_ (.A(_09906_),
    .B_N(_09876_),
    .X(_09993_));
 sky130_fd_sc_hd__a31oi_1 _16993_ (.A1(_08285_),
    .A2(_09869_),
    .A3(_09886_),
    .B1(_09885_),
    .Y(_09994_));
 sky130_fd_sc_hd__a21oi_1 _16994_ (.A1(_09904_),
    .A2(_09993_),
    .B1(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__and3_1 _16995_ (.A(_09904_),
    .B(_09993_),
    .C(_09994_),
    .X(_09996_));
 sky130_fd_sc_hd__nor2_1 _16996_ (.A(_09995_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(_09907_),
    .B(_09972_),
    .Y(_09998_));
 sky130_fd_sc_hd__a21o_1 _16998_ (.A1(_09889_),
    .A2(_09902_),
    .B1(_09900_),
    .X(_09999_));
 sky130_fd_sc_hd__or2b_1 _16999_ (.A(_09926_),
    .B_N(_09909_),
    .X(_10000_));
 sky130_fd_sc_hd__or2b_1 _17000_ (.A(_09927_),
    .B_N(_09908_),
    .X(_10001_));
 sky130_fd_sc_hd__nand2_1 _17001_ (.A(_10000_),
    .B(_10001_),
    .Y(_10002_));
 sky130_fd_sc_hd__or2_1 _17002_ (.A(_09127_),
    .B(_09341_),
    .X(_10003_));
 sky130_fd_sc_hd__or2_1 _17003_ (.A(_09128_),
    .B(_09341_),
    .X(_10004_));
 sky130_fd_sc_hd__o21ai_1 _17004_ (.A1(_09127_),
    .A2(_09227_),
    .B1(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__o31a_1 _17005_ (.A1(_09128_),
    .A2(_09227_),
    .A3(_10003_),
    .B1(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__nor2_1 _17006_ (.A(_08935_),
    .B(_09469_),
    .Y(_10007_));
 sky130_fd_sc_hd__nand2_1 _17007_ (.A(_10006_),
    .B(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__or2_1 _17008_ (.A(_10006_),
    .B(_10007_),
    .X(_10009_));
 sky130_fd_sc_hd__nand2_1 _17009_ (.A(_10008_),
    .B(_10009_),
    .Y(_10010_));
 sky130_fd_sc_hd__nand2_1 _17010_ (.A(_09879_),
    .B(_09880_),
    .Y(_10011_));
 sky130_fd_sc_hd__o31a_1 _17011_ (.A1(_08602_),
    .A2(_09469_),
    .A3(_09881_),
    .B1(_10011_),
    .X(_10012_));
 sky130_fd_sc_hd__xor2_1 _17012_ (.A(_10010_),
    .B(_10012_),
    .X(_10013_));
 sky130_fd_sc_hd__and2_1 _17013_ (.A(_08602_),
    .B(_09869_),
    .X(_10014_));
 sky130_fd_sc_hd__xor2_1 _17014_ (.A(_10013_),
    .B(_10014_),
    .X(_10015_));
 sky130_fd_sc_hd__o31ai_2 _17015_ (.A1(_09127_),
    .A2(_09111_),
    .A3(_09892_),
    .B1(_09893_),
    .Y(_10016_));
 sky130_fd_sc_hd__nor2_1 _17016_ (.A(_09369_),
    .B(_09055_),
    .Y(_10017_));
 sky130_fd_sc_hd__nor2_1 _17017_ (.A(_08649_),
    .B(_08599_),
    .Y(_10018_));
 sky130_fd_sc_hd__xnor2_1 _17018_ (.A(_10017_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__or3_1 _17019_ (.A(_09503_),
    .B(_09110_),
    .C(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__o21ai_1 _17020_ (.A1(_09503_),
    .A2(_09111_),
    .B1(_10019_),
    .Y(_10021_));
 sky130_fd_sc_hd__nand2_1 _17021_ (.A(_10020_),
    .B(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__o31ai_1 _17022_ (.A1(_09915_),
    .A2(_09132_),
    .A3(_09912_),
    .B1(_09913_),
    .Y(_10023_));
 sky130_fd_sc_hd__and2b_1 _17023_ (.A_N(_10022_),
    .B(_10023_),
    .X(_10024_));
 sky130_fd_sc_hd__and2b_1 _17024_ (.A_N(_10023_),
    .B(_10022_),
    .X(_10025_));
 sky130_fd_sc_hd__nor2_1 _17025_ (.A(_10024_),
    .B(_10025_),
    .Y(_10026_));
 sky130_fd_sc_hd__xnor2_1 _17026_ (.A(_10016_),
    .B(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__and2_1 _17027_ (.A(_09891_),
    .B(_09896_),
    .X(_10028_));
 sky130_fd_sc_hd__a21oi_1 _17028_ (.A1(_09890_),
    .A2(_09897_),
    .B1(_10028_),
    .Y(_10029_));
 sky130_fd_sc_hd__nor2_1 _17029_ (.A(_10027_),
    .B(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__and2_1 _17030_ (.A(_10027_),
    .B(_10029_),
    .X(_10031_));
 sky130_fd_sc_hd__nor2_1 _17031_ (.A(_10030_),
    .B(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__xor2_1 _17032_ (.A(_10015_),
    .B(_10032_),
    .X(_10033_));
 sky130_fd_sc_hd__xnor2_1 _17033_ (.A(_10002_),
    .B(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__xnor2_1 _17034_ (.A(_09999_),
    .B(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__a21o_1 _17035_ (.A1(_09917_),
    .A2(_09924_),
    .B1(_09923_),
    .X(_10036_));
 sky130_fd_sc_hd__a21o_1 _17036_ (.A1(_09930_),
    .A2(_09937_),
    .B1(_09936_),
    .X(_10037_));
 sky130_fd_sc_hd__clkbuf_4 _17037_ (.A(_08385_),
    .X(_10038_));
 sky130_fd_sc_hd__nor2_1 _17038_ (.A(_08126_),
    .B(_09910_),
    .Y(_10039_));
 sky130_fd_sc_hd__nor2_1 _17039_ (.A(_08148_),
    .B(_08368_),
    .Y(_10040_));
 sky130_fd_sc_hd__o22a_1 _17040_ (.A1(_08126_),
    .A2(_08368_),
    .B1(_09910_),
    .B2(_08148_),
    .X(_10041_));
 sky130_fd_sc_hd__a21o_1 _17041_ (.A1(_10039_),
    .A2(_10040_),
    .B1(_10041_),
    .X(_10042_));
 sky130_fd_sc_hd__or3_1 _17042_ (.A(_10038_),
    .B(_08534_),
    .C(_10042_),
    .X(_10043_));
 sky130_fd_sc_hd__o21ai_1 _17043_ (.A1(_10038_),
    .A2(_09132_),
    .B1(_10042_),
    .Y(_10044_));
 sky130_fd_sc_hd__and2_1 _17044_ (.A(_10043_),
    .B(_10044_),
    .X(_10045_));
 sky130_fd_sc_hd__nor2_1 _17045_ (.A(_08325_),
    .B(_08427_),
    .Y(_10046_));
 sky130_fd_sc_hd__a21oi_1 _17046_ (.A1(_08454_),
    .A2(_09025_),
    .B1(_08797_),
    .Y(_10047_));
 sky130_fd_sc_hd__xnor2_1 _17047_ (.A(_10046_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__nor2_1 _17048_ (.A(_09140_),
    .B(_08409_),
    .Y(_10049_));
 sky130_fd_sc_hd__xor2_1 _17049_ (.A(_10048_),
    .B(_10049_),
    .X(_10050_));
 sky130_fd_sc_hd__o2bb2a_1 _17050_ (.A1_N(_09636_),
    .A2_N(_09918_),
    .B1(_09919_),
    .B2(_09920_),
    .X(_10051_));
 sky130_fd_sc_hd__nor2_1 _17051_ (.A(_10050_),
    .B(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__nand2_1 _17052_ (.A(_10050_),
    .B(_10051_),
    .Y(_10053_));
 sky130_fd_sc_hd__and2b_1 _17053_ (.A_N(_10052_),
    .B(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__xor2_1 _17054_ (.A(_10045_),
    .B(_10054_),
    .X(_10055_));
 sky130_fd_sc_hd__xnor2_1 _17055_ (.A(_10037_),
    .B(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__xnor2_1 _17056_ (.A(_10036_),
    .B(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__a21oi_2 _17057_ (.A1(_09286_),
    .A2(_09287_),
    .B1(_08876_),
    .Y(_10058_));
 sky130_fd_sc_hd__o2bb2ai_1 _17058_ (.A1_N(_09653_),
    .A2_N(_10058_),
    .B1(_09933_),
    .B2(_09934_),
    .Y(_10059_));
 sky130_fd_sc_hd__a2bb2o_1 _17059_ (.A1_N(_09940_),
    .A2_N(_09943_),
    .B1(_09942_),
    .B2(_09941_),
    .X(_10060_));
 sky130_fd_sc_hd__a21oi_2 _17060_ (.A1(_09181_),
    .A2(_09402_),
    .B1(_08875_),
    .Y(_10061_));
 sky130_fd_sc_hd__xnor2_1 _17061_ (.A(_10058_),
    .B(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__nor2_1 _17062_ (.A(_08394_),
    .B(_09170_),
    .Y(_10063_));
 sky130_fd_sc_hd__xnor2_1 _17063_ (.A(_10062_),
    .B(_10063_),
    .Y(_10064_));
 sky130_fd_sc_hd__nand2_1 _17064_ (.A(_10060_),
    .B(_10064_),
    .Y(_10065_));
 sky130_fd_sc_hd__or2_1 _17065_ (.A(_10060_),
    .B(_10064_),
    .X(_10066_));
 sky130_fd_sc_hd__nand2_1 _17066_ (.A(_10065_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__xnor2_1 _17067_ (.A(_10059_),
    .B(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__buf_2 _17068_ (.A(_09540_),
    .X(_10069_));
 sky130_fd_sc_hd__nor2_1 _17069_ (.A(_08360_),
    .B(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__a21oi_1 _17070_ (.A1(_09951_),
    .A2(_09952_),
    .B1(_08911_),
    .Y(_10071_));
 sky130_fd_sc_hd__xor2_1 _17071_ (.A(_09942_),
    .B(_10071_),
    .X(_10072_));
 sky130_fd_sc_hd__xor2_1 _17072_ (.A(_10070_),
    .B(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__and2_1 _17073_ (.A(_09672_),
    .B(_09955_),
    .X(_10074_));
 sky130_fd_sc_hd__nor3_4 _17074_ (.A(_08447_),
    .B(_09672_),
    .C(_09950_),
    .Y(_10075_));
 sky130_fd_sc_hd__a21oi_4 _17075_ (.A1(_10074_),
    .A2(_09950_),
    .B1(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__xnor2_1 _17076_ (.A(_10073_),
    .B(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__and2_1 _17077_ (.A(_09946_),
    .B(_09957_),
    .X(_10078_));
 sky130_fd_sc_hd__a21oi_1 _17078_ (.A1(_09945_),
    .A2(_09958_),
    .B1(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__xor2_1 _17079_ (.A(_10077_),
    .B(_10079_),
    .X(_10080_));
 sky130_fd_sc_hd__xnor2_1 _17080_ (.A(_10068_),
    .B(_10080_),
    .Y(_10081_));
 sky130_fd_sc_hd__or2b_1 _17081_ (.A(_09959_),
    .B_N(_09961_),
    .X(_10082_));
 sky130_fd_sc_hd__a21bo_1 _17082_ (.A1(_09939_),
    .A2(_09962_),
    .B1_N(_10082_),
    .X(_10083_));
 sky130_fd_sc_hd__xnor2_1 _17083_ (.A(_10081_),
    .B(_10083_),
    .Y(_10084_));
 sky130_fd_sc_hd__xnor2_1 _17084_ (.A(_10057_),
    .B(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__or2b_1 _17085_ (.A(_09963_),
    .B_N(_09965_),
    .X(_10086_));
 sky130_fd_sc_hd__a21boi_1 _17086_ (.A1(_09928_),
    .A2(_09966_),
    .B1_N(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__nor2_1 _17087_ (.A(_10085_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__and2_1 _17088_ (.A(_10085_),
    .B(_10087_),
    .X(_10089_));
 sky130_fd_sc_hd__nor2_1 _17089_ (.A(_10088_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__xnor2_1 _17090_ (.A(_10035_),
    .B(_10090_),
    .Y(_10091_));
 sky130_fd_sc_hd__a21oi_1 _17091_ (.A1(_09970_),
    .A2(_09998_),
    .B1(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__and3_1 _17092_ (.A(_09970_),
    .B(_09998_),
    .C(_10091_),
    .X(_10093_));
 sky130_fd_sc_hd__nor2_1 _17093_ (.A(_10092_),
    .B(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__xnor2_1 _17094_ (.A(_09997_),
    .B(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__o21a_1 _17095_ (.A1(_09973_),
    .A2(_09974_),
    .B1(_09976_),
    .X(_10096_));
 sky130_fd_sc_hd__nor2_1 _17096_ (.A(_10095_),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__and2_1 _17097_ (.A(_10095_),
    .B(_10096_),
    .X(_10098_));
 sky130_fd_sc_hd__nor2_1 _17098_ (.A(_10097_),
    .B(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__xnor2_1 _17099_ (.A(_09873_),
    .B(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__a21oi_1 _17100_ (.A1(_09992_),
    .A2(_09981_),
    .B1(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__and3_1 _17101_ (.A(_09992_),
    .B(_09981_),
    .C(_10100_),
    .X(_10102_));
 sky130_fd_sc_hd__or2_2 _17102_ (.A(_10101_),
    .B(_10102_),
    .X(_10103_));
 sky130_fd_sc_hd__o21ai_2 _17103_ (.A1(_09986_),
    .A2(_09988_),
    .B1(_09984_),
    .Y(_10104_));
 sky130_fd_sc_hd__xnor2_4 _17104_ (.A(_10103_),
    .B(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__nand2_1 _17105_ (.A(_09824_),
    .B(_10105_),
    .Y(_10106_));
 sky130_fd_sc_hd__buf_6 _17106_ (.A(_09824_),
    .X(_10107_));
 sky130_fd_sc_hd__nand2_1 _17107_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_10108_));
 sky130_fd_sc_hd__or2_1 _17108_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_10109_));
 sky130_fd_sc_hd__a21o_1 _17109_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(\rbzero.wall_tracer.stepDistX[0] ),
    .B1(_09868_),
    .X(_10110_));
 sky130_fd_sc_hd__and3_1 _17110_ (.A(_10108_),
    .B(_10109_),
    .C(_10110_),
    .X(_10111_));
 sky130_fd_sc_hd__a21oi_1 _17111_ (.A1(_10108_),
    .A2(_10109_),
    .B1(_10110_),
    .Y(_10112_));
 sky130_fd_sc_hd__o31a_1 _17112_ (.A1(_10107_),
    .A2(_10111_),
    .A3(_10112_),
    .B1(_09794_),
    .X(_10113_));
 sky130_fd_sc_hd__o2bb2a_1 _17113_ (.A1_N(_10106_),
    .A2_N(_10113_),
    .B1(\rbzero.wall_tracer.trackDistX[1] ),
    .B2(_09805_),
    .X(_00540_));
 sky130_fd_sc_hd__nand2_1 _17114_ (.A(_10002_),
    .B(_10033_),
    .Y(_10114_));
 sky130_fd_sc_hd__or2b_1 _17115_ (.A(_10034_),
    .B_N(_09999_),
    .X(_10115_));
 sky130_fd_sc_hd__o2bb2a_1 _17116_ (.A1_N(_10013_),
    .A2_N(_10014_),
    .B1(_10010_),
    .B2(_10012_),
    .X(_10116_));
 sky130_fd_sc_hd__a21oi_1 _17117_ (.A1(_10114_),
    .A2(_10115_),
    .B1(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__and3_1 _17118_ (.A(_10114_),
    .B(_10115_),
    .C(_10116_),
    .X(_10118_));
 sky130_fd_sc_hd__nor2_1 _17119_ (.A(_10117_),
    .B(_10118_),
    .Y(_10119_));
 sky130_fd_sc_hd__a21o_1 _17120_ (.A1(_10015_),
    .A2(_10032_),
    .B1(_10030_),
    .X(_10120_));
 sky130_fd_sc_hd__or2b_1 _17121_ (.A(_10056_),
    .B_N(_10036_),
    .X(_10121_));
 sky130_fd_sc_hd__a21bo_1 _17122_ (.A1(_10037_),
    .A2(_10055_),
    .B1_N(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__o21ai_1 _17123_ (.A1(_09503_),
    .A2(_09227_),
    .B1(_10003_),
    .Y(_10123_));
 sky130_fd_sc_hd__or3_1 _17124_ (.A(_09503_),
    .B(_09227_),
    .C(_10003_),
    .X(_10124_));
 sky130_fd_sc_hd__nand2_1 _17125_ (.A(_10123_),
    .B(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__nor2_1 _17126_ (.A(_09128_),
    .B(_09469_),
    .Y(_10126_));
 sky130_fd_sc_hd__xor2_1 _17127_ (.A(_10125_),
    .B(_10126_),
    .X(_10127_));
 sky130_fd_sc_hd__o31a_1 _17128_ (.A1(_09127_),
    .A2(_09228_),
    .A3(_10004_),
    .B1(_10008_),
    .X(_10128_));
 sky130_fd_sc_hd__xor2_1 _17129_ (.A(_10127_),
    .B(_10128_),
    .X(_10129_));
 sky130_fd_sc_hd__and2_1 _17130_ (.A(_08935_),
    .B(_09869_),
    .X(_10130_));
 sky130_fd_sc_hd__xor2_1 _17131_ (.A(_10129_),
    .B(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__a21bo_1 _17132_ (.A1(_10017_),
    .A2(_10018_),
    .B1_N(_10020_),
    .X(_10132_));
 sky130_fd_sc_hd__o22ai_1 _17133_ (.A1(_10038_),
    .A2(_08600_),
    .B1(_09056_),
    .B2(_09915_),
    .Y(_10133_));
 sky130_fd_sc_hd__or4_1 _17134_ (.A(_08649_),
    .B(_08385_),
    .C(_08600_),
    .D(_09056_),
    .X(_10134_));
 sky130_fd_sc_hd__nand2_1 _17135_ (.A(_10133_),
    .B(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__nor2_1 _17136_ (.A(_09369_),
    .B(_09111_),
    .Y(_10136_));
 sky130_fd_sc_hd__xor2_1 _17137_ (.A(_10135_),
    .B(_10136_),
    .X(_10137_));
 sky130_fd_sc_hd__a21bo_1 _17138_ (.A1(_10039_),
    .A2(_10040_),
    .B1_N(_10043_),
    .X(_10138_));
 sky130_fd_sc_hd__and2b_1 _17139_ (.A_N(_10137_),
    .B(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__and2b_1 _17140_ (.A_N(_10138_),
    .B(_10137_),
    .X(_10140_));
 sky130_fd_sc_hd__nor2_1 _17141_ (.A(_10139_),
    .B(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__xnor2_1 _17142_ (.A(_10132_),
    .B(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__a21oi_1 _17143_ (.A1(_10016_),
    .A2(_10026_),
    .B1(_10024_),
    .Y(_10143_));
 sky130_fd_sc_hd__nor2_1 _17144_ (.A(_10142_),
    .B(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__and2_1 _17145_ (.A(_10142_),
    .B(_10143_),
    .X(_10145_));
 sky130_fd_sc_hd__nor2_1 _17146_ (.A(_10144_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__xor2_1 _17147_ (.A(_10131_),
    .B(_10146_),
    .X(_10147_));
 sky130_fd_sc_hd__xnor2_1 _17148_ (.A(_10122_),
    .B(_10147_),
    .Y(_10148_));
 sky130_fd_sc_hd__xnor2_1 _17149_ (.A(_10120_),
    .B(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__a21o_1 _17150_ (.A1(_10045_),
    .A2(_10053_),
    .B1(_10052_),
    .X(_10150_));
 sky130_fd_sc_hd__a21bo_1 _17151_ (.A1(_10059_),
    .A2(_10066_),
    .B1_N(_10065_),
    .X(_10151_));
 sky130_fd_sc_hd__nor2_1 _17152_ (.A(_08126_),
    .B(_08479_),
    .Y(_10152_));
 sky130_fd_sc_hd__xnor2_1 _17153_ (.A(_10040_),
    .B(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__or3_1 _17154_ (.A(_09911_),
    .B(_09132_),
    .C(_10153_),
    .X(_10154_));
 sky130_fd_sc_hd__o21ai_1 _17155_ (.A1(_09911_),
    .A2(_09132_),
    .B1(_10153_),
    .Y(_10155_));
 sky130_fd_sc_hd__and2_1 _17156_ (.A(_10154_),
    .B(_10155_),
    .X(_10156_));
 sky130_fd_sc_hd__a21oi_2 _17157_ (.A1(_08454_),
    .A2(_09025_),
    .B1(_08325_),
    .Y(_10157_));
 sky130_fd_sc_hd__a21oi_2 _17158_ (.A1(_09295_),
    .A2(_09168_),
    .B1(_08797_),
    .Y(_10158_));
 sky130_fd_sc_hd__xnor2_1 _17159_ (.A(_10157_),
    .B(_10158_),
    .Y(_10159_));
 sky130_fd_sc_hd__or2_1 _17160_ (.A(_09140_),
    .B(_08427_),
    .X(_10160_));
 sky130_fd_sc_hd__xnor2_1 _17161_ (.A(_10159_),
    .B(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__nand2_1 _17162_ (.A(_09636_),
    .B(_10157_),
    .Y(_10162_));
 sky130_fd_sc_hd__o31a_1 _17163_ (.A1(_09140_),
    .A2(_08409_),
    .A3(_10048_),
    .B1(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__nor2_1 _17164_ (.A(_10161_),
    .B(_10163_),
    .Y(_10164_));
 sky130_fd_sc_hd__nand2_1 _17165_ (.A(_10161_),
    .B(_10163_),
    .Y(_10165_));
 sky130_fd_sc_hd__and2b_1 _17166_ (.A_N(_10164_),
    .B(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__xor2_1 _17167_ (.A(_10156_),
    .B(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__xnor2_1 _17168_ (.A(_10151_),
    .B(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__xnor2_1 _17169_ (.A(_10150_),
    .B(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__nand2_1 _17170_ (.A(_10058_),
    .B(_10061_),
    .Y(_10170_));
 sky130_fd_sc_hd__o31ai_2 _17171_ (.A1(_09647_),
    .A2(_09170_),
    .A3(_10062_),
    .B1(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__or2_1 _17172_ (.A(_08911_),
    .B(_09663_),
    .X(_10172_));
 sky130_fd_sc_hd__a21o_1 _17173_ (.A1(_09951_),
    .A2(_09952_),
    .B1(_08941_),
    .X(_10173_));
 sky130_fd_sc_hd__a2bb2oi_1 _17174_ (.A1_N(_10172_),
    .A2_N(_10173_),
    .B1(_10072_),
    .B2(_10070_),
    .Y(_10174_));
 sky130_fd_sc_hd__or3b_1 _17175_ (.A(_08876_),
    .B(_10069_),
    .C_N(_10061_),
    .X(_10175_));
 sky130_fd_sc_hd__o22ai_1 _17176_ (.A1(_08876_),
    .A2(_09534_),
    .B1(_10069_),
    .B2(_08875_),
    .Y(_10176_));
 sky130_fd_sc_hd__nand2_1 _17177_ (.A(_10175_),
    .B(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__nor2_1 _17178_ (.A(_09647_),
    .B(_09533_),
    .Y(_10178_));
 sky130_fd_sc_hd__xnor2_1 _17179_ (.A(_10177_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__xnor2_1 _17180_ (.A(_10174_),
    .B(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__xor2_1 _17181_ (.A(_10171_),
    .B(_10180_),
    .X(_10181_));
 sky130_fd_sc_hd__nor2_1 _17182_ (.A(_08360_),
    .B(_09663_),
    .Y(_10182_));
 sky130_fd_sc_hd__a21oi_1 _17183_ (.A1(_09947_),
    .A2(_09949_),
    .B1(_08911_),
    .Y(_10183_));
 sky130_fd_sc_hd__xnor2_1 _17184_ (.A(_10173_),
    .B(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__xor2_1 _17185_ (.A(_10182_),
    .B(_10184_),
    .X(_10185_));
 sky130_fd_sc_hd__xor2_1 _17186_ (.A(_10076_),
    .B(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__a21o_1 _17187_ (.A1(_10073_),
    .A2(_10076_),
    .B1(_10075_),
    .X(_10187_));
 sky130_fd_sc_hd__xor2_1 _17188_ (.A(_10186_),
    .B(_10187_),
    .X(_10188_));
 sky130_fd_sc_hd__xnor2_1 _17189_ (.A(_10181_),
    .B(_10188_),
    .Y(_10189_));
 sky130_fd_sc_hd__nor2_1 _17190_ (.A(_10077_),
    .B(_10079_),
    .Y(_10190_));
 sky130_fd_sc_hd__a21o_1 _17191_ (.A1(_10068_),
    .A2(_10080_),
    .B1(_10190_),
    .X(_10191_));
 sky130_fd_sc_hd__xnor2_1 _17192_ (.A(_10189_),
    .B(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__xnor2_1 _17193_ (.A(_10169_),
    .B(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__and2b_1 _17194_ (.A_N(_10081_),
    .B(_10083_),
    .X(_10194_));
 sky130_fd_sc_hd__a21oi_1 _17195_ (.A1(_10057_),
    .A2(_10084_),
    .B1(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__nor2_1 _17196_ (.A(_10193_),
    .B(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__and2_1 _17197_ (.A(_10193_),
    .B(_10195_),
    .X(_10197_));
 sky130_fd_sc_hd__nor2_1 _17198_ (.A(_10196_),
    .B(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__xnor2_1 _17199_ (.A(_10149_),
    .B(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__a21oi_1 _17200_ (.A1(_10035_),
    .A2(_10090_),
    .B1(_10088_),
    .Y(_10200_));
 sky130_fd_sc_hd__nor2_1 _17201_ (.A(_10199_),
    .B(_10200_),
    .Y(_10201_));
 sky130_fd_sc_hd__and2_1 _17202_ (.A(_10199_),
    .B(_10200_),
    .X(_10202_));
 sky130_fd_sc_hd__nor2_1 _17203_ (.A(_10201_),
    .B(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__xnor2_1 _17204_ (.A(_10119_),
    .B(_10203_),
    .Y(_10204_));
 sky130_fd_sc_hd__a21oi_1 _17205_ (.A1(_09997_),
    .A2(_10094_),
    .B1(_10092_),
    .Y(_10205_));
 sky130_fd_sc_hd__xor2_1 _17206_ (.A(_10204_),
    .B(_10205_),
    .X(_10206_));
 sky130_fd_sc_hd__nand2_1 _17207_ (.A(_09995_),
    .B(_10206_),
    .Y(_10207_));
 sky130_fd_sc_hd__or2_1 _17208_ (.A(_09995_),
    .B(_10206_),
    .X(_10208_));
 sky130_fd_sc_hd__nand2_1 _17209_ (.A(_10207_),
    .B(_10208_),
    .Y(_10209_));
 sky130_fd_sc_hd__a21oi_1 _17210_ (.A1(_09873_),
    .A2(_10099_),
    .B1(_10097_),
    .Y(_10210_));
 sky130_fd_sc_hd__or2_1 _17211_ (.A(_10209_),
    .B(_10210_),
    .X(_10211_));
 sky130_fd_sc_hd__nand2_1 _17212_ (.A(_10209_),
    .B(_10210_),
    .Y(_10212_));
 sky130_fd_sc_hd__and2_2 _17213_ (.A(_10211_),
    .B(_10212_),
    .X(_10213_));
 sky130_fd_sc_hd__a21o_1 _17214_ (.A1(_09992_),
    .A2(_09981_),
    .B1(_10100_),
    .X(_10214_));
 sky130_fd_sc_hd__a21o_1 _17215_ (.A1(_09984_),
    .A2(_10214_),
    .B1(_10102_),
    .X(_10215_));
 sky130_fd_sc_hd__o31a_4 _17216_ (.A1(_09986_),
    .A2(_09988_),
    .A3(_10103_),
    .B1(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__xnor2_4 _17217_ (.A(_10213_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__nand2_1 _17218_ (.A(_06101_),
    .B(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__inv_2 _17219_ (.A(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__nand2_1 _17220_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .Y(_10220_));
 sky130_fd_sc_hd__or2_1 _17221_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_10221_));
 sky130_fd_sc_hd__inv_2 _17222_ (.A(_10108_),
    .Y(_10222_));
 sky130_fd_sc_hd__a211o_1 _17223_ (.A1(_10220_),
    .A2(_10221_),
    .B1(_10222_),
    .C1(_10111_),
    .X(_10223_));
 sky130_fd_sc_hd__o211ai_2 _17224_ (.A1(_10222_),
    .A2(_10111_),
    .B1(_10220_),
    .C1(_10221_),
    .Y(_10224_));
 sky130_fd_sc_hd__a31o_1 _17225_ (.A1(_08101_),
    .A2(_10223_),
    .A3(_10224_),
    .B1(_09761_),
    .X(_10225_));
 sky130_fd_sc_hd__o22a_1 _17226_ (.A1(\rbzero.wall_tracer.trackDistX[2] ),
    .A2(_09805_),
    .B1(_10219_),
    .B2(_10225_),
    .X(_00541_));
 sky130_fd_sc_hd__or2_1 _17227_ (.A(_10204_),
    .B(_10205_),
    .X(_10226_));
 sky130_fd_sc_hd__nand2_1 _17228_ (.A(_10122_),
    .B(_10147_),
    .Y(_10227_));
 sky130_fd_sc_hd__or2b_1 _17229_ (.A(_10148_),
    .B_N(_10120_),
    .X(_10228_));
 sky130_fd_sc_hd__o2bb2a_1 _17230_ (.A1_N(_10129_),
    .A2_N(_10130_),
    .B1(_10127_),
    .B2(_10128_),
    .X(_10229_));
 sky130_fd_sc_hd__a21oi_1 _17231_ (.A1(_10227_),
    .A2(_10228_),
    .B1(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__and3_1 _17232_ (.A(_10227_),
    .B(_10228_),
    .C(_10229_),
    .X(_10231_));
 sky130_fd_sc_hd__nor2_1 _17233_ (.A(_10230_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__a21o_1 _17234_ (.A1(_10131_),
    .A2(_10146_),
    .B1(_10144_),
    .X(_10233_));
 sky130_fd_sc_hd__or2b_1 _17235_ (.A(_10168_),
    .B_N(_10150_),
    .X(_10234_));
 sky130_fd_sc_hd__a21bo_1 _17236_ (.A1(_10151_),
    .A2(_10167_),
    .B1_N(_10234_),
    .X(_10235_));
 sky130_fd_sc_hd__nor2_1 _17237_ (.A(_09503_),
    .B(_09342_),
    .Y(_10236_));
 sky130_fd_sc_hd__or2_1 _17238_ (.A(_09369_),
    .B(_09226_),
    .X(_10237_));
 sky130_fd_sc_hd__xnor2_1 _17239_ (.A(_10236_),
    .B(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__nor2_1 _17240_ (.A(_09127_),
    .B(_09469_),
    .Y(_10239_));
 sky130_fd_sc_hd__nand2_1 _17241_ (.A(_10238_),
    .B(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__or2_1 _17242_ (.A(_10238_),
    .B(_10239_),
    .X(_10241_));
 sky130_fd_sc_hd__nand2_1 _17243_ (.A(_10240_),
    .B(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__o31a_1 _17244_ (.A1(_09128_),
    .A2(_09469_),
    .A3(_10125_),
    .B1(_10124_),
    .X(_10243_));
 sky130_fd_sc_hd__xnor2_1 _17245_ (.A(_10242_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__nor2_1 _17246_ (.A(_08512_),
    .B(_09589_),
    .Y(_10245_));
 sky130_fd_sc_hd__xnor2_1 _17247_ (.A(_10244_),
    .B(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__a21bo_1 _17248_ (.A1(_10133_),
    .A2(_10136_),
    .B1_N(_10134_),
    .X(_10247_));
 sky130_fd_sc_hd__nand2_1 _17249_ (.A(_10040_),
    .B(_10152_),
    .Y(_10248_));
 sky130_fd_sc_hd__o22ai_1 _17250_ (.A1(_09910_),
    .A2(_08600_),
    .B1(_09056_),
    .B2(_08385_),
    .Y(_10249_));
 sky130_fd_sc_hd__or4_1 _17251_ (.A(_09910_),
    .B(_08385_),
    .C(_08599_),
    .D(_09056_),
    .X(_10250_));
 sky130_fd_sc_hd__nand2_1 _17252_ (.A(_10249_),
    .B(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__nor2_1 _17253_ (.A(_08649_),
    .B(_09110_),
    .Y(_10252_));
 sky130_fd_sc_hd__xor2_1 _17254_ (.A(_10251_),
    .B(_10252_),
    .X(_10253_));
 sky130_fd_sc_hd__a21oi_1 _17255_ (.A1(_10248_),
    .A2(_10154_),
    .B1(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__and3_1 _17256_ (.A(_10248_),
    .B(_10154_),
    .C(_10253_),
    .X(_10255_));
 sky130_fd_sc_hd__nor2_1 _17257_ (.A(_10254_),
    .B(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__xnor2_1 _17258_ (.A(_10247_),
    .B(_10256_),
    .Y(_10257_));
 sky130_fd_sc_hd__a21oi_1 _17259_ (.A1(_10132_),
    .A2(_10141_),
    .B1(_10139_),
    .Y(_10258_));
 sky130_fd_sc_hd__nor2_1 _17260_ (.A(_10257_),
    .B(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__and2_1 _17261_ (.A(_10257_),
    .B(_10258_),
    .X(_10260_));
 sky130_fd_sc_hd__nor2_1 _17262_ (.A(_10259_),
    .B(_10260_),
    .Y(_10261_));
 sky130_fd_sc_hd__xor2_1 _17263_ (.A(_10246_),
    .B(_10261_),
    .X(_10262_));
 sky130_fd_sc_hd__xnor2_1 _17264_ (.A(_10235_),
    .B(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__xnor2_1 _17265_ (.A(_10233_),
    .B(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__a21o_1 _17266_ (.A1(_10156_),
    .A2(_10165_),
    .B1(_10164_),
    .X(_10265_));
 sky130_fd_sc_hd__and2b_1 _17267_ (.A_N(_10174_),
    .B(_10179_),
    .X(_10266_));
 sky130_fd_sc_hd__a21oi_1 _17268_ (.A1(_10171_),
    .A2(_10180_),
    .B1(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__clkbuf_4 _17269_ (.A(_08368_),
    .X(_10268_));
 sky130_fd_sc_hd__nand2_2 _17270_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08318_),
    .Y(_10269_));
 sky130_fd_sc_hd__or2_1 _17271_ (.A(_10269_),
    .B(_08405_),
    .X(_10270_));
 sky130_fd_sc_hd__and3_1 _17272_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08523_),
    .C(_08424_),
    .X(_10271_));
 sky130_fd_sc_hd__xor2_1 _17273_ (.A(_10270_),
    .B(_10271_),
    .X(_10272_));
 sky130_fd_sc_hd__or3_1 _17274_ (.A(_10268_),
    .B(_08534_),
    .C(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__o21ai_1 _17275_ (.A1(_10268_),
    .A2(_09132_),
    .B1(_10272_),
    .Y(_10274_));
 sky130_fd_sc_hd__and2_1 _17276_ (.A(_10273_),
    .B(_10274_),
    .X(_10275_));
 sky130_fd_sc_hd__nor2_1 _17277_ (.A(_09506_),
    .B(_09533_),
    .Y(_10276_));
 sky130_fd_sc_hd__o22a_1 _17278_ (.A1(_09506_),
    .A2(_09170_),
    .B1(_09533_),
    .B2(_08797_),
    .X(_10277_));
 sky130_fd_sc_hd__a21oi_1 _17279_ (.A1(_10158_),
    .A2(_10276_),
    .B1(_10277_),
    .Y(_10278_));
 sky130_fd_sc_hd__buf_2 _17280_ (.A(_08454_),
    .X(_10279_));
 sky130_fd_sc_hd__a21oi_1 _17281_ (.A1(_10279_),
    .A2(_09025_),
    .B1(_09140_),
    .Y(_10280_));
 sky130_fd_sc_hd__xnor2_1 _17282_ (.A(_10278_),
    .B(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__o2bb2a_1 _17283_ (.A1_N(_10157_),
    .A2_N(_10158_),
    .B1(_10159_),
    .B2(_10160_),
    .X(_10282_));
 sky130_fd_sc_hd__xor2_1 _17284_ (.A(_10281_),
    .B(_10282_),
    .X(_10283_));
 sky130_fd_sc_hd__xnor2_1 _17285_ (.A(_10275_),
    .B(_10283_),
    .Y(_10284_));
 sky130_fd_sc_hd__xnor2_1 _17286_ (.A(_10267_),
    .B(_10284_),
    .Y(_10285_));
 sky130_fd_sc_hd__xnor2_1 _17287_ (.A(_10265_),
    .B(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__a21bo_1 _17288_ (.A1(_10176_),
    .A2(_10178_),
    .B1_N(_10175_),
    .X(_10287_));
 sky130_fd_sc_hd__and2_1 _17289_ (.A(_09951_),
    .B(_09952_),
    .X(_10288_));
 sky130_fd_sc_hd__buf_2 _17290_ (.A(_10288_),
    .X(_10289_));
 sky130_fd_sc_hd__a211o_2 _17291_ (.A1(_09947_),
    .A2(_09949_),
    .B1(_08191_),
    .C1(_08171_),
    .X(_10290_));
 sky130_fd_sc_hd__a2bb2o_1 _17292_ (.A1_N(_10289_),
    .A2_N(_10290_),
    .B1(_10184_),
    .B2(_10182_),
    .X(_10291_));
 sky130_fd_sc_hd__nor2_1 _17293_ (.A(_08876_),
    .B(_09540_),
    .Y(_10292_));
 sky130_fd_sc_hd__nor2_1 _17294_ (.A(_08875_),
    .B(_09663_),
    .Y(_10293_));
 sky130_fd_sc_hd__xnor2_1 _17295_ (.A(_10292_),
    .B(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__nor2_1 _17296_ (.A(_08394_),
    .B(_09534_),
    .Y(_10295_));
 sky130_fd_sc_hd__xnor2_1 _17297_ (.A(_10294_),
    .B(_10295_),
    .Y(_10296_));
 sky130_fd_sc_hd__xnor2_1 _17298_ (.A(_10291_),
    .B(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__xnor2_1 _17299_ (.A(_10287_),
    .B(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__or2_1 _17300_ (.A(_08360_),
    .B(_10288_),
    .X(_10299_));
 sky130_fd_sc_hd__and2_1 _17301_ (.A(_08399_),
    .B(_08412_),
    .X(_10300_));
 sky130_fd_sc_hd__and2_1 _17302_ (.A(_09947_),
    .B(_09949_),
    .X(_10301_));
 sky130_fd_sc_hd__clkbuf_2 _17303_ (.A(_10301_),
    .X(_10302_));
 sky130_fd_sc_hd__or3b_1 _17304_ (.A(_10300_),
    .B(_10302_),
    .C_N(_10290_),
    .X(_10303_));
 sky130_fd_sc_hd__clkbuf_2 _17305_ (.A(_10303_),
    .X(_10304_));
 sky130_fd_sc_hd__xor2_1 _17306_ (.A(_10299_),
    .B(_10304_),
    .X(_10305_));
 sky130_fd_sc_hd__xnor2_1 _17307_ (.A(_10076_),
    .B(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__a21oi_1 _17308_ (.A1(_10076_),
    .A2(_10185_),
    .B1(_10075_),
    .Y(_10307_));
 sky130_fd_sc_hd__xor2_1 _17309_ (.A(_10306_),
    .B(_10307_),
    .X(_10308_));
 sky130_fd_sc_hd__xnor2_1 _17310_ (.A(_10298_),
    .B(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(_10186_),
    .B(_10187_),
    .Y(_10310_));
 sky130_fd_sc_hd__a21bo_1 _17312_ (.A1(_10181_),
    .A2(_10188_),
    .B1_N(_10310_),
    .X(_10311_));
 sky130_fd_sc_hd__xnor2_1 _17313_ (.A(_10309_),
    .B(_10311_),
    .Y(_10312_));
 sky130_fd_sc_hd__xnor2_1 _17314_ (.A(_10286_),
    .B(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__and2b_1 _17315_ (.A_N(_10189_),
    .B(_10191_),
    .X(_10314_));
 sky130_fd_sc_hd__a21oi_1 _17316_ (.A1(_10169_),
    .A2(_10192_),
    .B1(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__nor2_1 _17317_ (.A(_10313_),
    .B(_10315_),
    .Y(_10316_));
 sky130_fd_sc_hd__and2_1 _17318_ (.A(_10313_),
    .B(_10315_),
    .X(_10317_));
 sky130_fd_sc_hd__nor2_1 _17319_ (.A(_10316_),
    .B(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__xnor2_1 _17320_ (.A(_10264_),
    .B(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__a21oi_1 _17321_ (.A1(_10149_),
    .A2(_10198_),
    .B1(_10196_),
    .Y(_10320_));
 sky130_fd_sc_hd__xor2_1 _17322_ (.A(_10319_),
    .B(_10320_),
    .X(_10321_));
 sky130_fd_sc_hd__nand2_1 _17323_ (.A(_10232_),
    .B(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__or2_1 _17324_ (.A(_10232_),
    .B(_10321_),
    .X(_10323_));
 sky130_fd_sc_hd__nand2_1 _17325_ (.A(_10322_),
    .B(_10323_),
    .Y(_10324_));
 sky130_fd_sc_hd__a21oi_1 _17326_ (.A1(_10119_),
    .A2(_10203_),
    .B1(_10201_),
    .Y(_10325_));
 sky130_fd_sc_hd__xor2_1 _17327_ (.A(_10324_),
    .B(_10325_),
    .X(_10326_));
 sky130_fd_sc_hd__nand2_1 _17328_ (.A(_10117_),
    .B(_10326_),
    .Y(_10327_));
 sky130_fd_sc_hd__or2_1 _17329_ (.A(_10117_),
    .B(_10326_),
    .X(_10328_));
 sky130_fd_sc_hd__nand2_1 _17330_ (.A(_10327_),
    .B(_10328_),
    .Y(_10329_));
 sky130_fd_sc_hd__a21o_1 _17331_ (.A1(_10226_),
    .A2(_10207_),
    .B1(_10329_),
    .X(_10330_));
 sky130_fd_sc_hd__and3_1 _17332_ (.A(_10226_),
    .B(_10207_),
    .C(_10329_),
    .X(_10331_));
 sky130_fd_sc_hd__inv_2 _17333_ (.A(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__nand2_1 _17334_ (.A(_10330_),
    .B(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__inv_2 _17335_ (.A(_10213_),
    .Y(_10334_));
 sky130_fd_sc_hd__o21a_1 _17336_ (.A1(_10334_),
    .A2(_10216_),
    .B1(_10211_),
    .X(_10335_));
 sky130_fd_sc_hd__a21oi_1 _17337_ (.A1(_10333_),
    .A2(_10335_),
    .B1(_08101_),
    .Y(_10336_));
 sky130_fd_sc_hd__o21ai_4 _17338_ (.A1(_10333_),
    .A2(_10335_),
    .B1(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__clkbuf_4 _17339_ (.A(_09824_),
    .X(_10338_));
 sky130_fd_sc_hd__and2_1 _17340_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_10339_));
 sky130_fd_sc_hd__nor2_1 _17341_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_10340_));
 sky130_fd_sc_hd__o211a_1 _17342_ (.A1(_10339_),
    .A2(_10340_),
    .B1(_10220_),
    .C1(_10224_),
    .X(_10341_));
 sky130_fd_sc_hd__a211oi_2 _17343_ (.A1(_10220_),
    .A2(_10224_),
    .B1(_10339_),
    .C1(_10340_),
    .Y(_10342_));
 sky130_fd_sc_hd__o31a_1 _17344_ (.A1(_10338_),
    .A2(_10341_),
    .A3(_10342_),
    .B1(_09794_),
    .X(_10343_));
 sky130_fd_sc_hd__o2bb2a_1 _17345_ (.A1_N(_10337_),
    .A2_N(_10343_),
    .B1(\rbzero.wall_tracer.trackDistX[3] ),
    .B2(_09805_),
    .X(_00542_));
 sky130_fd_sc_hd__nand2_1 _17346_ (.A(_10235_),
    .B(_10262_),
    .Y(_10344_));
 sky130_fd_sc_hd__or2b_1 _17347_ (.A(_10263_),
    .B_N(_10233_),
    .X(_10345_));
 sky130_fd_sc_hd__o32a_1 _17348_ (.A1(_08512_),
    .A2(_09589_),
    .A3(_10244_),
    .B1(_10243_),
    .B2(_10242_),
    .X(_10346_));
 sky130_fd_sc_hd__a21oi_2 _17349_ (.A1(_10344_),
    .A2(_10345_),
    .B1(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__and3_1 _17350_ (.A(_10344_),
    .B(_10345_),
    .C(_10346_),
    .X(_10348_));
 sky130_fd_sc_hd__nor2_1 _17351_ (.A(_10347_),
    .B(_10348_),
    .Y(_10349_));
 sky130_fd_sc_hd__a21o_1 _17352_ (.A1(_10246_),
    .A2(_10261_),
    .B1(_10259_),
    .X(_10350_));
 sky130_fd_sc_hd__or2_1 _17353_ (.A(_10267_),
    .B(_10284_),
    .X(_10351_));
 sky130_fd_sc_hd__or2b_1 _17354_ (.A(_10285_),
    .B_N(_10265_),
    .X(_10352_));
 sky130_fd_sc_hd__o22a_1 _17355_ (.A1(_09915_),
    .A2(_09227_),
    .B1(_09341_),
    .B2(_09369_),
    .X(_10353_));
 sky130_fd_sc_hd__or3_1 _17356_ (.A(_09915_),
    .B(_09341_),
    .C(_10237_),
    .X(_10354_));
 sky130_fd_sc_hd__or2b_1 _17357_ (.A(_10353_),
    .B_N(_10354_),
    .X(_10355_));
 sky130_fd_sc_hd__nor2_1 _17358_ (.A(_09503_),
    .B(_09469_),
    .Y(_10356_));
 sky130_fd_sc_hd__xor2_1 _17359_ (.A(_10355_),
    .B(_10356_),
    .X(_10357_));
 sky130_fd_sc_hd__o31a_1 _17360_ (.A1(_09503_),
    .A2(_09342_),
    .A3(_10237_),
    .B1(_10240_),
    .X(_10358_));
 sky130_fd_sc_hd__xor2_1 _17361_ (.A(_10357_),
    .B(_10358_),
    .X(_10359_));
 sky130_fd_sc_hd__and2_1 _17362_ (.A(_09127_),
    .B(_09669_),
    .X(_10360_));
 sky130_fd_sc_hd__xor2_1 _17363_ (.A(_10359_),
    .B(_10360_),
    .X(_10361_));
 sky130_fd_sc_hd__a21bo_1 _17364_ (.A1(_10249_),
    .A2(_10252_),
    .B1_N(_10250_),
    .X(_10362_));
 sky130_fd_sc_hd__or2b_1 _17365_ (.A(_10270_),
    .B_N(_10271_),
    .X(_10363_));
 sky130_fd_sc_hd__nand2_1 _17366_ (.A(_10363_),
    .B(_10273_),
    .Y(_10364_));
 sky130_fd_sc_hd__or2_1 _17367_ (.A(_08374_),
    .B(_09055_),
    .X(_10365_));
 sky130_fd_sc_hd__or3_1 _17368_ (.A(_08368_),
    .B(_08600_),
    .C(_10365_),
    .X(_10366_));
 sky130_fd_sc_hd__o21ai_1 _17369_ (.A1(_08368_),
    .A2(_08600_),
    .B1(_10365_),
    .Y(_10367_));
 sky130_fd_sc_hd__nand2_1 _17370_ (.A(_10366_),
    .B(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__or2_1 _17371_ (.A(_10038_),
    .B(_09110_),
    .X(_10369_));
 sky130_fd_sc_hd__xnor2_1 _17372_ (.A(_10368_),
    .B(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__xnor2_1 _17373_ (.A(_10364_),
    .B(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__xnor2_1 _17374_ (.A(_10362_),
    .B(_10371_),
    .Y(_10372_));
 sky130_fd_sc_hd__a21oi_1 _17375_ (.A1(_10247_),
    .A2(_10256_),
    .B1(_10254_),
    .Y(_10373_));
 sky130_fd_sc_hd__nor2_1 _17376_ (.A(_10372_),
    .B(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__and2_1 _17377_ (.A(_10372_),
    .B(_10373_),
    .X(_10375_));
 sky130_fd_sc_hd__nor2_1 _17378_ (.A(_10374_),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__xnor2_1 _17379_ (.A(_10361_),
    .B(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__a21o_1 _17380_ (.A1(_10351_),
    .A2(_10352_),
    .B1(_10377_),
    .X(_10378_));
 sky130_fd_sc_hd__nand3_1 _17381_ (.A(_10351_),
    .B(_10352_),
    .C(_10377_),
    .Y(_10379_));
 sky130_fd_sc_hd__nand2_1 _17382_ (.A(_10378_),
    .B(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__xnor2_1 _17383_ (.A(_10350_),
    .B(_10380_),
    .Y(_10381_));
 sky130_fd_sc_hd__nor2_1 _17384_ (.A(_10281_),
    .B(_10282_),
    .Y(_10382_));
 sky130_fd_sc_hd__a21o_1 _17385_ (.A1(_10275_),
    .A2(_10283_),
    .B1(_10382_),
    .X(_10383_));
 sky130_fd_sc_hd__or2b_1 _17386_ (.A(_10297_),
    .B_N(_10287_),
    .X(_10384_));
 sky130_fd_sc_hd__a21bo_1 _17387_ (.A1(_10291_),
    .A2(_10296_),
    .B1_N(_10384_),
    .X(_10385_));
 sky130_fd_sc_hd__nand2_2 _17388_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08318_),
    .Y(_10386_));
 sky130_fd_sc_hd__nand2_1 _17389_ (.A(_08523_),
    .B(_08424_),
    .Y(_10387_));
 sky130_fd_sc_hd__or4_1 _17390_ (.A(_10386_),
    .B(_10269_),
    .C(_10387_),
    .D(_10279_),
    .X(_10388_));
 sky130_fd_sc_hd__and2_1 _17391_ (.A(_08523_),
    .B(_08424_),
    .X(_10389_));
 sky130_fd_sc_hd__nor2_1 _17392_ (.A(_10386_),
    .B(_08454_),
    .Y(_10390_));
 sky130_fd_sc_hd__a31o_1 _17393_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_08318_),
    .A3(_10389_),
    .B1(_10390_),
    .X(_10391_));
 sky130_fd_sc_hd__nand2_1 _17394_ (.A(_10388_),
    .B(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__or2_1 _17395_ (.A(_08479_),
    .B(_09132_),
    .X(_10393_));
 sky130_fd_sc_hd__xor2_2 _17396_ (.A(_10392_),
    .B(_10393_),
    .X(_10394_));
 sky130_fd_sc_hd__nor2_1 _17397_ (.A(_08797_),
    .B(_09534_),
    .Y(_10395_));
 sky130_fd_sc_hd__xnor2_1 _17398_ (.A(_10276_),
    .B(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__nor2_1 _17399_ (.A(_09140_),
    .B(_09170_),
    .Y(_10397_));
 sky130_fd_sc_hd__xor2_1 _17400_ (.A(_10396_),
    .B(_10397_),
    .X(_10398_));
 sky130_fd_sc_hd__a22oi_1 _17401_ (.A1(_10158_),
    .A2(_10276_),
    .B1(_10278_),
    .B2(_10280_),
    .Y(_10399_));
 sky130_fd_sc_hd__nor2_1 _17402_ (.A(_10398_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__and2_1 _17403_ (.A(_10398_),
    .B(_10399_),
    .X(_10401_));
 sky130_fd_sc_hd__nor2_1 _17404_ (.A(_10400_),
    .B(_10401_),
    .Y(_10402_));
 sky130_fd_sc_hd__xnor2_1 _17405_ (.A(_10394_),
    .B(_10402_),
    .Y(_10403_));
 sky130_fd_sc_hd__xor2_1 _17406_ (.A(_10385_),
    .B(_10403_),
    .X(_10404_));
 sky130_fd_sc_hd__xnor2_1 _17407_ (.A(_10383_),
    .B(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__or3_1 _17408_ (.A(_09647_),
    .B(_09534_),
    .C(_10294_),
    .X(_10406_));
 sky130_fd_sc_hd__a21bo_1 _17409_ (.A1(_10292_),
    .A2(_10293_),
    .B1_N(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__o21ai_1 _17410_ (.A1(_10299_),
    .A2(_10304_),
    .B1(_10290_),
    .Y(_10408_));
 sky130_fd_sc_hd__or2_1 _17411_ (.A(_08876_),
    .B(_09662_),
    .X(_10409_));
 sky130_fd_sc_hd__or3_1 _17412_ (.A(_08875_),
    .B(_10288_),
    .C(_10409_),
    .X(_10410_));
 sky130_fd_sc_hd__o21ai_1 _17413_ (.A1(_08875_),
    .A2(_10289_),
    .B1(_10409_),
    .Y(_10411_));
 sky130_fd_sc_hd__nand2_1 _17414_ (.A(_10410_),
    .B(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__or2_1 _17415_ (.A(_09647_),
    .B(_10069_),
    .X(_10413_));
 sky130_fd_sc_hd__xnor2_1 _17416_ (.A(_10412_),
    .B(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__xor2_1 _17417_ (.A(_10408_),
    .B(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__xnor2_1 _17418_ (.A(_10407_),
    .B(_10415_),
    .Y(_10416_));
 sky130_fd_sc_hd__a21o_1 _17419_ (.A1(_10076_),
    .A2(_10305_),
    .B1(_10075_),
    .X(_10417_));
 sky130_fd_sc_hd__nor2_1 _17420_ (.A(_08360_),
    .B(_10302_),
    .Y(_10418_));
 sky130_fd_sc_hd__mux2_2 _17421_ (.A0(_08360_),
    .A1(_10418_),
    .S(_10304_),
    .X(_10419_));
 sky130_fd_sc_hd__xor2_1 _17422_ (.A(_10076_),
    .B(_10419_),
    .X(_10420_));
 sky130_fd_sc_hd__and2_1 _17423_ (.A(_10417_),
    .B(_10420_),
    .X(_10421_));
 sky130_fd_sc_hd__nor2_1 _17424_ (.A(_10417_),
    .B(_10420_),
    .Y(_10422_));
 sky130_fd_sc_hd__nor2_1 _17425_ (.A(_10421_),
    .B(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__xnor2_1 _17426_ (.A(_10416_),
    .B(_10423_),
    .Y(_10424_));
 sky130_fd_sc_hd__nor2_1 _17427_ (.A(_10306_),
    .B(_10307_),
    .Y(_10425_));
 sky130_fd_sc_hd__a21oi_1 _17428_ (.A1(_10298_),
    .A2(_10308_),
    .B1(_10425_),
    .Y(_10426_));
 sky130_fd_sc_hd__xor2_1 _17429_ (.A(_10424_),
    .B(_10426_),
    .X(_10427_));
 sky130_fd_sc_hd__xnor2_1 _17430_ (.A(_10405_),
    .B(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__and2b_1 _17431_ (.A_N(_10309_),
    .B(_10311_),
    .X(_10429_));
 sky130_fd_sc_hd__a21oi_1 _17432_ (.A1(_10286_),
    .A2(_10312_),
    .B1(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__xor2_1 _17433_ (.A(_10428_),
    .B(_10430_),
    .X(_10431_));
 sky130_fd_sc_hd__xnor2_1 _17434_ (.A(_10381_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__a21oi_1 _17435_ (.A1(_10264_),
    .A2(_10318_),
    .B1(_10316_),
    .Y(_10433_));
 sky130_fd_sc_hd__nor2_1 _17436_ (.A(_10432_),
    .B(_10433_),
    .Y(_10434_));
 sky130_fd_sc_hd__nand2_1 _17437_ (.A(_10432_),
    .B(_10433_),
    .Y(_10435_));
 sky130_fd_sc_hd__and2b_1 _17438_ (.A_N(_10434_),
    .B(_10435_),
    .X(_10436_));
 sky130_fd_sc_hd__xnor2_1 _17439_ (.A(_10349_),
    .B(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__o21a_1 _17440_ (.A1(_10319_),
    .A2(_10320_),
    .B1(_10322_),
    .X(_10438_));
 sky130_fd_sc_hd__xor2_1 _17441_ (.A(_10437_),
    .B(_10438_),
    .X(_10439_));
 sky130_fd_sc_hd__nand2_1 _17442_ (.A(_10230_),
    .B(_10439_),
    .Y(_10440_));
 sky130_fd_sc_hd__or2_1 _17443_ (.A(_10230_),
    .B(_10439_),
    .X(_10441_));
 sky130_fd_sc_hd__nand2_1 _17444_ (.A(_10440_),
    .B(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__o21a_1 _17445_ (.A1(_10324_),
    .A2(_10325_),
    .B1(_10327_),
    .X(_10443_));
 sky130_fd_sc_hd__xor2_2 _17446_ (.A(_10442_),
    .B(_10443_),
    .X(_10444_));
 sky130_fd_sc_hd__nand3_1 _17447_ (.A(_10213_),
    .B(_10330_),
    .C(_10332_),
    .Y(_10445_));
 sky130_fd_sc_hd__a21oi_1 _17448_ (.A1(_10211_),
    .A2(_10330_),
    .B1(_10331_),
    .Y(_10446_));
 sky130_fd_sc_hd__o21bai_2 _17449_ (.A1(_10216_),
    .A2(_10445_),
    .B1_N(_10446_),
    .Y(_10447_));
 sky130_fd_sc_hd__a21oi_1 _17450_ (.A1(_10444_),
    .A2(_10447_),
    .B1(_08101_),
    .Y(_10448_));
 sky130_fd_sc_hd__o21ai_4 _17451_ (.A1(_10444_),
    .A2(_10447_),
    .B1(_10448_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _17452_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_01653_));
 sky130_fd_sc_hd__or2_1 _17453_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_01654_));
 sky130_fd_sc_hd__o211a_1 _17454_ (.A1(_10339_),
    .A2(_10342_),
    .B1(_01653_),
    .C1(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__a211oi_1 _17455_ (.A1(_01653_),
    .A2(_01654_),
    .B1(_10339_),
    .C1(_10342_),
    .Y(_01656_));
 sky130_fd_sc_hd__o31a_1 _17456_ (.A1(_10338_),
    .A2(_01655_),
    .A3(_01656_),
    .B1(_09794_),
    .X(_01657_));
 sky130_fd_sc_hd__o2bb2a_1 _17457_ (.A1_N(_01652_),
    .A2_N(_01657_),
    .B1(\rbzero.wall_tracer.trackDistX[4] ),
    .B2(_09805_),
    .X(_00543_));
 sky130_fd_sc_hd__or2_1 _17458_ (.A(_10437_),
    .B(_10438_),
    .X(_01658_));
 sky130_fd_sc_hd__or2b_1 _17459_ (.A(_10380_),
    .B_N(_10350_),
    .X(_01659_));
 sky130_fd_sc_hd__o2bb2a_1 _17460_ (.A1_N(_10359_),
    .A2_N(_10360_),
    .B1(_10357_),
    .B2(_10358_),
    .X(_01660_));
 sky130_fd_sc_hd__a21oi_1 _17461_ (.A1(_10378_),
    .A2(_01659_),
    .B1(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__and3_1 _17462_ (.A(_10378_),
    .B(_01659_),
    .C(_01660_),
    .X(_01662_));
 sky130_fd_sc_hd__nor2_1 _17463_ (.A(_01661_),
    .B(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__a21o_1 _17464_ (.A1(_10361_),
    .A2(_10376_),
    .B1(_10374_),
    .X(_01664_));
 sky130_fd_sc_hd__or2b_1 _17465_ (.A(_10403_),
    .B_N(_10385_),
    .X(_01665_));
 sky130_fd_sc_hd__or2b_1 _17466_ (.A(_10404_),
    .B_N(_10383_),
    .X(_01666_));
 sky130_fd_sc_hd__or2_1 _17467_ (.A(_10038_),
    .B(_09341_),
    .X(_01667_));
 sky130_fd_sc_hd__o22ai_1 _17468_ (.A1(_10038_),
    .A2(_09227_),
    .B1(_09342_),
    .B2(_09915_),
    .Y(_01668_));
 sky130_fd_sc_hd__o31a_1 _17469_ (.A1(_09915_),
    .A2(_09227_),
    .A3(_01667_),
    .B1(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__nor2_1 _17470_ (.A(_09369_),
    .B(_09469_),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _17471_ (.A(_01669_),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__or2_1 _17472_ (.A(_01669_),
    .B(_01670_),
    .X(_01672_));
 sky130_fd_sc_hd__nand2_1 _17473_ (.A(_01671_),
    .B(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__o31a_1 _17474_ (.A1(_09503_),
    .A2(_09605_),
    .A3(_10353_),
    .B1(_10354_),
    .X(_01674_));
 sky130_fd_sc_hd__xnor2_1 _17475_ (.A(_01673_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_1 _17476_ (.A(_09503_),
    .B(_09869_),
    .Y(_01676_));
 sky130_fd_sc_hd__xor2_1 _17477_ (.A(_01675_),
    .B(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__o31ai_2 _17478_ (.A1(_10038_),
    .A2(_09111_),
    .A3(_10368_),
    .B1(_10366_),
    .Y(_01678_));
 sky130_fd_sc_hd__o21ai_1 _17479_ (.A1(_10392_),
    .A2(_10393_),
    .B1(_10388_),
    .Y(_01679_));
 sky130_fd_sc_hd__or2_1 _17480_ (.A(_08479_),
    .B(_08600_),
    .X(_01680_));
 sky130_fd_sc_hd__or3_1 _17481_ (.A(_08368_),
    .B(_09056_),
    .C(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__o21ai_1 _17482_ (.A1(_10268_),
    .A2(_09056_),
    .B1(_01680_),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _17483_ (.A(_01681_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__nor2_1 _17484_ (.A(_09911_),
    .B(_09111_),
    .Y(_01684_));
 sky130_fd_sc_hd__xor2_1 _17485_ (.A(_01683_),
    .B(_01684_),
    .X(_01685_));
 sky130_fd_sc_hd__xnor2_1 _17486_ (.A(_01679_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__xnor2_1 _17487_ (.A(_01678_),
    .B(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__a21oi_1 _17488_ (.A1(_10363_),
    .A2(_10273_),
    .B1(_10370_),
    .Y(_01688_));
 sky130_fd_sc_hd__a21oi_1 _17489_ (.A1(_10362_),
    .A2(_10371_),
    .B1(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__nor2_1 _17490_ (.A(_01687_),
    .B(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__and2_1 _17491_ (.A(_01687_),
    .B(_01689_),
    .X(_01691_));
 sky130_fd_sc_hd__nor2_1 _17492_ (.A(_01690_),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__xnor2_1 _17493_ (.A(_01677_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__a21o_1 _17494_ (.A1(_01665_),
    .A2(_01666_),
    .B1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__nand3_1 _17495_ (.A(_01665_),
    .B(_01666_),
    .C(_01693_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _17496_ (.A(_01694_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__xnor2_1 _17497_ (.A(_01664_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__a21o_1 _17498_ (.A1(_10394_),
    .A2(_10402_),
    .B1(_10400_),
    .X(_01698_));
 sky130_fd_sc_hd__or2b_1 _17499_ (.A(_10414_),
    .B_N(_10408_),
    .X(_01699_));
 sky130_fd_sc_hd__or2b_1 _17500_ (.A(_10415_),
    .B_N(_10407_),
    .X(_01700_));
 sky130_fd_sc_hd__nor2_2 _17501_ (.A(_10269_),
    .B(_09295_),
    .Y(_01701_));
 sky130_fd_sc_hd__o22a_1 _17502_ (.A1(_10269_),
    .A2(_10279_),
    .B1(_09295_),
    .B2(_10386_),
    .X(_01702_));
 sky130_fd_sc_hd__a21oi_2 _17503_ (.A1(_10390_),
    .A2(_01701_),
    .B1(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__and3_1 _17504_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08523_),
    .C(_08424_),
    .X(_01704_));
 sky130_fd_sc_hd__xor2_2 _17505_ (.A(_01703_),
    .B(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__or4_1 _17506_ (.A(_08797_),
    .B(_09506_),
    .C(_09534_),
    .D(_10069_),
    .X(_01706_));
 sky130_fd_sc_hd__o22ai_1 _17507_ (.A1(_09506_),
    .A2(_09534_),
    .B1(_10069_),
    .B2(_08798_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _17508_ (.A(_01706_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__nor2_1 _17509_ (.A(_09512_),
    .B(_09533_),
    .Y(_01709_));
 sky130_fd_sc_hd__xor2_1 _17510_ (.A(_01708_),
    .B(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__nand2_1 _17511_ (.A(_10276_),
    .B(_10395_),
    .Y(_01711_));
 sky130_fd_sc_hd__o31a_1 _17512_ (.A1(_09512_),
    .A2(_09170_),
    .A3(_10396_),
    .B1(_01711_),
    .X(_01712_));
 sky130_fd_sc_hd__nor2_1 _17513_ (.A(_01710_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__and2_1 _17514_ (.A(_01710_),
    .B(_01712_),
    .X(_01714_));
 sky130_fd_sc_hd__nor2_1 _17515_ (.A(_01713_),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__xnor2_1 _17516_ (.A(_01705_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__a21o_1 _17517_ (.A1(_01699_),
    .A2(_01700_),
    .B1(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__nand3_1 _17518_ (.A(_01699_),
    .B(_01700_),
    .C(_01716_),
    .Y(_01718_));
 sky130_fd_sc_hd__nand2_1 _17519_ (.A(_01717_),
    .B(_01718_),
    .Y(_01719_));
 sky130_fd_sc_hd__xnor2_1 _17520_ (.A(_01698_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__o21ai_1 _17521_ (.A1(_10412_),
    .A2(_10413_),
    .B1(_10410_),
    .Y(_01721_));
 sky130_fd_sc_hd__o21ai_4 _17522_ (.A1(_08360_),
    .A2(_10304_),
    .B1(_10290_),
    .Y(_01722_));
 sky130_fd_sc_hd__or3_1 _17523_ (.A(_08875_),
    .B(_08876_),
    .C(_10302_),
    .X(_01723_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(_09951_),
    .B(_09952_),
    .Y(_01724_));
 sky130_fd_sc_hd__a2bb2o_1 _17525_ (.A1_N(_08875_),
    .A2_N(_10302_),
    .B1(_01724_),
    .B2(_08247_),
    .X(_01725_));
 sky130_fd_sc_hd__o21ai_1 _17526_ (.A1(_10289_),
    .A2(_01723_),
    .B1(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__nor2_1 _17527_ (.A(_09647_),
    .B(_09663_),
    .Y(_01727_));
 sky130_fd_sc_hd__xnor2_1 _17528_ (.A(_01726_),
    .B(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__xnor2_1 _17529_ (.A(_01722_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__xnor2_1 _17530_ (.A(_01721_),
    .B(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__nand2_1 _17531_ (.A(_10075_),
    .B(_10419_),
    .Y(_01731_));
 sky130_fd_sc_hd__nand3b_1 _17532_ (.A_N(_10419_),
    .B(_10074_),
    .C(_09950_),
    .Y(_01732_));
 sky130_fd_sc_hd__and2_1 _17533_ (.A(_01731_),
    .B(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__buf_2 _17534_ (.A(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__xnor2_1 _17535_ (.A(_01730_),
    .B(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__a21oi_1 _17536_ (.A1(_10416_),
    .A2(_10423_),
    .B1(_10421_),
    .Y(_01736_));
 sky130_fd_sc_hd__xor2_1 _17537_ (.A(_01735_),
    .B(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__xnor2_1 _17538_ (.A(_01720_),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__nor2_1 _17539_ (.A(_10424_),
    .B(_10426_),
    .Y(_01739_));
 sky130_fd_sc_hd__a21oi_1 _17540_ (.A1(_10405_),
    .A2(_10427_),
    .B1(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__xor2_1 _17541_ (.A(_01738_),
    .B(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__xnor2_1 _17542_ (.A(_01697_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__nor2_1 _17543_ (.A(_10428_),
    .B(_10430_),
    .Y(_01743_));
 sky130_fd_sc_hd__a21oi_1 _17544_ (.A1(_10381_),
    .A2(_10431_),
    .B1(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__xor2_1 _17545_ (.A(_01742_),
    .B(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__xnor2_1 _17546_ (.A(_01663_),
    .B(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__a21oi_1 _17547_ (.A1(_10349_),
    .A2(_10435_),
    .B1(_10434_),
    .Y(_01747_));
 sky130_fd_sc_hd__nor2_1 _17548_ (.A(_01746_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nand2_1 _17549_ (.A(_01746_),
    .B(_01747_),
    .Y(_01749_));
 sky130_fd_sc_hd__and2b_1 _17550_ (.A_N(_01748_),
    .B(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__xnor2_1 _17551_ (.A(_10347_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__and3_1 _17552_ (.A(_01658_),
    .B(_10440_),
    .C(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__a21oi_1 _17553_ (.A1(_01658_),
    .A2(_10440_),
    .B1(_01751_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_2 _17554_ (.A(_01752_),
    .B(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__or2_1 _17555_ (.A(_10442_),
    .B(_10443_),
    .X(_01755_));
 sky130_fd_sc_hd__a21boi_2 _17556_ (.A1(_10444_),
    .A2(_10447_),
    .B1_N(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__xnor2_4 _17557_ (.A(_01754_),
    .B(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_1 _17558_ (.A(_10107_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _17559_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_01759_));
 sky130_fd_sc_hd__and2_1 _17560_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_01760_));
 sky130_fd_sc_hd__a21oi_1 _17561_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(\rbzero.wall_tracer.stepDistX[4] ),
    .B1(_01655_),
    .Y(_01761_));
 sky130_fd_sc_hd__o21ai_1 _17562_ (.A1(_01759_),
    .A2(_01760_),
    .B1(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__o31a_1 _17563_ (.A1(_01759_),
    .A2(_01760_),
    .A3(_01761_),
    .B1(_08100_),
    .X(_01763_));
 sky130_fd_sc_hd__a21oi_1 _17564_ (.A1(_01762_),
    .A2(_01763_),
    .B1(_09763_),
    .Y(_01764_));
 sky130_fd_sc_hd__o2bb2a_1 _17565_ (.A1_N(_01758_),
    .A2_N(_01764_),
    .B1(\rbzero.wall_tracer.trackDistX[5] ),
    .B2(_09805_),
    .X(_00544_));
 sky130_fd_sc_hd__nor2_1 _17566_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01765_));
 sky130_fd_sc_hd__nand2_1 _17567_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01766_));
 sky130_fd_sc_hd__or2b_1 _17568_ (.A(_01765_),
    .B_N(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__o21ba_1 _17569_ (.A1(_01759_),
    .A2(_01761_),
    .B1_N(_01760_),
    .X(_01768_));
 sky130_fd_sc_hd__nor2_1 _17570_ (.A(_01767_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__a21o_1 _17571_ (.A1(_01767_),
    .A2(_01768_),
    .B1(_06102_),
    .X(_01770_));
 sky130_fd_sc_hd__or2b_1 _17572_ (.A(_01696_),
    .B_N(_01664_),
    .X(_01771_));
 sky130_fd_sc_hd__o22a_1 _17573_ (.A1(_01673_),
    .A2(_01674_),
    .B1(_01675_),
    .B2(_01676_),
    .X(_01772_));
 sky130_fd_sc_hd__a21oi_2 _17574_ (.A1(_01694_),
    .A2(_01771_),
    .B1(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__and3_1 _17575_ (.A(_01694_),
    .B(_01771_),
    .C(_01772_),
    .X(_01774_));
 sky130_fd_sc_hd__nor2_1 _17576_ (.A(_01773_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21o_1 _17577_ (.A1(_01677_),
    .A2(_01692_),
    .B1(_01690_),
    .X(_01776_));
 sky130_fd_sc_hd__or2b_1 _17578_ (.A(_01719_),
    .B_N(_01698_),
    .X(_01777_));
 sky130_fd_sc_hd__nor2_1 _17579_ (.A(_09911_),
    .B(_09228_),
    .Y(_01778_));
 sky130_fd_sc_hd__xnor2_1 _17580_ (.A(_01667_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__nor2_1 _17581_ (.A(_09915_),
    .B(_09605_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _17582_ (.A(_01779_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__or2_1 _17583_ (.A(_01779_),
    .B(_01780_),
    .X(_01782_));
 sky130_fd_sc_hd__nand2_1 _17584_ (.A(_01781_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__o31a_1 _17585_ (.A1(_09915_),
    .A2(_09228_),
    .A3(_01667_),
    .B1(_01671_),
    .X(_01784_));
 sky130_fd_sc_hd__nor2_1 _17586_ (.A(_01783_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__and2_1 _17587_ (.A(_01783_),
    .B(_01784_),
    .X(_01786_));
 sky130_fd_sc_hd__nor2_1 _17588_ (.A(_01785_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__and2_1 _17589_ (.A(_09369_),
    .B(_09869_),
    .X(_01788_));
 sky130_fd_sc_hd__xor2_1 _17590_ (.A(_01787_),
    .B(_01788_),
    .X(_01789_));
 sky130_fd_sc_hd__o31ai_2 _17591_ (.A1(_09911_),
    .A2(_09111_),
    .A3(_01683_),
    .B1(_01681_),
    .Y(_01790_));
 sky130_fd_sc_hd__nand2_1 _17592_ (.A(_10390_),
    .B(_01701_),
    .Y(_01791_));
 sky130_fd_sc_hd__nand2_1 _17593_ (.A(_01703_),
    .B(_01704_),
    .Y(_01792_));
 sky130_fd_sc_hd__or2_1 _17594_ (.A(_10268_),
    .B(_09111_),
    .X(_01793_));
 sky130_fd_sc_hd__nand2_1 _17595_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08318_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _17596_ (.A(_08405_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__a31o_1 _17597_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_08318_),
    .A3(_10389_),
    .B1(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__nand2_1 _17598_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_10389_),
    .Y(_01797_));
 sky130_fd_sc_hd__or2_1 _17599_ (.A(_01680_),
    .B(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__nand2_1 _17600_ (.A(_01796_),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__xnor2_1 _17601_ (.A(_01793_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__a21oi_1 _17602_ (.A1(_01791_),
    .A2(_01792_),
    .B1(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__and3_1 _17603_ (.A(_01791_),
    .B(_01792_),
    .C(_01800_),
    .X(_01802_));
 sky130_fd_sc_hd__nor2_1 _17604_ (.A(_01801_),
    .B(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__xnor2_1 _17605_ (.A(_01790_),
    .B(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__and2b_1 _17606_ (.A_N(_01685_),
    .B(_01679_),
    .X(_01805_));
 sky130_fd_sc_hd__a21oi_1 _17607_ (.A1(_01678_),
    .A2(_01686_),
    .B1(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__nor2_1 _17608_ (.A(_01804_),
    .B(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__and2_1 _17609_ (.A(_01804_),
    .B(_01806_),
    .X(_01808_));
 sky130_fd_sc_hd__nor2_1 _17610_ (.A(_01807_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__xnor2_1 _17611_ (.A(_01789_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__a21o_1 _17612_ (.A1(_01717_),
    .A2(_01777_),
    .B1(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__nand3_1 _17613_ (.A(_01717_),
    .B(_01777_),
    .C(_01810_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _17614_ (.A(_01811_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__xnor2_1 _17615_ (.A(_01776_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__a21o_1 _17616_ (.A1(_01705_),
    .A2(_01715_),
    .B1(_01713_),
    .X(_01815_));
 sky130_fd_sc_hd__or2b_1 _17617_ (.A(_01729_),
    .B_N(_01721_),
    .X(_01816_));
 sky130_fd_sc_hd__a21bo_1 _17618_ (.A1(_01722_),
    .A2(_01728_),
    .B1_N(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__nand2_2 _17619_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08318_),
    .Y(_01818_));
 sky130_fd_sc_hd__nor2_1 _17620_ (.A(_10386_),
    .B(_09286_),
    .Y(_01819_));
 sky130_fd_sc_hd__xnor2_1 _17621_ (.A(_01701_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__or3_1 _17622_ (.A(_10279_),
    .B(_01818_),
    .C(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__o21ai_1 _17623_ (.A1(_10279_),
    .A2(_01818_),
    .B1(_01820_),
    .Y(_01822_));
 sky130_fd_sc_hd__and2_1 _17624_ (.A(_01821_),
    .B(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__or2_1 _17625_ (.A(_09506_),
    .B(_09663_),
    .X(_01824_));
 sky130_fd_sc_hd__o22ai_1 _17626_ (.A1(_09506_),
    .A2(_10069_),
    .B1(_09663_),
    .B2(_08798_),
    .Y(_01825_));
 sky130_fd_sc_hd__o31ai_1 _17627_ (.A1(_08798_),
    .A2(_10069_),
    .A3(_01824_),
    .B1(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__or3_1 _17628_ (.A(_09512_),
    .B(_09534_),
    .C(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__o21ai_1 _17629_ (.A1(_09512_),
    .A2(_09534_),
    .B1(_01826_),
    .Y(_01828_));
 sky130_fd_sc_hd__nand2_1 _17630_ (.A(_01827_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__o31a_1 _17631_ (.A1(_09512_),
    .A2(_09533_),
    .A3(_01708_),
    .B1(_01706_),
    .X(_01830_));
 sky130_fd_sc_hd__nor2_1 _17632_ (.A(_01829_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__and2_1 _17633_ (.A(_01829_),
    .B(_01830_),
    .X(_01832_));
 sky130_fd_sc_hd__nor2_1 _17634_ (.A(_01831_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__xnor2_1 _17635_ (.A(_01823_),
    .B(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__xor2_1 _17636_ (.A(_01817_),
    .B(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__xnor2_1 _17637_ (.A(_01815_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__a2bb2o_1 _17638_ (.A1_N(_10289_),
    .A2_N(_01723_),
    .B1(_01727_),
    .B2(_01725_),
    .X(_01837_));
 sky130_fd_sc_hd__or2_1 _17639_ (.A(_09647_),
    .B(_10289_),
    .X(_01838_));
 sky130_fd_sc_hd__nand2_1 _17640_ (.A(_09947_),
    .B(_09949_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _17641_ (.A(_08875_),
    .B(_08876_),
    .Y(_01840_));
 sky130_fd_sc_hd__and3_1 _17642_ (.A(_01839_),
    .B(_01723_),
    .C(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__xnor2_1 _17643_ (.A(_01838_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__xor2_1 _17644_ (.A(_01722_),
    .B(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__nand2_1 _17645_ (.A(_01837_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__or2_1 _17646_ (.A(_01837_),
    .B(_01843_),
    .X(_01845_));
 sky130_fd_sc_hd__and2_1 _17647_ (.A(_01844_),
    .B(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__xnor2_1 _17648_ (.A(_01734_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__a21boi_1 _17649_ (.A1(_01730_),
    .A2(_01734_),
    .B1_N(_01731_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_1 _17650_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__and2_1 _17651_ (.A(_01847_),
    .B(_01848_),
    .X(_01850_));
 sky130_fd_sc_hd__nor2_1 _17652_ (.A(_01849_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__xnor2_1 _17653_ (.A(_01836_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _17654_ (.A(_01735_),
    .B(_01736_),
    .Y(_01853_));
 sky130_fd_sc_hd__a21oi_1 _17655_ (.A1(_01720_),
    .A2(_01737_),
    .B1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__xor2_1 _17656_ (.A(_01852_),
    .B(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__xnor2_1 _17657_ (.A(_01814_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _17658_ (.A(_01738_),
    .B(_01740_),
    .Y(_01857_));
 sky130_fd_sc_hd__a21oi_1 _17659_ (.A1(_01697_),
    .A2(_01741_),
    .B1(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__xor2_1 _17660_ (.A(_01856_),
    .B(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__xnor2_1 _17661_ (.A(_01775_),
    .B(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor2_1 _17662_ (.A(_01742_),
    .B(_01744_),
    .Y(_01861_));
 sky130_fd_sc_hd__a21oi_1 _17663_ (.A1(_01663_),
    .A2(_01745_),
    .B1(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__or2_1 _17664_ (.A(_01860_),
    .B(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__nand2_1 _17665_ (.A(_01860_),
    .B(_01862_),
    .Y(_01864_));
 sky130_fd_sc_hd__and2_1 _17666_ (.A(_01863_),
    .B(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__nand2_1 _17667_ (.A(_01661_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__or2_1 _17668_ (.A(_01661_),
    .B(_01865_),
    .X(_01867_));
 sky130_fd_sc_hd__nand2_1 _17669_ (.A(_01866_),
    .B(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__a21oi_1 _17670_ (.A1(_10347_),
    .A2(_01749_),
    .B1(_01748_),
    .Y(_01869_));
 sky130_fd_sc_hd__or2_4 _17671_ (.A(_01868_),
    .B(_01869_),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_1 _17672_ (.A(_01868_),
    .B(_01869_),
    .Y(_01871_));
 sky130_fd_sc_hd__nand2_1 _17673_ (.A(_01870_),
    .B(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__or3b_1 _17674_ (.A(_01752_),
    .B(_01753_),
    .C_N(_10444_),
    .X(_01873_));
 sky130_fd_sc_hd__or2b_1 _17675_ (.A(_01873_),
    .B_N(_10446_),
    .X(_01874_));
 sky130_fd_sc_hd__o31a_1 _17676_ (.A1(_10216_),
    .A2(_10445_),
    .A3(_01873_),
    .B1(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__o21ba_1 _17677_ (.A1(_01755_),
    .A2(_01752_),
    .B1_N(_01753_),
    .X(_01876_));
 sky130_fd_sc_hd__and3_2 _17678_ (.A(_01872_),
    .B(_01875_),
    .C(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__a21o_2 _17679_ (.A1(_01875_),
    .A2(_01876_),
    .B1(_01872_),
    .X(_01878_));
 sky130_fd_sc_hd__or3b_1 _17680_ (.A(_09784_),
    .B(_01877_),
    .C_N(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__o21ai_1 _17681_ (.A1(_01769_),
    .A2(_01770_),
    .B1(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__mux2_1 _17682_ (.A0(\rbzero.wall_tracer.trackDistX[6] ),
    .A1(_01880_),
    .S(_09826_),
    .X(_01881_));
 sky130_fd_sc_hd__clkbuf_1 _17683_ (.A(_01881_),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _17684_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_01882_));
 sky130_fd_sc_hd__nand2_1 _17685_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_01883_));
 sky130_fd_sc_hd__or2b_1 _17686_ (.A(_01882_),
    .B_N(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__o21a_1 _17687_ (.A1(_01765_),
    .A2(_01768_),
    .B1(_01766_),
    .X(_01885_));
 sky130_fd_sc_hd__nor2_1 _17688_ (.A(_01884_),
    .B(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__a21o_1 _17689_ (.A1(_01884_),
    .A2(_01885_),
    .B1(_06102_),
    .X(_01887_));
 sky130_fd_sc_hd__or2b_1 _17690_ (.A(_01813_),
    .B_N(_01776_),
    .X(_01888_));
 sky130_fd_sc_hd__a21oi_2 _17691_ (.A1(_01787_),
    .A2(_01788_),
    .B1(_01785_),
    .Y(_01889_));
 sky130_fd_sc_hd__a21oi_4 _17692_ (.A1(_01811_),
    .A2(_01888_),
    .B1(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__and3_1 _17693_ (.A(_01811_),
    .B(_01888_),
    .C(_01889_),
    .X(_01891_));
 sky130_fd_sc_hd__nor2_1 _17694_ (.A(_01890_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__a21o_1 _17695_ (.A1(_01789_),
    .A2(_01809_),
    .B1(_01807_),
    .X(_01893_));
 sky130_fd_sc_hd__or2b_1 _17696_ (.A(_01834_),
    .B_N(_01817_),
    .X(_01894_));
 sky130_fd_sc_hd__or2b_1 _17697_ (.A(_01835_),
    .B_N(_01815_),
    .X(_01895_));
 sky130_fd_sc_hd__nor2_1 _17698_ (.A(_08374_),
    .B(_09342_),
    .Y(_01896_));
 sky130_fd_sc_hd__nor2_1 _17699_ (.A(_10268_),
    .B(_09228_),
    .Y(_01897_));
 sky130_fd_sc_hd__xnor2_1 _17700_ (.A(_01896_),
    .B(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _17701_ (.A(_10038_),
    .B(_09605_),
    .Y(_01899_));
 sky130_fd_sc_hd__xor2_1 _17702_ (.A(_01898_),
    .B(_01899_),
    .X(_01900_));
 sky130_fd_sc_hd__o31a_1 _17703_ (.A1(_09911_),
    .A2(_09228_),
    .A3(_01667_),
    .B1(_01781_),
    .X(_01901_));
 sky130_fd_sc_hd__xor2_1 _17704_ (.A(_01900_),
    .B(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__and2_1 _17705_ (.A(_09915_),
    .B(_09869_),
    .X(_01903_));
 sky130_fd_sc_hd__xor2_1 _17706_ (.A(_01902_),
    .B(_01903_),
    .X(_01904_));
 sky130_fd_sc_hd__o21ai_1 _17707_ (.A1(_01793_),
    .A2(_01799_),
    .B1(_01798_),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_2 _17708_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08318_),
    .Y(_01906_));
 sky130_fd_sc_hd__or3_1 _17709_ (.A(_10279_),
    .B(_01906_),
    .C(_01797_),
    .X(_01907_));
 sky130_fd_sc_hd__o21ai_1 _17710_ (.A1(_10279_),
    .A2(_01906_),
    .B1(_01797_),
    .Y(_01908_));
 sky130_fd_sc_hd__nand2_1 _17711_ (.A(_01907_),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__nand2_2 _17712_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08318_),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _17713_ (.A(_08405_),
    .B(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__xor2_1 _17714_ (.A(_01909_),
    .B(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__a21bo_1 _17715_ (.A1(_01701_),
    .A2(_01819_),
    .B1_N(_01821_),
    .X(_01913_));
 sky130_fd_sc_hd__and2b_1 _17716_ (.A_N(_01912_),
    .B(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__and2b_1 _17717_ (.A_N(_01913_),
    .B(_01912_),
    .X(_01915_));
 sky130_fd_sc_hd__nor2_1 _17718_ (.A(_01914_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_1 _17719_ (.A(_01905_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__a21oi_1 _17720_ (.A1(_01790_),
    .A2(_01803_),
    .B1(_01801_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _17721_ (.A(_01917_),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__and2_1 _17722_ (.A(_01917_),
    .B(_01918_),
    .X(_01920_));
 sky130_fd_sc_hd__nor2_1 _17723_ (.A(_01919_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__xnor2_1 _17724_ (.A(_01904_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__a21o_1 _17725_ (.A1(_01894_),
    .A2(_01895_),
    .B1(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__nand3_1 _17726_ (.A(_01894_),
    .B(_01895_),
    .C(_01922_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _17727_ (.A(_01923_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__xnor2_1 _17728_ (.A(_01893_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__or2b_1 _17729_ (.A(_09647_),
    .B_N(_01841_),
    .X(_01927_));
 sky130_fd_sc_hd__o21ai_1 _17730_ (.A1(_10289_),
    .A2(_01927_),
    .B1(_01723_),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _17731_ (.A(_09647_),
    .B(_10302_),
    .Y(_01929_));
 sky130_fd_sc_hd__mux2_1 _17732_ (.A0(_01929_),
    .A1(_09647_),
    .S(_01841_),
    .X(_01930_));
 sky130_fd_sc_hd__nand2_1 _17733_ (.A(_01722_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__or2_1 _17734_ (.A(_01722_),
    .B(_01930_),
    .X(_01932_));
 sky130_fd_sc_hd__nand2_2 _17735_ (.A(_01931_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__xnor2_1 _17736_ (.A(_01928_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__xnor2_1 _17737_ (.A(_01734_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__a21boi_1 _17738_ (.A1(_01734_),
    .A2(_01846_),
    .B1_N(_01731_),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _17739_ (.A(_01935_),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__and2_1 _17740_ (.A(_01935_),
    .B(_01936_),
    .X(_01938_));
 sky130_fd_sc_hd__nor2_1 _17741_ (.A(_01937_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__a21o_1 _17742_ (.A1(_01823_),
    .A2(_01833_),
    .B1(_01831_),
    .X(_01940_));
 sky130_fd_sc_hd__nand2_1 _17743_ (.A(_01722_),
    .B(_01842_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor2_1 _17744_ (.A(_10269_),
    .B(_09181_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_1 _17745_ (.A(_10269_),
    .B(_09286_),
    .Y(_01943_));
 sky130_fd_sc_hd__nor2_1 _17746_ (.A(_10386_),
    .B(_09181_),
    .Y(_01944_));
 sky130_fd_sc_hd__nor2_1 _17747_ (.A(_01943_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__a21o_1 _17748_ (.A1(_01819_),
    .A2(_01942_),
    .B1(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__or3_1 _17749_ (.A(_09295_),
    .B(_01818_),
    .C(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__o21ai_1 _17750_ (.A1(_09295_),
    .A2(_01818_),
    .B1(_01946_),
    .Y(_01948_));
 sky130_fd_sc_hd__and2_1 _17751_ (.A(_01947_),
    .B(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__or3_1 _17752_ (.A(_08798_),
    .B(_10289_),
    .C(_01824_),
    .X(_01950_));
 sky130_fd_sc_hd__o21ai_1 _17753_ (.A1(_08798_),
    .A2(_10289_),
    .B1(_01824_),
    .Y(_01951_));
 sky130_fd_sc_hd__nand2_1 _17754_ (.A(_01950_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__or2_1 _17755_ (.A(_09512_),
    .B(_10069_),
    .X(_01953_));
 sky130_fd_sc_hd__xnor2_1 _17756_ (.A(_01952_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__o31a_1 _17757_ (.A1(_08798_),
    .A2(_10069_),
    .A3(_01824_),
    .B1(_01827_),
    .X(_01955_));
 sky130_fd_sc_hd__xor2_1 _17758_ (.A(_01954_),
    .B(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__xnor2_1 _17759_ (.A(_01949_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__a21o_1 _17760_ (.A1(_01941_),
    .A2(_01844_),
    .B1(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__nand3_1 _17761_ (.A(_01941_),
    .B(_01844_),
    .C(_01957_),
    .Y(_01959_));
 sky130_fd_sc_hd__nand2_1 _17762_ (.A(_01958_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__xnor2_1 _17763_ (.A(_01940_),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__xnor2_1 _17764_ (.A(_01939_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__a21oi_1 _17765_ (.A1(_01836_),
    .A2(_01851_),
    .B1(_01849_),
    .Y(_01963_));
 sky130_fd_sc_hd__xor2_1 _17766_ (.A(_01962_),
    .B(_01963_),
    .X(_01964_));
 sky130_fd_sc_hd__nand2_1 _17767_ (.A(_01926_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__or2_1 _17768_ (.A(_01926_),
    .B(_01964_),
    .X(_01966_));
 sky130_fd_sc_hd__nand2_1 _17769_ (.A(_01965_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _17770_ (.A(_01852_),
    .B(_01854_),
    .Y(_01968_));
 sky130_fd_sc_hd__a21oi_1 _17771_ (.A1(_01814_),
    .A2(_01855_),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__xor2_1 _17772_ (.A(_01967_),
    .B(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__xnor2_1 _17773_ (.A(_01892_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__nor2_1 _17774_ (.A(_01856_),
    .B(_01858_),
    .Y(_01972_));
 sky130_fd_sc_hd__a21oi_1 _17775_ (.A1(_01775_),
    .A2(_01859_),
    .B1(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_1 _17776_ (.A(_01971_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__and2_1 _17777_ (.A(_01971_),
    .B(_01973_),
    .X(_01975_));
 sky130_fd_sc_hd__nor2_1 _17778_ (.A(_01974_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__xnor2_1 _17779_ (.A(_01773_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__a21o_2 _17780_ (.A1(_01863_),
    .A2(_01866_),
    .B1(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__and3_2 _17781_ (.A(_01863_),
    .B(_01866_),
    .C(_01977_),
    .X(_01979_));
 sky130_fd_sc_hd__inv_2 _17782_ (.A(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__nand2_1 _17783_ (.A(_01978_),
    .B(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__a21oi_1 _17784_ (.A1(_01870_),
    .A2(_01878_),
    .B1(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__a31o_1 _17785_ (.A1(_01870_),
    .A2(_01878_),
    .A3(_01981_),
    .B1(_08099_),
    .X(_01983_));
 sky130_fd_sc_hd__or2_1 _17786_ (.A(_01982_),
    .B(_01983_),
    .X(_01984_));
 sky130_fd_sc_hd__o21ai_1 _17787_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__mux2_1 _17788_ (.A0(\rbzero.wall_tracer.trackDistX[7] ),
    .A1(_01985_),
    .S(_09826_),
    .X(_01986_));
 sky130_fd_sc_hd__clkbuf_1 _17789_ (.A(_01986_),
    .X(_00546_));
 sky130_fd_sc_hd__or2b_1 _17790_ (.A(_01925_),
    .B_N(_01893_),
    .X(_01987_));
 sky130_fd_sc_hd__o2bb2a_1 _17791_ (.A1_N(_01902_),
    .A2_N(_01903_),
    .B1(_01900_),
    .B2(_01901_),
    .X(_01988_));
 sky130_fd_sc_hd__a21o_1 _17792_ (.A1(_01923_),
    .A2(_01987_),
    .B1(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__nand3_1 _17793_ (.A(_01923_),
    .B(_01987_),
    .C(_01988_),
    .Y(_01990_));
 sky130_fd_sc_hd__and2_1 _17794_ (.A(_01989_),
    .B(_01990_),
    .X(_01991_));
 sky130_fd_sc_hd__a21bo_1 _17795_ (.A1(_01734_),
    .A2(_01934_),
    .B1_N(_01731_),
    .X(_01992_));
 sky130_fd_sc_hd__and2_1 _17796_ (.A(_01723_),
    .B(_01927_),
    .X(_01993_));
 sky130_fd_sc_hd__xor2_2 _17797_ (.A(_01933_),
    .B(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__xor2_1 _17798_ (.A(_01734_),
    .B(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__and2_1 _17799_ (.A(_01992_),
    .B(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__nor2_1 _17800_ (.A(_01992_),
    .B(_01995_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _17801_ (.A(_01996_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__nor2_1 _17802_ (.A(_01954_),
    .B(_01955_),
    .Y(_01999_));
 sky130_fd_sc_hd__a21o_1 _17803_ (.A1(_01949_),
    .A2(_01956_),
    .B1(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__a21bo_1 _17804_ (.A1(_01928_),
    .A2(_01932_),
    .B1_N(_01931_),
    .X(_02001_));
 sky130_fd_sc_hd__nor2_1 _17805_ (.A(_08127_),
    .B(_09409_),
    .Y(_02002_));
 sky130_fd_sc_hd__xnor2_1 _17806_ (.A(_01942_),
    .B(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__or3_1 _17807_ (.A(_01818_),
    .B(_09286_),
    .C(_02003_),
    .X(_02004_));
 sky130_fd_sc_hd__o21ai_1 _17808_ (.A1(_01818_),
    .A2(_09286_),
    .B1(_02003_),
    .Y(_02005_));
 sky130_fd_sc_hd__and2_1 _17809_ (.A(_02004_),
    .B(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__and3b_1 _17810_ (.A_N(_08798_),
    .B(_08513_),
    .C(_01839_),
    .X(_02007_));
 sky130_fd_sc_hd__o22a_1 _17811_ (.A1(_08798_),
    .A2(_10302_),
    .B1(_10289_),
    .B2(_09506_),
    .X(_02008_));
 sky130_fd_sc_hd__a21oi_1 _17812_ (.A1(_01724_),
    .A2(_02007_),
    .B1(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _17813_ (.A(_09512_),
    .B(_09663_),
    .Y(_02010_));
 sky130_fd_sc_hd__xnor2_1 _17814_ (.A(_02009_),
    .B(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__o21a_1 _17815_ (.A1(_01952_),
    .A2(_01953_),
    .B1(_01950_),
    .X(_02012_));
 sky130_fd_sc_hd__xor2_1 _17816_ (.A(_02011_),
    .B(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__nand2_1 _17817_ (.A(_02006_),
    .B(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__or2_1 _17818_ (.A(_02006_),
    .B(_02013_),
    .X(_02015_));
 sky130_fd_sc_hd__and2_1 _17819_ (.A(_02014_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__xnor2_1 _17820_ (.A(_02001_),
    .B(_02016_),
    .Y(_02017_));
 sky130_fd_sc_hd__xnor2_1 _17821_ (.A(_02000_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__xnor2_1 _17822_ (.A(_01998_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__a21oi_1 _17823_ (.A1(_01939_),
    .A2(_01961_),
    .B1(_01937_),
    .Y(_02020_));
 sky130_fd_sc_hd__xor2_1 _17824_ (.A(_02019_),
    .B(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__a21o_1 _17825_ (.A1(_01904_),
    .A2(_01921_),
    .B1(_01919_),
    .X(_02022_));
 sky130_fd_sc_hd__or2b_1 _17826_ (.A(_01960_),
    .B_N(_01940_),
    .X(_02023_));
 sky130_fd_sc_hd__or2_1 _17827_ (.A(_08479_),
    .B(_09228_),
    .X(_02024_));
 sky130_fd_sc_hd__or3_1 _17828_ (.A(_10268_),
    .B(_09342_),
    .C(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__o21ai_1 _17829_ (.A1(_10268_),
    .A2(_09342_),
    .B1(_02024_),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(_02025_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _17831_ (.A(_09911_),
    .B(_09605_),
    .Y(_02028_));
 sky130_fd_sc_hd__xor2_1 _17832_ (.A(_02027_),
    .B(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _17833_ (.A(_01896_),
    .B(_01897_),
    .Y(_02030_));
 sky130_fd_sc_hd__o31a_1 _17834_ (.A1(_10038_),
    .A2(_09605_),
    .A3(_01898_),
    .B1(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__xor2_1 _17835_ (.A(_02029_),
    .B(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__and2_1 _17836_ (.A(_10038_),
    .B(_09869_),
    .X(_02033_));
 sky130_fd_sc_hd__xor2_1 _17837_ (.A(_02032_),
    .B(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__o31ai_2 _17838_ (.A1(_08405_),
    .A2(_01910_),
    .A3(_01909_),
    .B1(_01907_),
    .Y(_02035_));
 sky130_fd_sc_hd__a21bo_1 _17839_ (.A1(_01943_),
    .A2(_01944_),
    .B1_N(_01947_),
    .X(_02036_));
 sky130_fd_sc_hd__or2_1 _17840_ (.A(_09295_),
    .B(_01794_),
    .X(_02037_));
 sky130_fd_sc_hd__or3_1 _17841_ (.A(_10279_),
    .B(_01906_),
    .C(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__o22ai_1 _17842_ (.A1(_09295_),
    .A2(_01906_),
    .B1(_01794_),
    .B2(_10279_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2_1 _17843_ (.A(_02038_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _17844_ (.A(_10387_),
    .B(_01910_),
    .Y(_02041_));
 sky130_fd_sc_hd__xor2_1 _17845_ (.A(_02040_),
    .B(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__xnor2_1 _17846_ (.A(_02036_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__xnor2_1 _17847_ (.A(_02035_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__a21oi_1 _17848_ (.A1(_01905_),
    .A2(_01916_),
    .B1(_01914_),
    .Y(_02045_));
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(_02044_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__and2_1 _17850_ (.A(_02044_),
    .B(_02045_),
    .X(_02047_));
 sky130_fd_sc_hd__nor2_1 _17851_ (.A(_02046_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__xnor2_1 _17852_ (.A(_02034_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__a21o_1 _17853_ (.A1(_01958_),
    .A2(_02023_),
    .B1(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__nand3_1 _17854_ (.A(_01958_),
    .B(_02023_),
    .C(_02049_),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _17855_ (.A(_02050_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__xnor2_1 _17856_ (.A(_02022_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_1 _17857_ (.A(_02021_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__or2_1 _17858_ (.A(_02021_),
    .B(_02053_),
    .X(_02055_));
 sky130_fd_sc_hd__nand2_1 _17859_ (.A(_02054_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__o21a_1 _17860_ (.A1(_01962_),
    .A2(_01963_),
    .B1(_01965_),
    .X(_02057_));
 sky130_fd_sc_hd__xor2_1 _17861_ (.A(_02056_),
    .B(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__nand2_1 _17862_ (.A(_01991_),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__or2_1 _17863_ (.A(_01991_),
    .B(_02058_),
    .X(_02060_));
 sky130_fd_sc_hd__nand2_1 _17864_ (.A(_02059_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__nor2_1 _17865_ (.A(_01967_),
    .B(_01969_),
    .Y(_02062_));
 sky130_fd_sc_hd__a21oi_2 _17866_ (.A1(_01892_),
    .A2(_01970_),
    .B1(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__xor2_1 _17867_ (.A(_02061_),
    .B(_02063_),
    .X(_02064_));
 sky130_fd_sc_hd__xnor2_1 _17868_ (.A(_01890_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__a21oi_2 _17869_ (.A1(_01773_),
    .A2(_01976_),
    .B1(_01974_),
    .Y(_02066_));
 sky130_fd_sc_hd__or2_1 _17870_ (.A(_02065_),
    .B(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__nand2_1 _17871_ (.A(_02065_),
    .B(_02066_),
    .Y(_02068_));
 sky130_fd_sc_hd__and2_1 _17872_ (.A(_02067_),
    .B(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__inv_2 _17873_ (.A(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__a311o_1 _17874_ (.A1(_01870_),
    .A2(_01878_),
    .A3(_01978_),
    .B1(_01979_),
    .C1(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__a31o_1 _17875_ (.A1(_01870_),
    .A2(_01878_),
    .A3(_01978_),
    .B1(_01979_),
    .X(_02072_));
 sky130_fd_sc_hd__a21oi_1 _17876_ (.A1(_02070_),
    .A2(_02072_),
    .B1(_08101_),
    .Y(_02073_));
 sky130_fd_sc_hd__nand2_1 _17877_ (.A(_02071_),
    .B(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__or2_1 _17878_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .X(_02075_));
 sky130_fd_sc_hd__nand2_1 _17879_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_1 _17880_ (.A(_02075_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__o21a_1 _17881_ (.A1(_01882_),
    .A2(_01885_),
    .B1(_01883_),
    .X(_02078_));
 sky130_fd_sc_hd__or2_1 _17882_ (.A(_02077_),
    .B(_02078_),
    .X(_02079_));
 sky130_fd_sc_hd__a21oi_1 _17883_ (.A1(_02077_),
    .A2(_02078_),
    .B1(_09789_),
    .Y(_02080_));
 sky130_fd_sc_hd__a21oi_1 _17884_ (.A1(_02079_),
    .A2(_02080_),
    .B1(_09763_),
    .Y(_02081_));
 sky130_fd_sc_hd__o2bb2a_1 _17885_ (.A1_N(_02074_),
    .A2_N(_02081_),
    .B1(\rbzero.wall_tracer.trackDistX[8] ),
    .B2(_09805_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _17886_ (.A(_02061_),
    .B(_02063_),
    .X(_02082_));
 sky130_fd_sc_hd__nand2_1 _17887_ (.A(_01890_),
    .B(_02064_),
    .Y(_02083_));
 sky130_fd_sc_hd__a21o_1 _17888_ (.A1(_01998_),
    .A2(_02018_),
    .B1(_01996_),
    .X(_02084_));
 sky130_fd_sc_hd__o21ai_1 _17889_ (.A1(_02011_),
    .A2(_02012_),
    .B1(_02014_),
    .Y(_02085_));
 sky130_fd_sc_hd__o21ai_2 _17890_ (.A1(_01933_),
    .A2(_01993_),
    .B1(_01931_),
    .Y(_02086_));
 sky130_fd_sc_hd__or2_1 _17891_ (.A(_06163_),
    .B(_09406_),
    .X(_02087_));
 sky130_fd_sc_hd__nor2_1 _17892_ (.A(_10269_),
    .B(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__o22a_1 _17893_ (.A1(_08286_),
    .A2(_09409_),
    .B1(_02087_),
    .B2(_10386_),
    .X(_02089_));
 sky130_fd_sc_hd__a21oi_1 _17894_ (.A1(_02002_),
    .A2(_02088_),
    .B1(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _17895_ (.A(_01818_),
    .B(_09181_),
    .Y(_02091_));
 sky130_fd_sc_hd__xnor2_1 _17896_ (.A(_02090_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__a22o_1 _17897_ (.A1(_01724_),
    .A2(_02007_),
    .B1(_02009_),
    .B2(_02010_),
    .X(_02093_));
 sky130_fd_sc_hd__nand2_1 _17898_ (.A(_08798_),
    .B(_09506_),
    .Y(_02094_));
 sky130_fd_sc_hd__or3b_1 _17899_ (.A(_10302_),
    .B(_02007_),
    .C_N(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__or2_1 _17900_ (.A(_09512_),
    .B(_10289_),
    .X(_02096_));
 sky130_fd_sc_hd__xor2_1 _17901_ (.A(_02095_),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__and2_1 _17902_ (.A(_02093_),
    .B(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__nor2_1 _17903_ (.A(_02093_),
    .B(_02097_),
    .Y(_02099_));
 sky130_fd_sc_hd__nor2_1 _17904_ (.A(_02098_),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__xnor2_1 _17905_ (.A(_02092_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__xor2_1 _17906_ (.A(_02086_),
    .B(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__nand2_1 _17907_ (.A(_02085_),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__or2_1 _17908_ (.A(_02085_),
    .B(_02102_),
    .X(_02104_));
 sky130_fd_sc_hd__nand2_1 _17909_ (.A(_02103_),
    .B(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__mux2_1 _17910_ (.A0(_01732_),
    .A1(_01731_),
    .S(_01994_),
    .X(_02106_));
 sky130_fd_sc_hd__xnor2_1 _17911_ (.A(_02105_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__xnor2_1 _17912_ (.A(_02084_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__a21o_1 _17913_ (.A1(_02034_),
    .A2(_02048_),
    .B1(_02046_),
    .X(_02109_));
 sky130_fd_sc_hd__or2b_1 _17914_ (.A(_02017_),
    .B_N(_02000_),
    .X(_02110_));
 sky130_fd_sc_hd__a21bo_1 _17915_ (.A1(_02001_),
    .A2(_02016_),
    .B1_N(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__or2_1 _17916_ (.A(_08479_),
    .B(_09342_),
    .X(_02112_));
 sky130_fd_sc_hd__nand2_1 _17917_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_10389_),
    .Y(_02113_));
 sky130_fd_sc_hd__xnor2_1 _17918_ (.A(_02112_),
    .B(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__or3_1 _17919_ (.A(_10268_),
    .B(_09605_),
    .C(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__o21ai_1 _17920_ (.A1(_10268_),
    .A2(_09605_),
    .B1(_02114_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2_1 _17921_ (.A(_02115_),
    .B(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__o31a_1 _17922_ (.A1(_09911_),
    .A2(_09605_),
    .A3(_02027_),
    .B1(_02025_),
    .X(_02118_));
 sky130_fd_sc_hd__xnor2_1 _17923_ (.A(_02117_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _17924_ (.A(_09911_),
    .B(_09869_),
    .Y(_02120_));
 sky130_fd_sc_hd__xnor2_1 _17925_ (.A(_02119_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__a21bo_1 _17926_ (.A1(_02039_),
    .A2(_02041_),
    .B1_N(_02038_),
    .X(_02122_));
 sky130_fd_sc_hd__a21bo_1 _17927_ (.A1(_01942_),
    .A2(_02002_),
    .B1_N(_02004_),
    .X(_02123_));
 sky130_fd_sc_hd__or3_1 _17928_ (.A(_01906_),
    .B(_09286_),
    .C(_02037_),
    .X(_02124_));
 sky130_fd_sc_hd__o21ai_1 _17929_ (.A1(_01906_),
    .A2(_09286_),
    .B1(_02037_),
    .Y(_02125_));
 sky130_fd_sc_hd__and2_1 _17930_ (.A(_02124_),
    .B(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__nor2_1 _17931_ (.A(_10279_),
    .B(_01910_),
    .Y(_02127_));
 sky130_fd_sc_hd__xor2_1 _17932_ (.A(_02126_),
    .B(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__nand2_1 _17933_ (.A(_02123_),
    .B(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__or2_1 _17934_ (.A(_02123_),
    .B(_02128_),
    .X(_02130_));
 sky130_fd_sc_hd__and2_1 _17935_ (.A(_02129_),
    .B(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__xnor2_1 _17936_ (.A(_02122_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__and2b_1 _17937_ (.A_N(_02042_),
    .B(_02036_),
    .X(_02133_));
 sky130_fd_sc_hd__a21oi_1 _17938_ (.A1(_02035_),
    .A2(_02043_),
    .B1(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__xor2_1 _17939_ (.A(_02132_),
    .B(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__xnor2_1 _17940_ (.A(_02121_),
    .B(_02135_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _17941_ (.A(_02111_),
    .B(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__or2_1 _17942_ (.A(_02111_),
    .B(_02136_),
    .X(_02138_));
 sky130_fd_sc_hd__and2_1 _17943_ (.A(_02137_),
    .B(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__xor2_1 _17944_ (.A(_02109_),
    .B(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__xor2_1 _17945_ (.A(_02108_),
    .B(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__o21a_1 _17946_ (.A1(_02019_),
    .A2(_02020_),
    .B1(_02054_),
    .X(_02142_));
 sky130_fd_sc_hd__xor2_1 _17947_ (.A(_02141_),
    .B(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__or2b_1 _17948_ (.A(_02052_),
    .B_N(_02022_),
    .X(_02144_));
 sky130_fd_sc_hd__o2bb2a_1 _17949_ (.A1_N(_02032_),
    .A2_N(_02033_),
    .B1(_02029_),
    .B2(_02031_),
    .X(_02145_));
 sky130_fd_sc_hd__a21o_1 _17950_ (.A1(_02050_),
    .A2(_02144_),
    .B1(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__nand3_1 _17951_ (.A(_02050_),
    .B(_02144_),
    .C(_02145_),
    .Y(_02147_));
 sky130_fd_sc_hd__and2_1 _17952_ (.A(_02146_),
    .B(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__nand2_1 _17953_ (.A(_02143_),
    .B(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__or2_1 _17954_ (.A(_02143_),
    .B(_02148_),
    .X(_02150_));
 sky130_fd_sc_hd__nand2_1 _17955_ (.A(_02149_),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__o21a_1 _17956_ (.A1(_02056_),
    .A2(_02057_),
    .B1(_02059_),
    .X(_02152_));
 sky130_fd_sc_hd__xor2_1 _17957_ (.A(_02151_),
    .B(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__xor2_1 _17958_ (.A(_01989_),
    .B(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__a21o_1 _17959_ (.A1(_02082_),
    .A2(_02083_),
    .B1(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__and3_1 _17960_ (.A(_02082_),
    .B(_02083_),
    .C(_02154_),
    .X(_02156_));
 sky130_fd_sc_hd__inv_2 _17961_ (.A(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_1 _17962_ (.A(_02155_),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21oi_1 _17963_ (.A1(_02067_),
    .A2(_02071_),
    .B1(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__a31o_1 _17964_ (.A1(_02067_),
    .A2(_02071_),
    .A3(_02158_),
    .B1(_08100_),
    .X(_02160_));
 sky130_fd_sc_hd__or2_1 _17965_ (.A(_02159_),
    .B(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__and2_1 _17966_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_02162_));
 sky130_fd_sc_hd__nor2_1 _17967_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_02163_));
 sky130_fd_sc_hd__nor2_1 _17968_ (.A(_02162_),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__nand2_1 _17969_ (.A(_02076_),
    .B(_02078_),
    .Y(_02165_));
 sky130_fd_sc_hd__and2_1 _17970_ (.A(_02075_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__xnor2_1 _17971_ (.A(_02164_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__o21a_1 _17972_ (.A1(_10107_),
    .A2(_02167_),
    .B1(_09805_),
    .X(_02168_));
 sky130_fd_sc_hd__o2bb2a_1 _17973_ (.A1_N(_02161_),
    .A2_N(_02168_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_09805_),
    .X(_00548_));
 sky130_fd_sc_hd__a21o_1 _17974_ (.A1(_02067_),
    .A2(_02155_),
    .B1(_02156_),
    .X(_02169_));
 sky130_fd_sc_hd__or2b_1 _17975_ (.A(_01989_),
    .B_N(_02153_),
    .X(_02170_));
 sky130_fd_sc_hd__o21a_1 _17976_ (.A1(_02151_),
    .A2(_02152_),
    .B1(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__o22a_1 _17977_ (.A1(_02117_),
    .A2(_02118_),
    .B1(_02119_),
    .B2(_02120_),
    .X(_02172_));
 sky130_fd_sc_hd__o21ai_1 _17978_ (.A1(_02141_),
    .A2(_02142_),
    .B1(_02149_),
    .Y(_02173_));
 sky130_fd_sc_hd__or2_1 _17979_ (.A(_01732_),
    .B(_01994_),
    .X(_02174_));
 sky130_fd_sc_hd__a32o_1 _17980_ (.A1(_10075_),
    .A2(_10419_),
    .A3(_01994_),
    .B1(_02174_),
    .B2(_02105_),
    .X(_02175_));
 sky130_fd_sc_hd__xnor2_1 _17981_ (.A(_02086_),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _17982_ (.A(_09512_),
    .B(_10302_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _17983_ (.A(_10386_),
    .B(_09951_),
    .Y(_02178_));
 sky130_fd_sc_hd__xor2_1 _17984_ (.A(_02088_),
    .B(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__xnor2_1 _17985_ (.A(_02177_),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _17986_ (.A(_01906_),
    .B(_09181_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _17987_ (.A(_02002_),
    .B(_02088_),
    .Y(_02182_));
 sky130_fd_sc_hd__o31a_1 _17988_ (.A1(_01818_),
    .A2(_09181_),
    .A3(_02089_),
    .B1(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__nand2_1 _17989_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_10389_),
    .Y(_02184_));
 sky130_fd_sc_hd__o21ai_1 _17990_ (.A1(_02024_),
    .A2(_02184_),
    .B1(_02115_),
    .Y(_02185_));
 sky130_fd_sc_hd__or2_1 _17991_ (.A(_08479_),
    .B(_09605_),
    .X(_02186_));
 sky130_fd_sc_hd__or2_1 _17992_ (.A(_08435_),
    .B(_09228_),
    .X(_02187_));
 sky130_fd_sc_hd__xnor2_1 _17993_ (.A(_02184_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__xnor2_1 _17994_ (.A(_02186_),
    .B(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__xnor2_1 _17995_ (.A(_02185_),
    .B(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__a21boi_1 _17996_ (.A1(_02126_),
    .A2(_02127_),
    .B1_N(_02124_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _17997_ (.A(_09295_),
    .B(_01910_),
    .Y(_02192_));
 sky130_fd_sc_hd__xor2_1 _17998_ (.A(_02191_),
    .B(_02192_),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_1 _17999_ (.A(_02190_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__xnor2_1 _18000_ (.A(_02183_),
    .B(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__xnor2_1 _18001_ (.A(_02181_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _18002_ (.A(_09286_),
    .B(_01794_),
    .Y(_02197_));
 sky130_fd_sc_hd__a21bo_1 _18003_ (.A1(_02122_),
    .A2(_02131_),
    .B1_N(_02129_),
    .X(_02198_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_02197_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__or2b_1 _18005_ (.A(_02121_),
    .B_N(_02135_),
    .X(_02200_));
 sky130_fd_sc_hd__o21a_1 _18006_ (.A1(_02132_),
    .A2(_02134_),
    .B1(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__xnor2_1 _18007_ (.A(_02199_),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__xnor2_1 _18008_ (.A(_02196_),
    .B(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__xnor2_1 _18009_ (.A(_02180_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__xnor2_1 _18010_ (.A(_02176_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__a21boi_1 _18011_ (.A1(_02086_),
    .A2(_02101_),
    .B1_N(_02103_),
    .Y(_02206_));
 sky130_fd_sc_hd__o21ba_1 _18012_ (.A1(_02092_),
    .A2(_02099_),
    .B1_N(_02098_),
    .X(_02207_));
 sky130_fd_sc_hd__nor2_1 _18013_ (.A(_09132_),
    .B(_09409_),
    .Y(_02208_));
 sky130_fd_sc_hd__xnor2_1 _18014_ (.A(_02207_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_1 _18015_ (.A(_10268_),
    .B(_09869_),
    .Y(_02210_));
 sky130_fd_sc_hd__xnor2_1 _18016_ (.A(_02209_),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__xnor2_1 _18017_ (.A(_02206_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__xnor2_1 _18018_ (.A(_02146_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__xnor2_1 _18019_ (.A(_02205_),
    .B(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__and2b_1 _18020_ (.A_N(_02108_),
    .B(_02140_),
    .X(_02215_));
 sky130_fd_sc_hd__a21o_1 _18021_ (.A1(_02084_),
    .A2(_02107_),
    .B1(_02215_),
    .X(_02216_));
 sky130_fd_sc_hd__a31o_1 _18022_ (.A1(_01839_),
    .A2(_02094_),
    .A3(_02096_),
    .B1(_02007_),
    .X(_02217_));
 sky130_fd_sc_hd__a21bo_1 _18023_ (.A1(_02109_),
    .A2(_02139_),
    .B1_N(_02137_),
    .X(_02218_));
 sky130_fd_sc_hd__xnor2_1 _18024_ (.A(_02217_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__xnor2_1 _18025_ (.A(_02216_),
    .B(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__xnor2_1 _18026_ (.A(_02214_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__xnor2_1 _18027_ (.A(_02173_),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__xnor2_1 _18028_ (.A(_02172_),
    .B(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__xor2_1 _18029_ (.A(_02171_),
    .B(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__o211a_1 _18030_ (.A1(_02071_),
    .A2(_02158_),
    .B1(_02169_),
    .C1(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__a311o_1 _18031_ (.A1(_02067_),
    .A2(_02071_),
    .A3(_02155_),
    .B1(_02156_),
    .C1(_02224_),
    .X(_02226_));
 sky130_fd_sc_hd__or3b_1 _18032_ (.A(_08100_),
    .B(_02225_),
    .C_N(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__a31o_1 _18033_ (.A1(_02075_),
    .A2(_02164_),
    .A3(_02165_),
    .B1(_02162_),
    .X(_02228_));
 sky130_fd_sc_hd__xnor2_1 _18034_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_02229_));
 sky130_fd_sc_hd__xnor2_1 _18035_ (.A(_02228_),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__a21oi_1 _18036_ (.A1(_08101_),
    .A2(_02230_),
    .B1(_09761_),
    .Y(_02231_));
 sky130_fd_sc_hd__o2bb2a_1 _18037_ (.A1_N(_02227_),
    .A2_N(_02231_),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_09805_),
    .X(_00549_));
 sky130_fd_sc_hd__and2_1 _18038_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_02232_));
 sky130_fd_sc_hd__nor2_1 _18039_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_02233_));
 sky130_fd_sc_hd__o21a_1 _18040_ (.A1(_06156_),
    .A2(_08406_),
    .B1(_06254_),
    .X(_02234_));
 sky130_fd_sc_hd__buf_4 _18041_ (.A(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__o31a_1 _18042_ (.A1(_10338_),
    .A2(_02232_),
    .A3(_02233_),
    .B1(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__buf_4 _18043_ (.A(_02234_),
    .X(_02237_));
 sky130_fd_sc_hd__clkbuf_4 _18044_ (.A(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__o2bb2a_1 _18045_ (.A1_N(_09785_),
    .A2_N(_02236_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-11] ),
    .X(_00550_));
 sky130_fd_sc_hd__nand2_1 _18046_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_02239_));
 sky130_fd_sc_hd__or2_1 _18047_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_02240_));
 sky130_fd_sc_hd__and4_1 _18048_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .C(_02239_),
    .D(_02240_),
    .X(_02241_));
 sky130_fd_sc_hd__a22oi_1 _18049_ (.A1(\rbzero.wall_tracer.trackDistY[-11] ),
    .A2(\rbzero.wall_tracer.stepDistY[-11] ),
    .B1(_02239_),
    .B2(_02240_),
    .Y(_02242_));
 sky130_fd_sc_hd__o31a_1 _18050_ (.A1(_10338_),
    .A2(_02241_),
    .A3(_02242_),
    .B1(_02235_),
    .X(_02243_));
 sky130_fd_sc_hd__o2bb2a_1 _18051_ (.A1_N(_09796_),
    .A2_N(_02243_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(_00551_));
 sky130_fd_sc_hd__a21oi_1 _18052_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(\rbzero.wall_tracer.stepDistY[-10] ),
    .B1(_02241_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_1 _18053_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_02245_));
 sky130_fd_sc_hd__and2_1 _18054_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_02246_));
 sky130_fd_sc_hd__nor3_1 _18055_ (.A(_02244_),
    .B(_02245_),
    .C(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__o21a_1 _18056_ (.A1(_02245_),
    .A2(_02246_),
    .B1(_02244_),
    .X(_02248_));
 sky130_fd_sc_hd__o31a_1 _18057_ (.A1(_10338_),
    .A2(_02247_),
    .A3(_02248_),
    .B1(_02235_),
    .X(_02249_));
 sky130_fd_sc_hd__o2bb2a_1 _18058_ (.A1_N(_09803_),
    .A2_N(_02249_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(_00552_));
 sky130_fd_sc_hd__buf_4 _18059_ (.A(_02234_),
    .X(_02250_));
 sky130_fd_sc_hd__or2_1 _18060_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_02251_));
 sky130_fd_sc_hd__nand2_1 _18061_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .Y(_02252_));
 sky130_fd_sc_hd__o21bai_1 _18062_ (.A1(_02244_),
    .A2(_02245_),
    .B1_N(_02246_),
    .Y(_02253_));
 sky130_fd_sc_hd__and3_1 _18063_ (.A(_02251_),
    .B(_02252_),
    .C(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__a21oi_1 _18064_ (.A1(_02251_),
    .A2(_02252_),
    .B1(_02253_),
    .Y(_02255_));
 sky130_fd_sc_hd__o31ai_1 _18065_ (.A1(_10107_),
    .A2(_02254_),
    .A3(_02255_),
    .B1(_02250_),
    .Y(_02256_));
 sky130_fd_sc_hd__o22a_1 _18066_ (.A1(\rbzero.wall_tracer.trackDistY[-8] ),
    .A2(_02250_),
    .B1(_02256_),
    .B2(_09811_),
    .X(_00553_));
 sky130_fd_sc_hd__nor2_1 _18067_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_1 _18068_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02258_));
 sky130_fd_sc_hd__or2b_1 _18069_ (.A(_02257_),
    .B_N(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__a21boi_1 _18070_ (.A1(_02251_),
    .A2(_02253_),
    .B1_N(_02252_),
    .Y(_02260_));
 sky130_fd_sc_hd__xnor2_1 _18071_ (.A(_02259_),
    .B(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__o21a_1 _18072_ (.A1(_10107_),
    .A2(_02261_),
    .B1(_02250_),
    .X(_02262_));
 sky130_fd_sc_hd__o2bb2a_1 _18073_ (.A1_N(_09818_),
    .A2_N(_02262_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-7] ),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _18074_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_02263_));
 sky130_fd_sc_hd__nand2_1 _18075_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .Y(_02264_));
 sky130_fd_sc_hd__o21ai_1 _18076_ (.A1(_02257_),
    .A2(_02260_),
    .B1(_02258_),
    .Y(_02265_));
 sky130_fd_sc_hd__and3_1 _18077_ (.A(_02263_),
    .B(_02264_),
    .C(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__a21oi_1 _18078_ (.A1(_02263_),
    .A2(_02264_),
    .B1(_02265_),
    .Y(_02267_));
 sky130_fd_sc_hd__o31a_1 _18079_ (.A1(_10338_),
    .A2(_02266_),
    .A3(_02267_),
    .B1(_02235_),
    .X(_02268_));
 sky130_fd_sc_hd__o2bb2a_1 _18080_ (.A1_N(_09827_),
    .A2_N(_02268_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(_00555_));
 sky130_fd_sc_hd__nor2_1 _18081_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02270_));
 sky130_fd_sc_hd__or2b_1 _18083_ (.A(_02269_),
    .B_N(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__a21boi_1 _18084_ (.A1(_02263_),
    .A2(_02265_),
    .B1_N(_02264_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _18085_ (.A(_02271_),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__a21o_1 _18086_ (.A1(_02271_),
    .A2(_02272_),
    .B1(_06102_),
    .X(_02274_));
 sky130_fd_sc_hd__o21ai_1 _18087_ (.A1(_02273_),
    .A2(_02274_),
    .B1(_09835_),
    .Y(_02275_));
 sky130_fd_sc_hd__mux2_1 _18088_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(_02275_),
    .S(_02237_),
    .X(_02276_));
 sky130_fd_sc_hd__clkbuf_1 _18089_ (.A(_02276_),
    .X(_00556_));
 sky130_fd_sc_hd__or2_1 _18090_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(_02277_));
 sky130_fd_sc_hd__nand2_1 _18091_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02278_));
 sky130_fd_sc_hd__o21ai_1 _18092_ (.A1(_02269_),
    .A2(_02272_),
    .B1(_02270_),
    .Y(_02279_));
 sky130_fd_sc_hd__and3_1 _18093_ (.A(_02277_),
    .B(_02278_),
    .C(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__a21oi_1 _18094_ (.A1(_02277_),
    .A2(_02278_),
    .B1(_02279_),
    .Y(_02281_));
 sky130_fd_sc_hd__o31a_1 _18095_ (.A1(_10338_),
    .A2(_02280_),
    .A3(_02281_),
    .B1(_02235_),
    .X(_02282_));
 sky130_fd_sc_hd__o2bb2a_1 _18096_ (.A1_N(_09842_),
    .A2_N(_02282_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-4] ),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _18097_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _18098_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02284_));
 sky130_fd_sc_hd__or2b_1 _18099_ (.A(_02283_),
    .B_N(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__a21boi_1 _18100_ (.A1(_02277_),
    .A2(_02279_),
    .B1_N(_02278_),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _18101_ (.A(_02285_),
    .B(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__o21a_1 _18102_ (.A1(_10107_),
    .A2(_02287_),
    .B1(_02250_),
    .X(_02288_));
 sky130_fd_sc_hd__o2bb2a_1 _18103_ (.A1_N(_09849_),
    .A2_N(_02288_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-3] ),
    .X(_00558_));
 sky130_fd_sc_hd__or2_1 _18104_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_02289_));
 sky130_fd_sc_hd__nand2_1 _18105_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02290_));
 sky130_fd_sc_hd__o21ai_1 _18106_ (.A1(_02283_),
    .A2(_02286_),
    .B1(_02284_),
    .Y(_02291_));
 sky130_fd_sc_hd__a21oi_1 _18107_ (.A1(_02289_),
    .A2(_02290_),
    .B1(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__a31o_1 _18108_ (.A1(_02289_),
    .A2(_02290_),
    .A3(_02291_),
    .B1(_09824_),
    .X(_02293_));
 sky130_fd_sc_hd__o21a_1 _18109_ (.A1(_02292_),
    .A2(_02293_),
    .B1(_02235_),
    .X(_02294_));
 sky130_fd_sc_hd__o2bb2a_1 _18110_ (.A1_N(_09856_),
    .A2_N(_02294_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_00559_));
 sky130_fd_sc_hd__nor2_1 _18111_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_02295_));
 sky130_fd_sc_hd__and2_1 _18112_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .X(_02296_));
 sky130_fd_sc_hd__or2_1 _18113_ (.A(_02295_),
    .B(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__a21boi_1 _18114_ (.A1(_02289_),
    .A2(_02291_),
    .B1_N(_02290_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _18115_ (.A(_02297_),
    .B(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__a21o_1 _18116_ (.A1(_02297_),
    .A2(_02298_),
    .B1(_06102_),
    .X(_02300_));
 sky130_fd_sc_hd__o21ai_1 _18117_ (.A1(_02299_),
    .A2(_02300_),
    .B1(_09863_),
    .Y(_02301_));
 sky130_fd_sc_hd__mux2_1 _18118_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(_02301_),
    .S(_02237_),
    .X(_02302_));
 sky130_fd_sc_hd__clkbuf_1 _18119_ (.A(_02302_),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _18120_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .X(_02303_));
 sky130_fd_sc_hd__nand2_1 _18121_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_02304_));
 sky130_fd_sc_hd__o211a_1 _18122_ (.A1(_02296_),
    .A2(_02299_),
    .B1(_02303_),
    .C1(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__a211oi_1 _18123_ (.A1(_02303_),
    .A2(_02304_),
    .B1(_02296_),
    .C1(_02299_),
    .Y(_02306_));
 sky130_fd_sc_hd__o31a_1 _18124_ (.A1(_10338_),
    .A2(_02305_),
    .A3(_02306_),
    .B1(_02237_),
    .X(_02307_));
 sky130_fd_sc_hd__o2bb2a_1 _18125_ (.A1_N(_09990_),
    .A2_N(_02307_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[0] ),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_1 _18126_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_02308_));
 sky130_fd_sc_hd__or2_1 _18127_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__a21o_1 _18128_ (.A1(\rbzero.wall_tracer.trackDistY[0] ),
    .A2(\rbzero.wall_tracer.stepDistY[0] ),
    .B1(_02305_),
    .X(_02310_));
 sky130_fd_sc_hd__and3_1 _18129_ (.A(_02308_),
    .B(_02309_),
    .C(_02310_),
    .X(_02311_));
 sky130_fd_sc_hd__a21o_1 _18130_ (.A1(_02308_),
    .A2(_02309_),
    .B1(_02310_),
    .X(_02312_));
 sky130_fd_sc_hd__or3b_1 _18131_ (.A(_06101_),
    .B(_02311_),
    .C_N(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__nand2_1 _18132_ (.A(_10106_),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__mux2_1 _18133_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(_02314_),
    .S(_02237_),
    .X(_02315_));
 sky130_fd_sc_hd__clkbuf_1 _18134_ (.A(_02315_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _18135_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_02316_));
 sky130_fd_sc_hd__or2_1 _18136_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_02317_));
 sky130_fd_sc_hd__inv_2 _18137_ (.A(_02308_),
    .Y(_02318_));
 sky130_fd_sc_hd__a211o_1 _18138_ (.A1(_02316_),
    .A2(_02317_),
    .B1(_02318_),
    .C1(_02311_),
    .X(_02319_));
 sky130_fd_sc_hd__o211ai_2 _18139_ (.A1(_02318_),
    .A2(_02311_),
    .B1(_02316_),
    .C1(_02317_),
    .Y(_02320_));
 sky130_fd_sc_hd__a31o_1 _18140_ (.A1(_08100_),
    .A2(_02319_),
    .A3(_02320_),
    .B1(_10219_),
    .X(_02321_));
 sky130_fd_sc_hd__mux2_1 _18141_ (.A0(\rbzero.wall_tracer.trackDistY[2] ),
    .A1(_02321_),
    .S(_02237_),
    .X(_02322_));
 sky130_fd_sc_hd__clkbuf_1 _18142_ (.A(_02322_),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _18143_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_02323_));
 sky130_fd_sc_hd__nor2_1 _18144_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_02324_));
 sky130_fd_sc_hd__o211a_1 _18145_ (.A1(_02323_),
    .A2(_02324_),
    .B1(_02316_),
    .C1(_02320_),
    .X(_02325_));
 sky130_fd_sc_hd__a211oi_2 _18146_ (.A1(_02316_),
    .A2(_02320_),
    .B1(_02323_),
    .C1(_02324_),
    .Y(_02326_));
 sky130_fd_sc_hd__o31a_1 _18147_ (.A1(_10338_),
    .A2(_02325_),
    .A3(_02326_),
    .B1(_02237_),
    .X(_02327_));
 sky130_fd_sc_hd__o2bb2a_1 _18148_ (.A1_N(_10337_),
    .A2_N(_02327_),
    .B1(_02238_),
    .B2(\rbzero.wall_tracer.trackDistY[3] ),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _18149_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .Y(_02328_));
 sky130_fd_sc_hd__or2_1 _18150_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_02329_));
 sky130_fd_sc_hd__o211a_1 _18151_ (.A1(_02323_),
    .A2(_02326_),
    .B1(_02328_),
    .C1(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__a211oi_1 _18152_ (.A1(_02328_),
    .A2(_02329_),
    .B1(_02323_),
    .C1(_02326_),
    .Y(_02331_));
 sky130_fd_sc_hd__o31a_1 _18153_ (.A1(_10338_),
    .A2(_02330_),
    .A3(_02331_),
    .B1(_02237_),
    .X(_02332_));
 sky130_fd_sc_hd__o2bb2a_1 _18154_ (.A1_N(_01652_),
    .A2_N(_02332_),
    .B1(_02250_),
    .B2(\rbzero.wall_tracer.trackDistY[4] ),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _18155_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_02333_));
 sky130_fd_sc_hd__and2_1 _18156_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_02334_));
 sky130_fd_sc_hd__a21oi_1 _18157_ (.A1(\rbzero.wall_tracer.trackDistY[4] ),
    .A2(\rbzero.wall_tracer.stepDistY[4] ),
    .B1(_02330_),
    .Y(_02335_));
 sky130_fd_sc_hd__nor3_1 _18158_ (.A(_02333_),
    .B(_02334_),
    .C(_02335_),
    .Y(_02336_));
 sky130_fd_sc_hd__o21a_1 _18159_ (.A1(_02333_),
    .A2(_02334_),
    .B1(_02335_),
    .X(_02337_));
 sky130_fd_sc_hd__o31a_1 _18160_ (.A1(_09789_),
    .A2(_02336_),
    .A3(_02337_),
    .B1(_02237_),
    .X(_02338_));
 sky130_fd_sc_hd__o2bb2a_1 _18161_ (.A1_N(_01758_),
    .A2_N(_02338_),
    .B1(_02250_),
    .B2(\rbzero.wall_tracer.trackDistY[5] ),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_1 _18162_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02339_));
 sky130_fd_sc_hd__nand2_1 _18163_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02340_));
 sky130_fd_sc_hd__or2b_1 _18164_ (.A(_02339_),
    .B_N(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__o21ba_1 _18165_ (.A1(_02333_),
    .A2(_02335_),
    .B1_N(_02334_),
    .X(_02342_));
 sky130_fd_sc_hd__nor2_1 _18166_ (.A(_02341_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__a21o_1 _18167_ (.A1(_02341_),
    .A2(_02342_),
    .B1(_06102_),
    .X(_02344_));
 sky130_fd_sc_hd__o21ai_1 _18168_ (.A1(_02343_),
    .A2(_02344_),
    .B1(_01879_),
    .Y(_02345_));
 sky130_fd_sc_hd__mux2_1 _18169_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(_02345_),
    .S(_02237_),
    .X(_02346_));
 sky130_fd_sc_hd__clkbuf_1 _18170_ (.A(_02346_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _18171_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _18172_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02348_));
 sky130_fd_sc_hd__or2b_1 _18173_ (.A(_02347_),
    .B_N(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__o21a_1 _18174_ (.A1(_02339_),
    .A2(_02342_),
    .B1(_02340_),
    .X(_02350_));
 sky130_fd_sc_hd__xnor2_1 _18175_ (.A(_02349_),
    .B(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__o21a_1 _18176_ (.A1(_10107_),
    .A2(_02351_),
    .B1(_02235_),
    .X(_02352_));
 sky130_fd_sc_hd__o2bb2a_1 _18177_ (.A1_N(_01984_),
    .A2_N(_02352_),
    .B1(_02250_),
    .B2(\rbzero.wall_tracer.trackDistY[7] ),
    .X(_00568_));
 sky130_fd_sc_hd__or2_1 _18178_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .X(_02353_));
 sky130_fd_sc_hd__nand2_1 _18179_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _18180_ (.A(_02353_),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__o21a_1 _18181_ (.A1(_02347_),
    .A2(_02350_),
    .B1(_02348_),
    .X(_02356_));
 sky130_fd_sc_hd__nor2_1 _18182_ (.A(_02355_),
    .B(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__a21o_1 _18183_ (.A1(_02355_),
    .A2(_02356_),
    .B1(_09760_),
    .X(_02358_));
 sky130_fd_sc_hd__o21a_1 _18184_ (.A1(_02357_),
    .A2(_02358_),
    .B1(_02235_),
    .X(_02359_));
 sky130_fd_sc_hd__o2bb2a_1 _18185_ (.A1_N(_02074_),
    .A2_N(_02359_),
    .B1(_02250_),
    .B2(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_00569_));
 sky130_fd_sc_hd__and2_1 _18186_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_02360_));
 sky130_fd_sc_hd__nor2_1 _18187_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_02361_));
 sky130_fd_sc_hd__nor2_1 _18188_ (.A(_02360_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand2_1 _18189_ (.A(_02354_),
    .B(_02356_),
    .Y(_02363_));
 sky130_fd_sc_hd__and2_1 _18190_ (.A(_02353_),
    .B(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__xnor2_1 _18191_ (.A(_02362_),
    .B(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__o21a_1 _18192_ (.A1(_10107_),
    .A2(_02365_),
    .B1(_02235_),
    .X(_02366_));
 sky130_fd_sc_hd__o2bb2a_1 _18193_ (.A1_N(_02161_),
    .A2_N(_02366_),
    .B1(_02250_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .X(_00570_));
 sky130_fd_sc_hd__a31o_1 _18194_ (.A1(_02353_),
    .A2(_02362_),
    .A3(_02363_),
    .B1(_02360_),
    .X(_02367_));
 sky130_fd_sc_hd__xor2_1 _18195_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .X(_02368_));
 sky130_fd_sc_hd__xnor2_1 _18196_ (.A(_02367_),
    .B(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__o21a_1 _18197_ (.A1(_10107_),
    .A2(_02369_),
    .B1(_02235_),
    .X(_02370_));
 sky130_fd_sc_hd__o2bb2a_1 _18198_ (.A1_N(_02227_),
    .A2_N(_02370_),
    .B1(_02250_),
    .B2(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_00571_));
 sky130_fd_sc_hd__buf_4 _18199_ (.A(_08091_),
    .X(_02371_));
 sky130_fd_sc_hd__and2_1 _18200_ (.A(net43),
    .B(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__clkbuf_1 _18201_ (.A(_02372_),
    .X(_00572_));
 sky130_fd_sc_hd__and2_1 _18202_ (.A(\rbzero.spi_registers.ss_buffer[0] ),
    .B(_02371_),
    .X(_02373_));
 sky130_fd_sc_hd__clkbuf_1 _18203_ (.A(_02373_),
    .X(_00573_));
 sky130_fd_sc_hd__buf_4 _18204_ (.A(\rbzero.spi_registers.spi_done ),
    .X(_02374_));
 sky130_fd_sc_hd__nor2b_2 _18205_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B_N(\rbzero.spi_registers.spi_cmd[2] ),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2b_2 _18206_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B_N(\rbzero.spi_registers.spi_cmd[1] ),
    .Y(_02376_));
 sky130_fd_sc_hd__or2b_1 _18207_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B_N(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_02377_));
 sky130_fd_sc_hd__nor2b_4 _18208_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .B_N(\rbzero.spi_registers.spi_cmd[3] ),
    .Y(_02378_));
 sky130_fd_sc_hd__clkinv_2 _18209_ (.A(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__nand2_4 _18210_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .Y(_02380_));
 sky130_fd_sc_hd__mux2_1 _18211_ (.A0(_02377_),
    .A1(_02379_),
    .S(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__a21bo_1 _18212_ (.A1(_02375_),
    .A2(_02376_),
    .B1_N(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__xor2_1 _18213_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__nor2_2 _18214_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .Y(_02384_));
 sky130_fd_sc_hd__and2_2 _18215_ (.A(_02375_),
    .B(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__nor2_4 _18216_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .Y(_02386_));
 sky130_fd_sc_hd__or3b_1 _18217_ (.A(_02385_),
    .B(_02386_),
    .C_N(_02381_),
    .X(_02387_));
 sky130_fd_sc_hd__xor2_1 _18218_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__or2_1 _18219_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(\rbzero.spi_registers.spi_counter[5] ),
    .X(_02389_));
 sky130_fd_sc_hd__nor4_4 _18220_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(\rbzero.spi_registers.spi_counter[3] ),
    .C(\rbzero.spi_registers.spi_counter[2] ),
    .D(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__or4_1 _18221_ (.A(_02383_),
    .B(_02388_),
    .C(_02389_),
    .D(_02390_),
    .X(_02391_));
 sky130_fd_sc_hd__a21oi_1 _18222_ (.A1(_02375_),
    .A2(_02376_),
    .B1(_02387_),
    .Y(_02392_));
 sky130_fd_sc_hd__a211o_1 _18223_ (.A1(_02386_),
    .A2(_02380_),
    .B1(_02392_),
    .C1(_02385_),
    .X(_02393_));
 sky130_fd_sc_hd__xnor2_1 _18224_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__or2_2 _18225_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .B(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_02395_));
 sky130_fd_sc_hd__o21a_1 _18226_ (.A1(_02395_),
    .A2(_02380_),
    .B1(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02396_));
 sky130_fd_sc_hd__a22oi_1 _18227_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02392_),
    .B1(_02396_),
    .B2(\rbzero.spi_registers.spi_counter[2] ),
    .Y(_02397_));
 sky130_fd_sc_hd__o221a_1 _18228_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02392_),
    .B1(_02396_),
    .B2(\rbzero.spi_registers.spi_counter[2] ),
    .C1(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__or3b_1 _18229_ (.A(_02391_),
    .B(_02394_),
    .C_N(_02398_),
    .X(_02399_));
 sky130_fd_sc_hd__and2b_1 _18230_ (.A_N(\rbzero.spi_registers.sclk_buffer[2] ),
    .B(\rbzero.spi_registers.sclk_buffer[1] ),
    .X(_02400_));
 sky130_fd_sc_hd__nor2_1 _18231_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_04094_),
    .Y(_02401_));
 sky130_fd_sc_hd__and4bb_1 _18232_ (.A_N(_02374_),
    .B_N(_02399_),
    .C(_02400_),
    .D(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__clkbuf_1 _18233_ (.A(_02402_),
    .X(_00574_));
 sky130_fd_sc_hd__and2_1 _18234_ (.A(net44),
    .B(_02371_),
    .X(_02403_));
 sky130_fd_sc_hd__clkbuf_1 _18235_ (.A(_02403_),
    .X(_00575_));
 sky130_fd_sc_hd__and2_1 _18236_ (.A(\rbzero.spi_registers.mosi_buffer[0] ),
    .B(_02371_),
    .X(_02404_));
 sky130_fd_sc_hd__clkbuf_1 _18237_ (.A(_02404_),
    .X(_00576_));
 sky130_fd_sc_hd__clkbuf_4 _18238_ (.A(_09723_),
    .X(_02405_));
 sky130_fd_sc_hd__clkbuf_4 _18239_ (.A(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__nor2_1 _18240_ (.A(_05291_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _18241_ (.A(_05291_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02408_));
 sky130_fd_sc_hd__or2b_1 _18242_ (.A(_02407_),
    .B_N(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__or2_1 _18243_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .X(_02410_));
 sky130_fd_sc_hd__nor2_1 _18244_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02411_));
 sky130_fd_sc_hd__nand2_1 _18245_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_02412_));
 sky130_fd_sc_hd__or2_1 _18246_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_02413_));
 sky130_fd_sc_hd__and4_1 _18247_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .C(_02412_),
    .D(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__a21oi_1 _18248_ (.A1(\rbzero.debug_overlay.vplaneX[-8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-8] ),
    .B1(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__nand2_1 _18249_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02416_));
 sky130_fd_sc_hd__o21ai_1 _18250_ (.A1(_02411_),
    .A2(_02415_),
    .B1(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__nand2_1 _18251_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .Y(_02418_));
 sky130_fd_sc_hd__a21boi_1 _18252_ (.A1(_02410_),
    .A2(_02417_),
    .B1_N(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__xnor2_1 _18253_ (.A(_02409_),
    .B(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__nor2_1 _18254_ (.A(_09731_),
    .B(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__a221o_1 _18255_ (.A1(_05290_),
    .A2(_08113_),
    .B1(_02406_),
    .B2(\rbzero.wall_tracer.rayAddendX[-5] ),
    .C1(_02421_),
    .X(_00577_));
 sky130_fd_sc_hd__xnor2_1 _18256_ (.A(_05292_),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .Y(_02422_));
 sky130_fd_sc_hd__o21ai_1 _18257_ (.A1(_02407_),
    .A2(_02419_),
    .B1(_02408_),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_1 _18258_ (.A(_02422_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__clkbuf_4 _18259_ (.A(_08112_),
    .X(_02425_));
 sky130_fd_sc_hd__a211o_1 _18260_ (.A1(_02422_),
    .A2(_02423_),
    .B1(_02424_),
    .C1(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__nand2_1 _18261_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(_05290_),
    .Y(_02427_));
 sky130_fd_sc_hd__or2_1 _18262_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(_05290_),
    .X(_02428_));
 sky130_fd_sc_hd__a31o_1 _18263_ (.A1(_02425_),
    .A2(_02427_),
    .A3(_02428_),
    .B1(_09728_),
    .X(_02429_));
 sky130_fd_sc_hd__a22o_1 _18264_ (.A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_09738_),
    .B1(_02426_),
    .B2(_02429_),
    .X(_00578_));
 sky130_fd_sc_hd__or2_1 _18265_ (.A(_08111_),
    .B(_09722_),
    .X(_02430_));
 sky130_fd_sc_hd__clkbuf_4 _18266_ (.A(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__buf_4 _18267_ (.A(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__nor2_1 _18268_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02433_));
 sky130_fd_sc_hd__and2_1 _18269_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .X(_02434_));
 sky130_fd_sc_hd__a21o_1 _18270_ (.A1(_05292_),
    .A2(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B1(_02423_),
    .X(_02435_));
 sky130_fd_sc_hd__o21ai_1 _18271_ (.A1(_05292_),
    .A2(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B1(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__o21ai_1 _18272_ (.A1(_02433_),
    .A2(_02434_),
    .B1(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__o311a_1 _18273_ (.A1(_02433_),
    .A2(_02434_),
    .A3(_02436_),
    .B1(_02437_),
    .C1(_04478_),
    .X(_02438_));
 sky130_fd_sc_hd__clkbuf_4 _18274_ (.A(_08112_),
    .X(_02439_));
 sky130_fd_sc_hd__or2_1 _18275_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02428_),
    .X(_02440_));
 sky130_fd_sc_hd__nand2_1 _18276_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02428_),
    .Y(_02441_));
 sky130_fd_sc_hd__a31o_1 _18277_ (.A1(_02439_),
    .A2(_02440_),
    .A3(_02441_),
    .B1(_09724_),
    .X(_02442_));
 sky130_fd_sc_hd__o22a_1 _18278_ (.A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A2(_02432_),
    .B1(_02438_),
    .B2(_02442_),
    .X(_00579_));
 sky130_fd_sc_hd__clkbuf_4 _18279_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_02443_));
 sky130_fd_sc_hd__nor2_1 _18280_ (.A(_02443_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_02444_));
 sky130_fd_sc_hd__and2_1 _18281_ (.A(_02443_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02445_));
 sky130_fd_sc_hd__nand2_1 _18282_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02446_));
 sky130_fd_sc_hd__o21ai_1 _18283_ (.A1(_02433_),
    .A2(_02436_),
    .B1(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__or3_1 _18284_ (.A(_02444_),
    .B(_02445_),
    .C(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__o21ai_1 _18285_ (.A1(_02444_),
    .A2(_02445_),
    .B1(_02447_),
    .Y(_02449_));
 sky130_fd_sc_hd__a21oi_1 _18286_ (.A1(_02448_),
    .A2(_02449_),
    .B1(_08113_),
    .Y(_02450_));
 sky130_fd_sc_hd__nand2_1 _18287_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_02440_),
    .Y(_02451_));
 sky130_fd_sc_hd__or2_1 _18288_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_02440_),
    .X(_02452_));
 sky130_fd_sc_hd__a31o_1 _18289_ (.A1(_02439_),
    .A2(_02451_),
    .A3(_02452_),
    .B1(_09724_),
    .X(_02453_));
 sky130_fd_sc_hd__o22a_1 _18290_ (.A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A2(_02432_),
    .B1(_02450_),
    .B2(_02453_),
    .X(_00580_));
 sky130_fd_sc_hd__or2_1 _18291_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02454_));
 sky130_fd_sc_hd__nand2_1 _18292_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_02455_));
 sky130_fd_sc_hd__or2_1 _18293_ (.A(_02443_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02456_));
 sky130_fd_sc_hd__a21o_1 _18294_ (.A1(_02456_),
    .A2(_02447_),
    .B1(_02445_),
    .X(_02457_));
 sky130_fd_sc_hd__a21oi_1 _18295_ (.A1(_02454_),
    .A2(_02455_),
    .B1(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__a31o_1 _18296_ (.A1(_02454_),
    .A2(_02455_),
    .A3(_02457_),
    .B1(_09730_),
    .X(_02459_));
 sky130_fd_sc_hd__inv_2 _18297_ (.A(_05290_),
    .Y(_02460_));
 sky130_fd_sc_hd__o31a_1 _18298_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(\rbzero.debug_overlay.vplaneX[-7] ),
    .A3(\rbzero.debug_overlay.vplaneX[-8] ),
    .B1(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__xnor2_1 _18299_ (.A(_05291_),
    .B(_02461_),
    .Y(_02462_));
 sky130_fd_sc_hd__o2bb2a_1 _18300_ (.A1_N(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A2_N(_02405_),
    .B1(_02462_),
    .B2(_04469_),
    .X(_02463_));
 sky130_fd_sc_hd__o21ai_1 _18301_ (.A1(_02458_),
    .A2(_02459_),
    .B1(_02463_),
    .Y(_00581_));
 sky130_fd_sc_hd__a21bo_1 _18302_ (.A1(_02454_),
    .A2(_02457_),
    .B1_N(_02455_),
    .X(_02464_));
 sky130_fd_sc_hd__clkbuf_4 _18303_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_02465_));
 sky130_fd_sc_hd__nor2_1 _18304_ (.A(_02465_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_02466_));
 sky130_fd_sc_hd__and2_1 _18305_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_02467_));
 sky130_fd_sc_hd__or2_1 _18306_ (.A(_02466_),
    .B(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__xnor2_1 _18307_ (.A(_02464_),
    .B(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__or2_1 _18308_ (.A(_05292_),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_02470_));
 sky130_fd_sc_hd__nand2_1 _18309_ (.A(_05292_),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .Y(_02471_));
 sky130_fd_sc_hd__nand2_1 _18310_ (.A(_02470_),
    .B(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__nor2_1 _18311_ (.A(_05291_),
    .B(_02452_),
    .Y(_02473_));
 sky130_fd_sc_hd__a21oi_1 _18312_ (.A1(_05291_),
    .A2(_05290_),
    .B1(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__xnor2_1 _18313_ (.A(_02472_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__mux2_1 _18314_ (.A0(_02469_),
    .A1(_02475_),
    .S(_08112_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _18315_ (.A0(\rbzero.wall_tracer.rayAddendX[0] ),
    .A1(_02476_),
    .S(_02431_),
    .X(_02477_));
 sky130_fd_sc_hd__clkbuf_1 _18316_ (.A(_02477_),
    .X(_00582_));
 sky130_fd_sc_hd__buf_4 _18317_ (.A(_09728_),
    .X(_02478_));
 sky130_fd_sc_hd__nand2_1 _18318_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_02479_));
 sky130_fd_sc_hd__or2_1 _18319_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02480_));
 sky130_fd_sc_hd__o21a_1 _18320_ (.A1(_02465_),
    .A2(\rbzero.wall_tracer.rayAddendX[0] ),
    .B1(_02464_),
    .X(_02481_));
 sky130_fd_sc_hd__a211o_1 _18321_ (.A1(_02479_),
    .A2(_02480_),
    .B1(_02481_),
    .C1(_02467_),
    .X(_02482_));
 sky130_fd_sc_hd__o211ai_2 _18322_ (.A1(_02467_),
    .A2(_02481_),
    .B1(_02480_),
    .C1(_02479_),
    .Y(_02483_));
 sky130_fd_sc_hd__a21oi_1 _18323_ (.A1(_05291_),
    .A2(_05290_),
    .B1(_02472_),
    .Y(_02484_));
 sky130_fd_sc_hd__nor2_1 _18324_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_02485_));
 sky130_fd_sc_hd__and2_1 _18325_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_02486_));
 sky130_fd_sc_hd__nor2_1 _18326_ (.A(_02485_),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__xnor2_1 _18327_ (.A(_02470_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__o21a_1 _18328_ (.A1(_02473_),
    .A2(_02484_),
    .B1(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__inv_2 _18329_ (.A(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__or3_1 _18330_ (.A(_02473_),
    .B(_02488_),
    .C(_02484_),
    .X(_02491_));
 sky130_fd_sc_hd__a32o_1 _18331_ (.A1(_02425_),
    .A2(_02490_),
    .A3(_02491_),
    .B1(_02406_),
    .B2(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02492_));
 sky130_fd_sc_hd__a31o_1 _18332_ (.A1(_02478_),
    .A2(_02482_),
    .A3(_02483_),
    .B1(_02492_),
    .X(_00583_));
 sky130_fd_sc_hd__buf_2 _18333_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_02493_));
 sky130_fd_sc_hd__buf_2 _18334_ (.A(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__clkbuf_4 _18335_ (.A(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__xnor2_1 _18336_ (.A(_02495_),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_02496_));
 sky130_fd_sc_hd__a21oi_1 _18337_ (.A1(_02479_),
    .A2(_02483_),
    .B1(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__a311oi_1 _18338_ (.A1(_02479_),
    .A2(_02483_),
    .A3(_02496_),
    .B1(_02497_),
    .C1(_08113_),
    .Y(_02498_));
 sky130_fd_sc_hd__xor2_1 _18339_ (.A(_02443_),
    .B(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_02499_));
 sky130_fd_sc_hd__o31ai_1 _18340_ (.A1(_02470_),
    .A2(_02485_),
    .A3(_02486_),
    .B1(_02490_),
    .Y(_02500_));
 sky130_fd_sc_hd__xnor2_1 _18341_ (.A(_02499_),
    .B(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__xnor2_1 _18342_ (.A(_02485_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__a21o_1 _18343_ (.A1(_08113_),
    .A2(_02502_),
    .B1(_02406_),
    .X(_02503_));
 sky130_fd_sc_hd__o22a_1 _18344_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(_02432_),
    .B1(_02498_),
    .B2(_02503_),
    .X(_00584_));
 sky130_fd_sc_hd__and2_1 _18345_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02504_));
 sky130_fd_sc_hd__nor2_1 _18346_ (.A(_02493_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02505_));
 sky130_fd_sc_hd__o21ai_1 _18347_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[1] ),
    .B1(_02493_),
    .Y(_02506_));
 sky130_fd_sc_hd__o21bai_1 _18348_ (.A1(_02493_),
    .A2(\rbzero.wall_tracer.rayAddendX[2] ),
    .B1_N(_02483_),
    .Y(_02507_));
 sky130_fd_sc_hd__o211ai_1 _18349_ (.A1(_02504_),
    .A2(_02505_),
    .B1(_02506_),
    .C1(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__a211o_1 _18350_ (.A1(_02506_),
    .A2(_02507_),
    .B1(_02504_),
    .C1(_02505_),
    .X(_02509_));
 sky130_fd_sc_hd__or2_1 _18351_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05291_),
    .X(_02510_));
 sky130_fd_sc_hd__nand2_1 _18352_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05291_),
    .Y(_02511_));
 sky130_fd_sc_hd__and4bb_1 _18353_ (.A_N(_02443_),
    .B_N(\rbzero.debug_overlay.vplaneX[-6] ),
    .C(_02510_),
    .D(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__a2bb2o_1 _18354_ (.A1_N(_02443_),
    .A2_N(\rbzero.debug_overlay.vplaneX[-6] ),
    .B1(_02510_),
    .B2(_02511_),
    .X(_02513_));
 sky130_fd_sc_hd__and2b_1 _18355_ (.A_N(_02512_),
    .B(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__o21a_1 _18356_ (.A1(_02489_),
    .A2(_02499_),
    .B1(_02485_),
    .X(_02515_));
 sky130_fd_sc_hd__a21o_1 _18357_ (.A1(_02499_),
    .A2(_02500_),
    .B1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__and2_1 _18358_ (.A(_02514_),
    .B(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__o21ai_1 _18359_ (.A1(_02514_),
    .A2(_02516_),
    .B1(_02425_),
    .Y(_02518_));
 sky130_fd_sc_hd__a2bb2o_1 _18360_ (.A1_N(_02517_),
    .A2_N(_02518_),
    .B1(\rbzero.wall_tracer.rayAddendX[3] ),
    .B2(_02405_),
    .X(_02519_));
 sky130_fd_sc_hd__a31o_1 _18361_ (.A1(_02478_),
    .A2(_02508_),
    .A3(_02509_),
    .B1(_02519_),
    .X(_00585_));
 sky130_fd_sc_hd__nand2_1 _18362_ (.A(_02495_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02520_));
 sky130_fd_sc_hd__xor2_1 _18363_ (.A(_02493_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_02521_));
 sky130_fd_sc_hd__a21oi_1 _18364_ (.A1(_02520_),
    .A2(_02509_),
    .B1(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__a31o_1 _18365_ (.A1(_02520_),
    .A2(_02509_),
    .A3(_02521_),
    .B1(_08111_),
    .X(_02523_));
 sky130_fd_sc_hd__xor2_1 _18366_ (.A(_02465_),
    .B(_05292_),
    .X(_02524_));
 sky130_fd_sc_hd__o21ai_1 _18367_ (.A1(_02512_),
    .A2(_02517_),
    .B1(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__or3_1 _18368_ (.A(_02512_),
    .B(_02517_),
    .C(_02524_),
    .X(_02526_));
 sky130_fd_sc_hd__and2_1 _18369_ (.A(_02525_),
    .B(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__xnor2_1 _18370_ (.A(_02510_),
    .B(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__o22a_1 _18371_ (.A1(_02522_),
    .A2(_02523_),
    .B1(_02528_),
    .B2(_04469_),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _18372_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02529_),
    .S(_02431_),
    .X(_02530_));
 sky130_fd_sc_hd__clkbuf_1 _18373_ (.A(_02530_),
    .X(_00586_));
 sky130_fd_sc_hd__or2b_1 _18374_ (.A(_02509_),
    .B_N(_02521_),
    .X(_02531_));
 sky130_fd_sc_hd__o21ai_1 _18375_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02495_),
    .Y(_02532_));
 sky130_fd_sc_hd__nand2_1 _18376_ (.A(_02493_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02533_));
 sky130_fd_sc_hd__or2_1 _18377_ (.A(_02493_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_02534_));
 sky130_fd_sc_hd__nand2_1 _18378_ (.A(_02533_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__a21o_1 _18379_ (.A1(_02531_),
    .A2(_02532_),
    .B1(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__nand3_1 _18380_ (.A(_02535_),
    .B(_02531_),
    .C(_02532_),
    .Y(_02537_));
 sky130_fd_sc_hd__nor2_1 _18381_ (.A(_02493_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .Y(_02538_));
 sky130_fd_sc_hd__and2_1 _18382_ (.A(_02493_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_02539_));
 sky130_fd_sc_hd__o22a_1 _18383_ (.A1(_02465_),
    .A2(_05292_),
    .B1(_02538_),
    .B2(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__nor4_1 _18384_ (.A(_02465_),
    .B(_05292_),
    .C(_02538_),
    .D(_02539_),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _18385_ (.A(_02540_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__a2bb2o_1 _18386_ (.A1_N(_02517_),
    .A2_N(_02524_),
    .B1(_02525_),
    .B2(_02510_),
    .X(_02543_));
 sky130_fd_sc_hd__xnor2_1 _18387_ (.A(_02542_),
    .B(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__a22o_1 _18388_ (.A1(\rbzero.wall_tracer.rayAddendX[5] ),
    .A2(_02405_),
    .B1(_02544_),
    .B2(_02439_),
    .X(_02545_));
 sky130_fd_sc_hd__a31o_1 _18389_ (.A1(_02478_),
    .A2(_02536_),
    .A3(_02537_),
    .B1(_02545_),
    .X(_00587_));
 sky130_fd_sc_hd__xnor2_1 _18390_ (.A(_02494_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_02546_));
 sky130_fd_sc_hd__a21o_1 _18391_ (.A1(_02533_),
    .A2(_02536_),
    .B1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__nand3_1 _18392_ (.A(_02533_),
    .B(_02536_),
    .C(_02546_),
    .Y(_02548_));
 sky130_fd_sc_hd__or2_1 _18393_ (.A(_02493_),
    .B(_02443_),
    .X(_02549_));
 sky130_fd_sc_hd__nand2_1 _18394_ (.A(_02494_),
    .B(_02443_),
    .Y(_02550_));
 sky130_fd_sc_hd__a21o_1 _18395_ (.A1(_02549_),
    .A2(_02550_),
    .B1(_02538_),
    .X(_02551_));
 sky130_fd_sc_hd__nand2_1 _18396_ (.A(_02443_),
    .B(_02538_),
    .Y(_02552_));
 sky130_fd_sc_hd__nand2_1 _18397_ (.A(_02551_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__o21bai_1 _18398_ (.A1(_02540_),
    .A2(_02543_),
    .B1_N(_02541_),
    .Y(_02554_));
 sky130_fd_sc_hd__xnor2_1 _18399_ (.A(_02553_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__a22o_1 _18400_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(_02405_),
    .B1(_02555_),
    .B2(_02439_),
    .X(_02556_));
 sky130_fd_sc_hd__a31o_1 _18401_ (.A1(_02478_),
    .A2(_02547_),
    .A3(_02548_),
    .B1(_02556_),
    .X(_00588_));
 sky130_fd_sc_hd__nand2_1 _18402_ (.A(_02494_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_02557_));
 sky130_fd_sc_hd__or2_1 _18403_ (.A(_02494_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02558_));
 sky130_fd_sc_hd__nor3_1 _18404_ (.A(_02535_),
    .B(_02531_),
    .C(_02546_),
    .Y(_02559_));
 sky130_fd_sc_hd__o41a_1 _18405_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .A3(\rbzero.wall_tracer.rayAddendX[4] ),
    .A4(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02494_),
    .X(_02560_));
 sky130_fd_sc_hd__a211o_1 _18406_ (.A1(_02557_),
    .A2(_02558_),
    .B1(_02559_),
    .C1(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__o211ai_2 _18407_ (.A1(_02559_),
    .A2(_02560_),
    .B1(_02557_),
    .C1(_02558_),
    .Y(_02562_));
 sky130_fd_sc_hd__inv_2 _18408_ (.A(_02552_),
    .Y(_02563_));
 sky130_fd_sc_hd__and3_1 _18409_ (.A(_02551_),
    .B(_02552_),
    .C(_02554_),
    .X(_02564_));
 sky130_fd_sc_hd__nor2_1 _18410_ (.A(_02494_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .Y(_02565_));
 sky130_fd_sc_hd__and2_1 _18411_ (.A(_02494_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_02566_));
 sky130_fd_sc_hd__o21ai_1 _18412_ (.A1(_02565_),
    .A2(_02566_),
    .B1(_02549_),
    .Y(_02567_));
 sky130_fd_sc_hd__or3_1 _18413_ (.A(_02549_),
    .B(_02565_),
    .C(_02566_),
    .X(_02568_));
 sky130_fd_sc_hd__o211ai_2 _18414_ (.A1(_02563_),
    .A2(_02564_),
    .B1(_02567_),
    .C1(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__a211o_1 _18415_ (.A1(_02567_),
    .A2(_02568_),
    .B1(_02563_),
    .C1(_02564_),
    .X(_02570_));
 sky130_fd_sc_hd__a32o_1 _18416_ (.A1(_02425_),
    .A2(_02569_),
    .A3(_02570_),
    .B1(_02406_),
    .B2(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02571_));
 sky130_fd_sc_hd__a31o_1 _18417_ (.A1(_02478_),
    .A2(_02561_),
    .A3(_02562_),
    .B1(_02571_),
    .X(_00589_));
 sky130_fd_sc_hd__xnor2_1 _18418_ (.A(_02494_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_02572_));
 sky130_fd_sc_hd__a21oi_1 _18419_ (.A1(_02557_),
    .A2(_02562_),
    .B1(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__a31o_1 _18420_ (.A1(_02557_),
    .A2(_02562_),
    .A3(_02572_),
    .B1(_08112_),
    .X(_02574_));
 sky130_fd_sc_hd__nor2_1 _18421_ (.A(_02573_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__inv_2 _18422_ (.A(_02465_),
    .Y(_02576_));
 sky130_fd_sc_hd__a21oi_1 _18423_ (.A1(_02465_),
    .A2(\rbzero.debug_overlay.vplaneX[-1] ),
    .B1(_02494_),
    .Y(_02577_));
 sky130_fd_sc_hd__a21oi_1 _18424_ (.A1(_02495_),
    .A2(_02465_),
    .B1(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__a21oi_1 _18425_ (.A1(_02576_),
    .A2(_02565_),
    .B1(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__a21o_1 _18426_ (.A1(_02568_),
    .A2(_02569_),
    .B1(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__nand3_1 _18427_ (.A(_02568_),
    .B(_02569_),
    .C(_02579_),
    .Y(_02581_));
 sky130_fd_sc_hd__a31o_1 _18428_ (.A1(_02439_),
    .A2(_02580_),
    .A3(_02581_),
    .B1(_09724_),
    .X(_02582_));
 sky130_fd_sc_hd__o22a_1 _18429_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(_02432_),
    .B1(_02575_),
    .B2(_02582_),
    .X(_00590_));
 sky130_fd_sc_hd__or2_1 _18430_ (.A(_02495_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_1 _18431_ (.A(_02495_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_1 _18432_ (.A(_02583_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__o21ai_1 _18433_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[7] ),
    .B1(_02495_),
    .Y(_02586_));
 sky130_fd_sc_hd__o21ai_1 _18434_ (.A1(_02562_),
    .A2(_02572_),
    .B1(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__xnor2_1 _18435_ (.A(_02585_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__inv_2 _18436_ (.A(_02495_),
    .Y(_02589_));
 sky130_fd_sc_hd__a21oi_1 _18437_ (.A1(_02589_),
    .A2(_02576_),
    .B1(_02580_),
    .Y(_02590_));
 sky130_fd_sc_hd__a211o_1 _18438_ (.A1(_02577_),
    .A2(_02580_),
    .B1(_02590_),
    .C1(_04469_),
    .X(_02591_));
 sky130_fd_sc_hd__o221a_1 _18439_ (.A1(\rbzero.wall_tracer.rayAddendX[9] ),
    .A2(_02432_),
    .B1(_09731_),
    .B2(_02588_),
    .C1(_02591_),
    .X(_00591_));
 sky130_fd_sc_hd__a21bo_1 _18440_ (.A1(_02583_),
    .A2(_02587_),
    .B1_N(_02584_),
    .X(_02592_));
 sky130_fd_sc_hd__xnor2_1 _18441_ (.A(_02495_),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_02593_));
 sky130_fd_sc_hd__xnor2_1 _18442_ (.A(_02592_),
    .B(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__o211a_1 _18443_ (.A1(_02465_),
    .A2(_02580_),
    .B1(_08112_),
    .C1(_02589_),
    .X(_02595_));
 sky130_fd_sc_hd__o22a_1 _18444_ (.A1(_02439_),
    .A2(_02594_),
    .B1(_02595_),
    .B2(_09728_),
    .X(_02596_));
 sky130_fd_sc_hd__a21o_1 _18445_ (.A1(\rbzero.wall_tracer.rayAddendX[10] ),
    .A2(_09725_),
    .B1(_02596_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _18446_ (.A0(\rbzero.debug_overlay.playerY[0] ),
    .A1(_06113_),
    .S(_09784_),
    .X(_02597_));
 sky130_fd_sc_hd__o21a_2 _18447_ (.A1(_06156_),
    .A2(_06163_),
    .B1(_06254_),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _18448_ (.A0(_06086_),
    .A1(_02597_),
    .S(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__clkbuf_1 _18449_ (.A(_02599_),
    .X(_00593_));
 sky130_fd_sc_hd__nor2_1 _18450_ (.A(_06086_),
    .B(_06088_),
    .Y(_02600_));
 sky130_fd_sc_hd__nand2_1 _18451_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(_09760_),
    .Y(_02601_));
 sky130_fd_sc_hd__o311a_1 _18452_ (.A1(_09760_),
    .A2(_06089_),
    .A3(_02600_),
    .B1(_02601_),
    .C1(_02598_),
    .X(_02602_));
 sky130_fd_sc_hd__a21oi_1 _18453_ (.A1(_06084_),
    .A2(_06255_),
    .B1(_02602_),
    .Y(_00594_));
 sky130_fd_sc_hd__or3_1 _18454_ (.A(_06085_),
    .B(_06089_),
    .C(_06090_),
    .X(_02603_));
 sky130_fd_sc_hd__and3_1 _18455_ (.A(_08100_),
    .B(_06091_),
    .C(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__a211o_1 _18456_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_10107_),
    .B1(_06255_),
    .C1(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__o21a_1 _18457_ (.A1(\rbzero.map_rom.b6 ),
    .A2(_02598_),
    .B1(_02605_),
    .X(_00595_));
 sky130_fd_sc_hd__or2_1 _18458_ (.A(_06080_),
    .B(_06082_),
    .X(_02606_));
 sky130_fd_sc_hd__xnor2_1 _18459_ (.A(_06092_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__mux2_1 _18460_ (.A0(\rbzero.debug_overlay.playerY[3] ),
    .A1(_02607_),
    .S(_09784_),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _18461_ (.A0(\rbzero.map_rom.a6 ),
    .A1(_02608_),
    .S(_02598_),
    .X(_02609_));
 sky130_fd_sc_hd__clkbuf_1 _18462_ (.A(_02609_),
    .X(_00596_));
 sky130_fd_sc_hd__or3_1 _18463_ (.A(_06094_),
    .B(_06080_),
    .C(_06093_),
    .X(_02610_));
 sky130_fd_sc_hd__nor2_1 _18464_ (.A(_09760_),
    .B(_06095_),
    .Y(_02611_));
 sky130_fd_sc_hd__a221o_1 _18465_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_09789_),
    .B1(_02610_),
    .B2(_02611_),
    .C1(_06255_),
    .X(_02612_));
 sky130_fd_sc_hd__o21a_1 _18466_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(_02598_),
    .B1(_02612_),
    .X(_00597_));
 sky130_fd_sc_hd__a21oi_1 _18467_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(_06081_),
    .B1(_06095_),
    .Y(_02613_));
 sky130_fd_sc_hd__xnor2_1 _18468_ (.A(_06078_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__mux2_1 _18469_ (.A0(\rbzero.debug_overlay.playerY[5] ),
    .A1(_02614_),
    .S(_09784_),
    .X(_02615_));
 sky130_fd_sc_hd__mux2_1 _18470_ (.A0(\rbzero.wall_tracer.mapY[5] ),
    .A1(_02615_),
    .S(_02598_),
    .X(_02616_));
 sky130_fd_sc_hd__clkbuf_1 _18471_ (.A(_02616_),
    .X(_00598_));
 sky130_fd_sc_hd__and3_1 _18472_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .B(_02399_),
    .C(_02400_),
    .X(_02617_));
 sky130_fd_sc_hd__a21o_1 _18473_ (.A1(_02399_),
    .A2(_02400_),
    .B1(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02618_));
 sky130_fd_sc_hd__and3b_1 _18474_ (.A_N(_02617_),
    .B(_02618_),
    .C(_02401_),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _18475_ (.A(_02619_),
    .X(_00599_));
 sky130_fd_sc_hd__and2_1 _18476_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(_02617_),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_2 _18477_ (.A(_02401_),
    .X(_02621_));
 sky130_fd_sc_hd__o21ai_1 _18478_ (.A1(\rbzero.spi_registers.spi_counter[1] ),
    .A2(_02617_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__nor2_1 _18479_ (.A(_02620_),
    .B(_02622_),
    .Y(_00600_));
 sky130_fd_sc_hd__and3_1 _18480_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(\rbzero.spi_registers.spi_counter[1] ),
    .C(_02617_),
    .X(_02623_));
 sky130_fd_sc_hd__o21ai_1 _18481_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(_02620_),
    .B1(_02621_),
    .Y(_02624_));
 sky130_fd_sc_hd__nor2_1 _18482_ (.A(_02623_),
    .B(_02624_),
    .Y(_00601_));
 sky130_fd_sc_hd__and2_1 _18483_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02623_),
    .X(_02625_));
 sky130_fd_sc_hd__o21ai_1 _18484_ (.A1(\rbzero.spi_registers.spi_counter[3] ),
    .A2(_02623_),
    .B1(_02621_),
    .Y(_02626_));
 sky130_fd_sc_hd__nor2_1 _18485_ (.A(_02625_),
    .B(_02626_),
    .Y(_00602_));
 sky130_fd_sc_hd__and3_1 _18486_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(\rbzero.spi_registers.spi_counter[3] ),
    .C(_02623_),
    .X(_02627_));
 sky130_fd_sc_hd__o21ai_1 _18487_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_02625_),
    .B1(_02621_),
    .Y(_02628_));
 sky130_fd_sc_hd__nor2_1 _18488_ (.A(_02627_),
    .B(_02628_),
    .Y(_00603_));
 sky130_fd_sc_hd__and2_1 _18489_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(_02627_),
    .X(_02629_));
 sky130_fd_sc_hd__o21ai_1 _18490_ (.A1(\rbzero.spi_registers.spi_counter[5] ),
    .A2(_02627_),
    .B1(_02621_),
    .Y(_02630_));
 sky130_fd_sc_hd__nor2_1 _18491_ (.A(_02629_),
    .B(_02630_),
    .Y(_00604_));
 sky130_fd_sc_hd__o21ai_1 _18492_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02629_),
    .B1(_02621_),
    .Y(_02631_));
 sky130_fd_sc_hd__a21oi_1 _18493_ (.A1(\rbzero.spi_registers.spi_counter[6] ),
    .A2(_02629_),
    .B1(_02631_),
    .Y(_00605_));
 sky130_fd_sc_hd__buf_4 _18494_ (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .X(_02632_));
 sky130_fd_sc_hd__nor3b_4 _18495_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_02390_),
    .C_N(_02400_),
    .Y(_02633_));
 sky130_fd_sc_hd__clkbuf_4 _18496_ (.A(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__or3b_4 _18497_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_02390_),
    .C_N(_02400_),
    .X(_02635_));
 sky130_fd_sc_hd__buf_2 _18498_ (.A(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__or2_1 _18499_ (.A(\rbzero.spi_registers.mosi ),
    .B(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__buf_4 _18500_ (.A(_08091_),
    .X(_02638_));
 sky130_fd_sc_hd__buf_4 _18501_ (.A(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__o211a_1 _18502_ (.A1(_02632_),
    .A2(_02634_),
    .B1(_02637_),
    .C1(_02639_),
    .X(_00606_));
 sky130_fd_sc_hd__buf_4 _18503_ (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .X(_02640_));
 sky130_fd_sc_hd__or2_1 _18504_ (.A(_02632_),
    .B(_02636_),
    .X(_02641_));
 sky130_fd_sc_hd__o211a_1 _18505_ (.A1(_02640_),
    .A2(_02634_),
    .B1(_02641_),
    .C1(_02639_),
    .X(_00607_));
 sky130_fd_sc_hd__buf_4 _18506_ (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .X(_02642_));
 sky130_fd_sc_hd__or2_1 _18507_ (.A(_02640_),
    .B(_02636_),
    .X(_02643_));
 sky130_fd_sc_hd__o211a_1 _18508_ (.A1(_02642_),
    .A2(_02634_),
    .B1(_02643_),
    .C1(_02639_),
    .X(_00608_));
 sky130_fd_sc_hd__buf_4 _18509_ (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .X(_02644_));
 sky130_fd_sc_hd__or2_1 _18510_ (.A(_02642_),
    .B(_02636_),
    .X(_02645_));
 sky130_fd_sc_hd__o211a_1 _18511_ (.A1(_02644_),
    .A2(_02634_),
    .B1(_02645_),
    .C1(_02639_),
    .X(_00609_));
 sky130_fd_sc_hd__buf_4 _18512_ (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .X(_02646_));
 sky130_fd_sc_hd__or2_1 _18513_ (.A(_02644_),
    .B(_02636_),
    .X(_02647_));
 sky130_fd_sc_hd__o211a_1 _18514_ (.A1(_02646_),
    .A2(_02634_),
    .B1(_02647_),
    .C1(_02639_),
    .X(_00610_));
 sky130_fd_sc_hd__buf_4 _18515_ (.A(\rbzero.spi_registers.spi_buffer[5] ),
    .X(_02648_));
 sky130_fd_sc_hd__or2_1 _18516_ (.A(_02646_),
    .B(_02636_),
    .X(_02649_));
 sky130_fd_sc_hd__o211a_1 _18517_ (.A1(_02648_),
    .A2(_02634_),
    .B1(_02649_),
    .C1(_02639_),
    .X(_00611_));
 sky130_fd_sc_hd__or2_1 _18518_ (.A(_02648_),
    .B(_02636_),
    .X(_02650_));
 sky130_fd_sc_hd__o211a_1 _18519_ (.A1(\rbzero.spi_registers.spi_buffer[6] ),
    .A2(_02634_),
    .B1(_02650_),
    .C1(_02639_),
    .X(_00612_));
 sky130_fd_sc_hd__or2_1 _18520_ (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .B(_02636_),
    .X(_02651_));
 sky130_fd_sc_hd__o211a_1 _18521_ (.A1(\rbzero.spi_registers.spi_buffer[7] ),
    .A2(_02634_),
    .B1(_02651_),
    .C1(_02639_),
    .X(_00613_));
 sky130_fd_sc_hd__or2_1 _18522_ (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .B(_02636_),
    .X(_02652_));
 sky130_fd_sc_hd__clkbuf_8 _18523_ (.A(_08092_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_4 _18524_ (.A(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__o211a_1 _18525_ (.A1(\rbzero.spi_registers.spi_buffer[8] ),
    .A2(_02634_),
    .B1(_02652_),
    .C1(_02654_),
    .X(_00614_));
 sky130_fd_sc_hd__or2_1 _18526_ (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .B(_02636_),
    .X(_02655_));
 sky130_fd_sc_hd__o211a_1 _18527_ (.A1(\rbzero.spi_registers.spi_buffer[9] ),
    .A2(_02634_),
    .B1(_02655_),
    .C1(_02654_),
    .X(_00615_));
 sky130_fd_sc_hd__buf_2 _18528_ (.A(_02633_),
    .X(_02656_));
 sky130_fd_sc_hd__clkbuf_2 _18529_ (.A(_02635_),
    .X(_02657_));
 sky130_fd_sc_hd__or2_1 _18530_ (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .B(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__o211a_1 _18531_ (.A1(\rbzero.spi_registers.spi_buffer[10] ),
    .A2(_02656_),
    .B1(_02658_),
    .C1(_02654_),
    .X(_00616_));
 sky130_fd_sc_hd__or2_1 _18532_ (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .B(_02657_),
    .X(_02659_));
 sky130_fd_sc_hd__o211a_1 _18533_ (.A1(\rbzero.spi_registers.spi_buffer[11] ),
    .A2(_02656_),
    .B1(_02659_),
    .C1(_02654_),
    .X(_00617_));
 sky130_fd_sc_hd__or2_1 _18534_ (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .B(_02657_),
    .X(_02660_));
 sky130_fd_sc_hd__o211a_1 _18535_ (.A1(\rbzero.spi_registers.spi_buffer[12] ),
    .A2(_02656_),
    .B1(_02660_),
    .C1(_02654_),
    .X(_00618_));
 sky130_fd_sc_hd__or2_1 _18536_ (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .B(_02657_),
    .X(_02661_));
 sky130_fd_sc_hd__o211a_1 _18537_ (.A1(\rbzero.spi_registers.spi_buffer[13] ),
    .A2(_02656_),
    .B1(_02661_),
    .C1(_02654_),
    .X(_00619_));
 sky130_fd_sc_hd__or2_1 _18538_ (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .B(_02657_),
    .X(_02662_));
 sky130_fd_sc_hd__o211a_1 _18539_ (.A1(\rbzero.spi_registers.spi_buffer[14] ),
    .A2(_02656_),
    .B1(_02662_),
    .C1(_02654_),
    .X(_00620_));
 sky130_fd_sc_hd__or2_1 _18540_ (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .B(_02657_),
    .X(_02663_));
 sky130_fd_sc_hd__o211a_1 _18541_ (.A1(\rbzero.spi_registers.spi_buffer[15] ),
    .A2(_02656_),
    .B1(_02663_),
    .C1(_02654_),
    .X(_00621_));
 sky130_fd_sc_hd__or2_1 _18542_ (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .B(_02657_),
    .X(_02664_));
 sky130_fd_sc_hd__o211a_1 _18543_ (.A1(\rbzero.spi_registers.spi_buffer[16] ),
    .A2(_02656_),
    .B1(_02664_),
    .C1(_02654_),
    .X(_00622_));
 sky130_fd_sc_hd__or2_1 _18544_ (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .B(_02657_),
    .X(_02665_));
 sky130_fd_sc_hd__o211a_1 _18545_ (.A1(\rbzero.spi_registers.spi_buffer[17] ),
    .A2(_02656_),
    .B1(_02665_),
    .C1(_02654_),
    .X(_00623_));
 sky130_fd_sc_hd__or2_1 _18546_ (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .B(_02657_),
    .X(_02666_));
 sky130_fd_sc_hd__clkbuf_4 _18547_ (.A(_02653_),
    .X(_02667_));
 sky130_fd_sc_hd__o211a_1 _18548_ (.A1(\rbzero.spi_registers.spi_buffer[18] ),
    .A2(_02656_),
    .B1(_02666_),
    .C1(_02667_),
    .X(_00624_));
 sky130_fd_sc_hd__or2_1 _18549_ (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .B(_02657_),
    .X(_02668_));
 sky130_fd_sc_hd__o211a_1 _18550_ (.A1(\rbzero.spi_registers.spi_buffer[19] ),
    .A2(_02656_),
    .B1(_02668_),
    .C1(_02667_),
    .X(_00625_));
 sky130_fd_sc_hd__or2_1 _18551_ (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .B(_02635_),
    .X(_02669_));
 sky130_fd_sc_hd__o211a_1 _18552_ (.A1(\rbzero.spi_registers.spi_buffer[20] ),
    .A2(_02633_),
    .B1(_02669_),
    .C1(_02667_),
    .X(_00626_));
 sky130_fd_sc_hd__or2_1 _18553_ (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .B(_02635_),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_1 _18554_ (.A1(\rbzero.spi_registers.spi_buffer[21] ),
    .A2(_02633_),
    .B1(_02670_),
    .C1(_02667_),
    .X(_00627_));
 sky130_fd_sc_hd__or2_1 _18555_ (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .B(_02635_),
    .X(_02671_));
 sky130_fd_sc_hd__o211a_1 _18556_ (.A1(\rbzero.spi_registers.spi_buffer[22] ),
    .A2(_02633_),
    .B1(_02671_),
    .C1(_02667_),
    .X(_00628_));
 sky130_fd_sc_hd__or2_1 _18557_ (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .B(_02635_),
    .X(_02672_));
 sky130_fd_sc_hd__o211a_1 _18558_ (.A1(\rbzero.spi_registers.spi_buffer[23] ),
    .A2(_02633_),
    .B1(_02672_),
    .C1(_02667_),
    .X(_00629_));
 sky130_fd_sc_hd__and2_1 _18559_ (.A(net57),
    .B(_02371_),
    .X(_02673_));
 sky130_fd_sc_hd__clkbuf_1 _18560_ (.A(_02673_),
    .X(_00630_));
 sky130_fd_sc_hd__and2_1 _18561_ (.A(\rbzero.pov.sclk_buffer[0] ),
    .B(_09712_),
    .X(_02674_));
 sky130_fd_sc_hd__clkbuf_1 _18562_ (.A(_02674_),
    .X(_00631_));
 sky130_fd_sc_hd__and2_1 _18563_ (.A(\rbzero.pov.sclk_buffer[1] ),
    .B(_09712_),
    .X(_02675_));
 sky130_fd_sc_hd__clkbuf_1 _18564_ (.A(_02675_),
    .X(_00632_));
 sky130_fd_sc_hd__nor2_1 _18565_ (.A(_05001_),
    .B(_05014_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _18566_ (.A(_05186_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__or4b_2 _18567_ (.A(_05716_),
    .B(_05016_),
    .C(_02677_),
    .D_N(_05715_),
    .X(_02678_));
 sky130_fd_sc_hd__and4_1 _18568_ (.A(_05711_),
    .B(_04675_),
    .C(\gpout0.vpos[1] ),
    .D(\gpout0.vpos[0] ),
    .X(_02679_));
 sky130_fd_sc_hd__nand2_2 _18569_ (.A(_09708_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__nor2_1 _18570_ (.A(_02678_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__buf_4 _18571_ (.A(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__buf_4 _18572_ (.A(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__buf_2 _18573_ (.A(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__or2_4 _18574_ (.A(_02678_),
    .B(_02680_),
    .X(_02685_));
 sky130_fd_sc_hd__buf_4 _18575_ (.A(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__clkbuf_2 _18576_ (.A(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__or2_1 _18577_ (.A(\rbzero.spi_registers.buf_otherx[0] ),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__o211a_1 _18578_ (.A1(\rbzero.map_overlay.i_otherx[0] ),
    .A2(_02684_),
    .B1(_02688_),
    .C1(_02667_),
    .X(_00633_));
 sky130_fd_sc_hd__or2_1 _18579_ (.A(\rbzero.spi_registers.buf_otherx[1] ),
    .B(_02687_),
    .X(_02689_));
 sky130_fd_sc_hd__o211a_1 _18580_ (.A1(\rbzero.map_overlay.i_otherx[1] ),
    .A2(_02684_),
    .B1(_02689_),
    .C1(_02667_),
    .X(_00634_));
 sky130_fd_sc_hd__or2_1 _18581_ (.A(\rbzero.spi_registers.buf_otherx[2] ),
    .B(_02687_),
    .X(_02690_));
 sky130_fd_sc_hd__o211a_1 _18582_ (.A1(\rbzero.map_overlay.i_otherx[2] ),
    .A2(_02684_),
    .B1(_02690_),
    .C1(_02667_),
    .X(_00635_));
 sky130_fd_sc_hd__or2_1 _18583_ (.A(\rbzero.spi_registers.buf_otherx[3] ),
    .B(_02687_),
    .X(_02691_));
 sky130_fd_sc_hd__o211a_1 _18584_ (.A1(\rbzero.map_overlay.i_otherx[3] ),
    .A2(_02684_),
    .B1(_02691_),
    .C1(_02667_),
    .X(_00636_));
 sky130_fd_sc_hd__or2_1 _18585_ (.A(\rbzero.spi_registers.buf_otherx[4] ),
    .B(_02687_),
    .X(_02692_));
 sky130_fd_sc_hd__buf_4 _18586_ (.A(_08091_),
    .X(_02693_));
 sky130_fd_sc_hd__buf_2 _18587_ (.A(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__o211a_1 _18588_ (.A1(\rbzero.map_overlay.i_otherx[4] ),
    .A2(_02684_),
    .B1(_02692_),
    .C1(_02694_),
    .X(_00637_));
 sky130_fd_sc_hd__or2_1 _18589_ (.A(\rbzero.spi_registers.buf_othery[0] ),
    .B(_02687_),
    .X(_02695_));
 sky130_fd_sc_hd__o211a_1 _18590_ (.A1(\rbzero.map_overlay.i_othery[0] ),
    .A2(_02684_),
    .B1(_02695_),
    .C1(_02694_),
    .X(_00638_));
 sky130_fd_sc_hd__or2_1 _18591_ (.A(\rbzero.spi_registers.buf_othery[1] ),
    .B(_02687_),
    .X(_02696_));
 sky130_fd_sc_hd__o211a_1 _18592_ (.A1(\rbzero.map_overlay.i_othery[1] ),
    .A2(_02684_),
    .B1(_02696_),
    .C1(_02694_),
    .X(_00639_));
 sky130_fd_sc_hd__or2_1 _18593_ (.A(\rbzero.spi_registers.buf_othery[2] ),
    .B(_02687_),
    .X(_02697_));
 sky130_fd_sc_hd__o211a_1 _18594_ (.A1(\rbzero.map_overlay.i_othery[2] ),
    .A2(_02684_),
    .B1(_02697_),
    .C1(_02694_),
    .X(_00640_));
 sky130_fd_sc_hd__or2_1 _18595_ (.A(\rbzero.spi_registers.buf_othery[3] ),
    .B(_02687_),
    .X(_02698_));
 sky130_fd_sc_hd__o211a_1 _18596_ (.A1(\rbzero.map_overlay.i_othery[3] ),
    .A2(_02684_),
    .B1(_02698_),
    .C1(_02694_),
    .X(_00641_));
 sky130_fd_sc_hd__or2_1 _18597_ (.A(\rbzero.spi_registers.buf_othery[4] ),
    .B(_02687_),
    .X(_02699_));
 sky130_fd_sc_hd__o211a_1 _18598_ (.A1(\rbzero.map_overlay.i_othery[4] ),
    .A2(_02684_),
    .B1(_02699_),
    .C1(_02694_),
    .X(_00642_));
 sky130_fd_sc_hd__buf_2 _18599_ (.A(_02683_),
    .X(_02700_));
 sky130_fd_sc_hd__clkbuf_2 _18600_ (.A(_02686_),
    .X(_02701_));
 sky130_fd_sc_hd__or2_1 _18601_ (.A(\rbzero.spi_registers.buf_vinf ),
    .B(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__o211a_1 _18602_ (.A1(\rbzero.row_render.vinf ),
    .A2(_02700_),
    .B1(_02702_),
    .C1(_02694_),
    .X(_00643_));
 sky130_fd_sc_hd__or2_1 _18603_ (.A(\rbzero.spi_registers.buf_mapdx[0] ),
    .B(_02701_),
    .X(_02703_));
 sky130_fd_sc_hd__o211a_1 _18604_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_02700_),
    .B1(_02703_),
    .C1(_02694_),
    .X(_00644_));
 sky130_fd_sc_hd__or2_1 _18605_ (.A(\rbzero.spi_registers.buf_mapdx[1] ),
    .B(_02701_),
    .X(_02704_));
 sky130_fd_sc_hd__o211a_1 _18606_ (.A1(\rbzero.map_overlay.i_mapdx[1] ),
    .A2(_02700_),
    .B1(_02704_),
    .C1(_02694_),
    .X(_00645_));
 sky130_fd_sc_hd__or2_1 _18607_ (.A(\rbzero.spi_registers.buf_mapdx[2] ),
    .B(_02701_),
    .X(_02705_));
 sky130_fd_sc_hd__o211a_1 _18608_ (.A1(\rbzero.map_overlay.i_mapdx[2] ),
    .A2(_02700_),
    .B1(_02705_),
    .C1(_02694_),
    .X(_00646_));
 sky130_fd_sc_hd__or2_1 _18609_ (.A(\rbzero.spi_registers.buf_mapdx[3] ),
    .B(_02701_),
    .X(_02706_));
 sky130_fd_sc_hd__buf_2 _18610_ (.A(_02693_),
    .X(_02707_));
 sky130_fd_sc_hd__o211a_1 _18611_ (.A1(\rbzero.map_overlay.i_mapdx[3] ),
    .A2(_02700_),
    .B1(_02706_),
    .C1(_02707_),
    .X(_00647_));
 sky130_fd_sc_hd__or2_1 _18612_ (.A(\rbzero.spi_registers.buf_mapdx[4] ),
    .B(_02701_),
    .X(_02708_));
 sky130_fd_sc_hd__o211a_1 _18613_ (.A1(\rbzero.map_overlay.i_mapdx[4] ),
    .A2(_02700_),
    .B1(_02708_),
    .C1(_02707_),
    .X(_00648_));
 sky130_fd_sc_hd__or2_1 _18614_ (.A(\rbzero.spi_registers.buf_mapdx[5] ),
    .B(_02701_),
    .X(_02709_));
 sky130_fd_sc_hd__o211a_1 _18615_ (.A1(\rbzero.map_overlay.i_mapdx[5] ),
    .A2(_02700_),
    .B1(_02709_),
    .C1(_02707_),
    .X(_00649_));
 sky130_fd_sc_hd__or2_1 _18616_ (.A(\rbzero.spi_registers.buf_mapdy[0] ),
    .B(_02701_),
    .X(_02710_));
 sky130_fd_sc_hd__o211a_1 _18617_ (.A1(\rbzero.map_overlay.i_mapdy[0] ),
    .A2(_02700_),
    .B1(_02710_),
    .C1(_02707_),
    .X(_00650_));
 sky130_fd_sc_hd__or2_1 _18618_ (.A(\rbzero.spi_registers.buf_mapdy[1] ),
    .B(_02701_),
    .X(_02711_));
 sky130_fd_sc_hd__o211a_1 _18619_ (.A1(\rbzero.map_overlay.i_mapdy[1] ),
    .A2(_02700_),
    .B1(_02711_),
    .C1(_02707_),
    .X(_00651_));
 sky130_fd_sc_hd__or2_1 _18620_ (.A(\rbzero.spi_registers.buf_mapdy[2] ),
    .B(_02701_),
    .X(_02712_));
 sky130_fd_sc_hd__o211a_1 _18621_ (.A1(\rbzero.map_overlay.i_mapdy[2] ),
    .A2(_02700_),
    .B1(_02712_),
    .C1(_02707_),
    .X(_00652_));
 sky130_fd_sc_hd__clkbuf_4 _18622_ (.A(_02683_),
    .X(_02713_));
 sky130_fd_sc_hd__buf_2 _18623_ (.A(_02686_),
    .X(_02714_));
 sky130_fd_sc_hd__or2_1 _18624_ (.A(\rbzero.spi_registers.buf_mapdy[3] ),
    .B(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__o211a_1 _18625_ (.A1(\rbzero.map_overlay.i_mapdy[3] ),
    .A2(_02713_),
    .B1(_02715_),
    .C1(_02707_),
    .X(_00653_));
 sky130_fd_sc_hd__or2_1 _18626_ (.A(\rbzero.spi_registers.buf_mapdy[4] ),
    .B(_02714_),
    .X(_02716_));
 sky130_fd_sc_hd__o211a_1 _18627_ (.A1(\rbzero.map_overlay.i_mapdy[4] ),
    .A2(_02713_),
    .B1(_02716_),
    .C1(_02707_),
    .X(_00654_));
 sky130_fd_sc_hd__or2_1 _18628_ (.A(\rbzero.spi_registers.buf_mapdy[5] ),
    .B(_02714_),
    .X(_02717_));
 sky130_fd_sc_hd__o211a_1 _18629_ (.A1(\rbzero.map_overlay.i_mapdy[5] ),
    .A2(_02713_),
    .B1(_02717_),
    .C1(_02707_),
    .X(_00655_));
 sky130_fd_sc_hd__or2_1 _18630_ (.A(\rbzero.spi_registers.buf_mapdxw[0] ),
    .B(_02714_),
    .X(_02718_));
 sky130_fd_sc_hd__o211a_1 _18631_ (.A1(\rbzero.mapdxw[0] ),
    .A2(_02713_),
    .B1(_02718_),
    .C1(_02707_),
    .X(_00656_));
 sky130_fd_sc_hd__or2_1 _18632_ (.A(\rbzero.spi_registers.buf_mapdxw[1] ),
    .B(_02714_),
    .X(_02719_));
 sky130_fd_sc_hd__clkbuf_4 _18633_ (.A(_02693_),
    .X(_02720_));
 sky130_fd_sc_hd__o211a_1 _18634_ (.A1(\rbzero.mapdxw[1] ),
    .A2(_02713_),
    .B1(_02719_),
    .C1(_02720_),
    .X(_00657_));
 sky130_fd_sc_hd__or2_1 _18635_ (.A(\rbzero.spi_registers.buf_mapdyw[0] ),
    .B(_02714_),
    .X(_02721_));
 sky130_fd_sc_hd__o211a_1 _18636_ (.A1(\rbzero.mapdyw[0] ),
    .A2(_02713_),
    .B1(_02721_),
    .C1(_02720_),
    .X(_00658_));
 sky130_fd_sc_hd__or2_1 _18637_ (.A(\rbzero.spi_registers.buf_mapdyw[1] ),
    .B(_02714_),
    .X(_02722_));
 sky130_fd_sc_hd__o211a_1 _18638_ (.A1(\rbzero.mapdyw[1] ),
    .A2(_02713_),
    .B1(_02722_),
    .C1(_02720_),
    .X(_00659_));
 sky130_fd_sc_hd__or2_1 _18639_ (.A(\rbzero.spi_registers.buf_leak[0] ),
    .B(_02714_),
    .X(_02723_));
 sky130_fd_sc_hd__o211a_1 _18640_ (.A1(\rbzero.floor_leak[0] ),
    .A2(_02713_),
    .B1(_02723_),
    .C1(_02720_),
    .X(_00660_));
 sky130_fd_sc_hd__or2_1 _18641_ (.A(\rbzero.spi_registers.buf_leak[1] ),
    .B(_02714_),
    .X(_02724_));
 sky130_fd_sc_hd__o211a_1 _18642_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_02713_),
    .B1(_02724_),
    .C1(_02720_),
    .X(_00661_));
 sky130_fd_sc_hd__or2_1 _18643_ (.A(\rbzero.spi_registers.buf_leak[2] ),
    .B(_02714_),
    .X(_02725_));
 sky130_fd_sc_hd__o211a_1 _18644_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_02713_),
    .B1(_02725_),
    .C1(_02720_),
    .X(_00662_));
 sky130_fd_sc_hd__buf_2 _18645_ (.A(_02683_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_2 _18646_ (.A(_02686_),
    .X(_02727_));
 sky130_fd_sc_hd__or2_1 _18647_ (.A(\rbzero.spi_registers.buf_leak[3] ),
    .B(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__o211a_1 _18648_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_02726_),
    .B1(_02728_),
    .C1(_02720_),
    .X(_00663_));
 sky130_fd_sc_hd__or2_1 _18649_ (.A(\rbzero.spi_registers.buf_leak[4] ),
    .B(_02727_),
    .X(_02729_));
 sky130_fd_sc_hd__o211a_1 _18650_ (.A1(\rbzero.floor_leak[4] ),
    .A2(_02726_),
    .B1(_02729_),
    .C1(_02720_),
    .X(_00664_));
 sky130_fd_sc_hd__or2_1 _18651_ (.A(\rbzero.spi_registers.buf_leak[5] ),
    .B(_02727_),
    .X(_02730_));
 sky130_fd_sc_hd__o211a_1 _18652_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_02726_),
    .B1(_02730_),
    .C1(_02720_),
    .X(_00665_));
 sky130_fd_sc_hd__buf_4 _18653_ (.A(_04094_),
    .X(_02731_));
 sky130_fd_sc_hd__clkbuf_8 _18654_ (.A(_02685_),
    .X(_02732_));
 sky130_fd_sc_hd__mux2_1 _18655_ (.A0(\rbzero.spi_registers.buf_sky[0] ),
    .A1(\rbzero.color_sky[0] ),
    .S(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__or2_1 _18656_ (.A(_02731_),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_1 _18657_ (.A(_02734_),
    .X(_00666_));
 sky130_fd_sc_hd__or2_1 _18658_ (.A(\rbzero.spi_registers.buf_sky[1] ),
    .B(_02727_),
    .X(_02735_));
 sky130_fd_sc_hd__o211a_1 _18659_ (.A1(\rbzero.color_sky[1] ),
    .A2(_02726_),
    .B1(_02735_),
    .C1(_02720_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _18660_ (.A0(\rbzero.spi_registers.buf_sky[2] ),
    .A1(\rbzero.color_sky[2] ),
    .S(_02732_),
    .X(_02736_));
 sky130_fd_sc_hd__or2_1 _18661_ (.A(_02731_),
    .B(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__clkbuf_1 _18662_ (.A(_02737_),
    .X(_00668_));
 sky130_fd_sc_hd__or2_1 _18663_ (.A(\rbzero.spi_registers.buf_sky[3] ),
    .B(_02727_),
    .X(_02738_));
 sky130_fd_sc_hd__clkbuf_4 _18664_ (.A(_02693_),
    .X(_02739_));
 sky130_fd_sc_hd__o211a_1 _18665_ (.A1(\rbzero.color_sky[3] ),
    .A2(_02726_),
    .B1(_02738_),
    .C1(_02739_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _18666_ (.A0(\rbzero.spi_registers.buf_sky[4] ),
    .A1(\rbzero.color_sky[4] ),
    .S(_02732_),
    .X(_02740_));
 sky130_fd_sc_hd__or2_1 _18667_ (.A(_02731_),
    .B(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__clkbuf_1 _18668_ (.A(_02741_),
    .X(_00670_));
 sky130_fd_sc_hd__or2_1 _18669_ (.A(\rbzero.spi_registers.buf_sky[5] ),
    .B(_02727_),
    .X(_02742_));
 sky130_fd_sc_hd__o211a_1 _18670_ (.A1(\rbzero.color_sky[5] ),
    .A2(_02726_),
    .B1(_02742_),
    .C1(_02739_),
    .X(_00671_));
 sky130_fd_sc_hd__or2_1 _18671_ (.A(\rbzero.spi_registers.buf_floor[0] ),
    .B(_02727_),
    .X(_02743_));
 sky130_fd_sc_hd__o211a_1 _18672_ (.A1(\rbzero.color_floor[0] ),
    .A2(_02726_),
    .B1(_02743_),
    .C1(_02739_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _18673_ (.A0(\rbzero.spi_registers.buf_floor[1] ),
    .A1(\rbzero.color_floor[1] ),
    .S(_02732_),
    .X(_02744_));
 sky130_fd_sc_hd__or2_1 _18674_ (.A(_02731_),
    .B(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__clkbuf_1 _18675_ (.A(_02745_),
    .X(_00673_));
 sky130_fd_sc_hd__or2_1 _18676_ (.A(\rbzero.spi_registers.buf_floor[2] ),
    .B(_02727_),
    .X(_02746_));
 sky130_fd_sc_hd__o211a_1 _18677_ (.A1(\rbzero.color_floor[2] ),
    .A2(_02726_),
    .B1(_02746_),
    .C1(_02739_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _18678_ (.A0(\rbzero.spi_registers.buf_floor[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_02685_),
    .X(_02747_));
 sky130_fd_sc_hd__or2_1 _18679_ (.A(_02731_),
    .B(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__clkbuf_1 _18680_ (.A(_02748_),
    .X(_00675_));
 sky130_fd_sc_hd__or2_1 _18681_ (.A(\rbzero.spi_registers.buf_floor[4] ),
    .B(_02727_),
    .X(_02749_));
 sky130_fd_sc_hd__o211a_1 _18682_ (.A1(\rbzero.color_floor[4] ),
    .A2(_02726_),
    .B1(_02749_),
    .C1(_02739_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _18683_ (.A0(\rbzero.spi_registers.buf_floor[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_02685_),
    .X(_02750_));
 sky130_fd_sc_hd__or2_1 _18684_ (.A(_02731_),
    .B(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__clkbuf_1 _18685_ (.A(_02751_),
    .X(_00677_));
 sky130_fd_sc_hd__or2_1 _18686_ (.A(\rbzero.spi_registers.buf_vshift[0] ),
    .B(_02727_),
    .X(_02752_));
 sky130_fd_sc_hd__o211a_1 _18687_ (.A1(\rbzero.spi_registers.vshift[0] ),
    .A2(_02726_),
    .B1(_02752_),
    .C1(_02739_),
    .X(_00678_));
 sky130_fd_sc_hd__buf_2 _18688_ (.A(_02683_),
    .X(_02753_));
 sky130_fd_sc_hd__clkbuf_2 _18689_ (.A(_02686_),
    .X(_02754_));
 sky130_fd_sc_hd__or2_1 _18690_ (.A(\rbzero.spi_registers.buf_vshift[1] ),
    .B(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__o211a_1 _18691_ (.A1(\rbzero.spi_registers.vshift[1] ),
    .A2(_02753_),
    .B1(_02755_),
    .C1(_02739_),
    .X(_00679_));
 sky130_fd_sc_hd__or2_1 _18692_ (.A(\rbzero.spi_registers.buf_vshift[2] ),
    .B(_02754_),
    .X(_02756_));
 sky130_fd_sc_hd__o211a_1 _18693_ (.A1(\rbzero.spi_registers.vshift[2] ),
    .A2(_02753_),
    .B1(_02756_),
    .C1(_02739_),
    .X(_00680_));
 sky130_fd_sc_hd__or2_1 _18694_ (.A(\rbzero.spi_registers.buf_vshift[3] ),
    .B(_02754_),
    .X(_02757_));
 sky130_fd_sc_hd__o211a_1 _18695_ (.A1(\rbzero.spi_registers.vshift[3] ),
    .A2(_02753_),
    .B1(_02757_),
    .C1(_02739_),
    .X(_00681_));
 sky130_fd_sc_hd__or2_1 _18696_ (.A(\rbzero.spi_registers.buf_vshift[4] ),
    .B(_02754_),
    .X(_02758_));
 sky130_fd_sc_hd__o211a_1 _18697_ (.A1(\rbzero.spi_registers.vshift[4] ),
    .A2(_02753_),
    .B1(_02758_),
    .C1(_02739_),
    .X(_00682_));
 sky130_fd_sc_hd__or2_1 _18698_ (.A(\rbzero.spi_registers.buf_vshift[5] ),
    .B(_02754_),
    .X(_02759_));
 sky130_fd_sc_hd__buf_2 _18699_ (.A(_02693_),
    .X(_02760_));
 sky130_fd_sc_hd__o211a_1 _18700_ (.A1(\rbzero.spi_registers.vshift[5] ),
    .A2(_02753_),
    .B1(_02759_),
    .C1(_02760_),
    .X(_00683_));
 sky130_fd_sc_hd__or2_1 _18701_ (.A(\rbzero.spi_registers.buf_texadd0[0] ),
    .B(_02754_),
    .X(_02761_));
 sky130_fd_sc_hd__o211a_1 _18702_ (.A1(\rbzero.spi_registers.texadd0[0] ),
    .A2(_02753_),
    .B1(_02761_),
    .C1(_02760_),
    .X(_00684_));
 sky130_fd_sc_hd__or2_1 _18703_ (.A(\rbzero.spi_registers.buf_texadd0[1] ),
    .B(_02754_),
    .X(_02762_));
 sky130_fd_sc_hd__o211a_1 _18704_ (.A1(\rbzero.spi_registers.texadd0[1] ),
    .A2(_02753_),
    .B1(_02762_),
    .C1(_02760_),
    .X(_00685_));
 sky130_fd_sc_hd__or2_1 _18705_ (.A(\rbzero.spi_registers.buf_texadd0[2] ),
    .B(_02754_),
    .X(_02763_));
 sky130_fd_sc_hd__o211a_1 _18706_ (.A1(\rbzero.spi_registers.texadd0[2] ),
    .A2(_02753_),
    .B1(_02763_),
    .C1(_02760_),
    .X(_00686_));
 sky130_fd_sc_hd__or2_1 _18707_ (.A(\rbzero.spi_registers.buf_texadd0[3] ),
    .B(_02754_),
    .X(_02764_));
 sky130_fd_sc_hd__o211a_1 _18708_ (.A1(\rbzero.spi_registers.texadd0[3] ),
    .A2(_02753_),
    .B1(_02764_),
    .C1(_02760_),
    .X(_00687_));
 sky130_fd_sc_hd__or2_1 _18709_ (.A(\rbzero.spi_registers.buf_texadd0[4] ),
    .B(_02754_),
    .X(_02765_));
 sky130_fd_sc_hd__o211a_1 _18710_ (.A1(\rbzero.spi_registers.texadd0[4] ),
    .A2(_02753_),
    .B1(_02765_),
    .C1(_02760_),
    .X(_00688_));
 sky130_fd_sc_hd__clkbuf_4 _18711_ (.A(_02683_),
    .X(_02766_));
 sky130_fd_sc_hd__buf_2 _18712_ (.A(_02686_),
    .X(_02767_));
 sky130_fd_sc_hd__or2_1 _18713_ (.A(\rbzero.spi_registers.buf_texadd0[5] ),
    .B(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__o211a_1 _18714_ (.A1(\rbzero.spi_registers.texadd0[5] ),
    .A2(_02766_),
    .B1(_02768_),
    .C1(_02760_),
    .X(_00689_));
 sky130_fd_sc_hd__or2_1 _18715_ (.A(\rbzero.spi_registers.buf_texadd0[6] ),
    .B(_02767_),
    .X(_02769_));
 sky130_fd_sc_hd__o211a_1 _18716_ (.A1(\rbzero.spi_registers.texadd0[6] ),
    .A2(_02766_),
    .B1(_02769_),
    .C1(_02760_),
    .X(_00690_));
 sky130_fd_sc_hd__or2_1 _18717_ (.A(\rbzero.spi_registers.buf_texadd0[7] ),
    .B(_02767_),
    .X(_02770_));
 sky130_fd_sc_hd__o211a_1 _18718_ (.A1(\rbzero.spi_registers.texadd0[7] ),
    .A2(_02766_),
    .B1(_02770_),
    .C1(_02760_),
    .X(_00691_));
 sky130_fd_sc_hd__or2_1 _18719_ (.A(\rbzero.spi_registers.buf_texadd0[8] ),
    .B(_02767_),
    .X(_02771_));
 sky130_fd_sc_hd__o211a_1 _18720_ (.A1(\rbzero.spi_registers.texadd0[8] ),
    .A2(_02766_),
    .B1(_02771_),
    .C1(_02760_),
    .X(_00692_));
 sky130_fd_sc_hd__or2_1 _18721_ (.A(\rbzero.spi_registers.buf_texadd0[9] ),
    .B(_02767_),
    .X(_02772_));
 sky130_fd_sc_hd__buf_2 _18722_ (.A(_02693_),
    .X(_02773_));
 sky130_fd_sc_hd__o211a_1 _18723_ (.A1(\rbzero.spi_registers.texadd0[9] ),
    .A2(_02766_),
    .B1(_02772_),
    .C1(_02773_),
    .X(_00693_));
 sky130_fd_sc_hd__or2_1 _18724_ (.A(\rbzero.spi_registers.buf_texadd0[10] ),
    .B(_02767_),
    .X(_02774_));
 sky130_fd_sc_hd__o211a_1 _18725_ (.A1(\rbzero.spi_registers.texadd0[10] ),
    .A2(_02766_),
    .B1(_02774_),
    .C1(_02773_),
    .X(_00694_));
 sky130_fd_sc_hd__or2_1 _18726_ (.A(\rbzero.spi_registers.buf_texadd0[11] ),
    .B(_02767_),
    .X(_02775_));
 sky130_fd_sc_hd__o211a_1 _18727_ (.A1(\rbzero.spi_registers.texadd0[11] ),
    .A2(_02766_),
    .B1(_02775_),
    .C1(_02773_),
    .X(_00695_));
 sky130_fd_sc_hd__or2_1 _18728_ (.A(\rbzero.spi_registers.buf_texadd0[12] ),
    .B(_02767_),
    .X(_02776_));
 sky130_fd_sc_hd__o211a_1 _18729_ (.A1(\rbzero.spi_registers.texadd0[12] ),
    .A2(_02766_),
    .B1(_02776_),
    .C1(_02773_),
    .X(_00696_));
 sky130_fd_sc_hd__or2_1 _18730_ (.A(\rbzero.spi_registers.buf_texadd0[13] ),
    .B(_02767_),
    .X(_02777_));
 sky130_fd_sc_hd__o211a_1 _18731_ (.A1(\rbzero.spi_registers.texadd0[13] ),
    .A2(_02766_),
    .B1(_02777_),
    .C1(_02773_),
    .X(_00697_));
 sky130_fd_sc_hd__or2_1 _18732_ (.A(\rbzero.spi_registers.buf_texadd0[14] ),
    .B(_02767_),
    .X(_02778_));
 sky130_fd_sc_hd__o211a_1 _18733_ (.A1(\rbzero.spi_registers.texadd0[14] ),
    .A2(_02766_),
    .B1(_02778_),
    .C1(_02773_),
    .X(_00698_));
 sky130_fd_sc_hd__clkbuf_4 _18734_ (.A(_02683_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_2 _18735_ (.A(_02686_),
    .X(_02780_));
 sky130_fd_sc_hd__or2_1 _18736_ (.A(\rbzero.spi_registers.buf_texadd0[15] ),
    .B(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__o211a_1 _18737_ (.A1(\rbzero.spi_registers.texadd0[15] ),
    .A2(_02779_),
    .B1(_02781_),
    .C1(_02773_),
    .X(_00699_));
 sky130_fd_sc_hd__or2_1 _18738_ (.A(\rbzero.spi_registers.buf_texadd0[16] ),
    .B(_02780_),
    .X(_02782_));
 sky130_fd_sc_hd__o211a_1 _18739_ (.A1(\rbzero.spi_registers.texadd0[16] ),
    .A2(_02779_),
    .B1(_02782_),
    .C1(_02773_),
    .X(_00700_));
 sky130_fd_sc_hd__or2_1 _18740_ (.A(\rbzero.spi_registers.buf_texadd0[17] ),
    .B(_02780_),
    .X(_02783_));
 sky130_fd_sc_hd__o211a_1 _18741_ (.A1(\rbzero.spi_registers.texadd0[17] ),
    .A2(_02779_),
    .B1(_02783_),
    .C1(_02773_),
    .X(_00701_));
 sky130_fd_sc_hd__or2_1 _18742_ (.A(\rbzero.spi_registers.buf_texadd0[18] ),
    .B(_02780_),
    .X(_02784_));
 sky130_fd_sc_hd__o211a_1 _18743_ (.A1(\rbzero.spi_registers.texadd0[18] ),
    .A2(_02779_),
    .B1(_02784_),
    .C1(_02773_),
    .X(_00702_));
 sky130_fd_sc_hd__or2_1 _18744_ (.A(\rbzero.spi_registers.buf_texadd0[19] ),
    .B(_02780_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_4 _18745_ (.A(_02693_),
    .X(_02786_));
 sky130_fd_sc_hd__o211a_1 _18746_ (.A1(\rbzero.spi_registers.texadd0[19] ),
    .A2(_02779_),
    .B1(_02785_),
    .C1(_02786_),
    .X(_00703_));
 sky130_fd_sc_hd__or2_1 _18747_ (.A(\rbzero.spi_registers.buf_texadd0[20] ),
    .B(_02780_),
    .X(_02787_));
 sky130_fd_sc_hd__o211a_1 _18748_ (.A1(\rbzero.spi_registers.texadd0[20] ),
    .A2(_02779_),
    .B1(_02787_),
    .C1(_02786_),
    .X(_00704_));
 sky130_fd_sc_hd__or2_1 _18749_ (.A(\rbzero.spi_registers.buf_texadd0[21] ),
    .B(_02780_),
    .X(_02788_));
 sky130_fd_sc_hd__o211a_1 _18750_ (.A1(\rbzero.spi_registers.texadd0[21] ),
    .A2(_02779_),
    .B1(_02788_),
    .C1(_02786_),
    .X(_00705_));
 sky130_fd_sc_hd__or2_1 _18751_ (.A(\rbzero.spi_registers.buf_texadd0[22] ),
    .B(_02780_),
    .X(_02789_));
 sky130_fd_sc_hd__o211a_1 _18752_ (.A1(\rbzero.spi_registers.texadd0[22] ),
    .A2(_02779_),
    .B1(_02789_),
    .C1(_02786_),
    .X(_00706_));
 sky130_fd_sc_hd__or2_1 _18753_ (.A(\rbzero.spi_registers.buf_texadd0[23] ),
    .B(_02780_),
    .X(_02790_));
 sky130_fd_sc_hd__o211a_1 _18754_ (.A1(\rbzero.spi_registers.texadd0[23] ),
    .A2(_02779_),
    .B1(_02790_),
    .C1(_02786_),
    .X(_00707_));
 sky130_fd_sc_hd__or2_1 _18755_ (.A(\rbzero.spi_registers.buf_texadd1[0] ),
    .B(_02780_),
    .X(_02791_));
 sky130_fd_sc_hd__o211a_1 _18756_ (.A1(\rbzero.spi_registers.texadd1[0] ),
    .A2(_02779_),
    .B1(_02791_),
    .C1(_02786_),
    .X(_00708_));
 sky130_fd_sc_hd__buf_2 _18757_ (.A(_02683_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_2 _18758_ (.A(_02686_),
    .X(_02793_));
 sky130_fd_sc_hd__or2_1 _18759_ (.A(\rbzero.spi_registers.buf_texadd1[1] ),
    .B(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__o211a_1 _18760_ (.A1(\rbzero.spi_registers.texadd1[1] ),
    .A2(_02792_),
    .B1(_02794_),
    .C1(_02786_),
    .X(_00709_));
 sky130_fd_sc_hd__or2_1 _18761_ (.A(\rbzero.spi_registers.buf_texadd1[2] ),
    .B(_02793_),
    .X(_02795_));
 sky130_fd_sc_hd__o211a_1 _18762_ (.A1(\rbzero.spi_registers.texadd1[2] ),
    .A2(_02792_),
    .B1(_02795_),
    .C1(_02786_),
    .X(_00710_));
 sky130_fd_sc_hd__or2_1 _18763_ (.A(\rbzero.spi_registers.buf_texadd1[3] ),
    .B(_02793_),
    .X(_02796_));
 sky130_fd_sc_hd__o211a_1 _18764_ (.A1(\rbzero.spi_registers.texadd1[3] ),
    .A2(_02792_),
    .B1(_02796_),
    .C1(_02786_),
    .X(_00711_));
 sky130_fd_sc_hd__or2_1 _18765_ (.A(\rbzero.spi_registers.buf_texadd1[4] ),
    .B(_02793_),
    .X(_02797_));
 sky130_fd_sc_hd__o211a_1 _18766_ (.A1(\rbzero.spi_registers.texadd1[4] ),
    .A2(_02792_),
    .B1(_02797_),
    .C1(_02786_),
    .X(_00712_));
 sky130_fd_sc_hd__or2_1 _18767_ (.A(\rbzero.spi_registers.buf_texadd1[5] ),
    .B(_02793_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_4 _18768_ (.A(_02693_),
    .X(_02799_));
 sky130_fd_sc_hd__o211a_1 _18769_ (.A1(\rbzero.spi_registers.texadd1[5] ),
    .A2(_02792_),
    .B1(_02798_),
    .C1(_02799_),
    .X(_00713_));
 sky130_fd_sc_hd__or2_1 _18770_ (.A(\rbzero.spi_registers.buf_texadd1[6] ),
    .B(_02793_),
    .X(_02800_));
 sky130_fd_sc_hd__o211a_1 _18771_ (.A1(\rbzero.spi_registers.texadd1[6] ),
    .A2(_02792_),
    .B1(_02800_),
    .C1(_02799_),
    .X(_00714_));
 sky130_fd_sc_hd__or2_1 _18772_ (.A(\rbzero.spi_registers.buf_texadd1[7] ),
    .B(_02793_),
    .X(_02801_));
 sky130_fd_sc_hd__o211a_1 _18773_ (.A1(\rbzero.spi_registers.texadd1[7] ),
    .A2(_02792_),
    .B1(_02801_),
    .C1(_02799_),
    .X(_00715_));
 sky130_fd_sc_hd__or2_1 _18774_ (.A(\rbzero.spi_registers.buf_texadd1[8] ),
    .B(_02793_),
    .X(_02802_));
 sky130_fd_sc_hd__o211a_1 _18775_ (.A1(\rbzero.spi_registers.texadd1[8] ),
    .A2(_02792_),
    .B1(_02802_),
    .C1(_02799_),
    .X(_00716_));
 sky130_fd_sc_hd__or2_1 _18776_ (.A(\rbzero.spi_registers.buf_texadd1[9] ),
    .B(_02793_),
    .X(_02803_));
 sky130_fd_sc_hd__o211a_1 _18777_ (.A1(\rbzero.spi_registers.texadd1[9] ),
    .A2(_02792_),
    .B1(_02803_),
    .C1(_02799_),
    .X(_00717_));
 sky130_fd_sc_hd__or2_1 _18778_ (.A(\rbzero.spi_registers.buf_texadd1[10] ),
    .B(_02793_),
    .X(_02804_));
 sky130_fd_sc_hd__o211a_1 _18779_ (.A1(\rbzero.spi_registers.texadd1[10] ),
    .A2(_02792_),
    .B1(_02804_),
    .C1(_02799_),
    .X(_00718_));
 sky130_fd_sc_hd__clkbuf_4 _18780_ (.A(_02683_),
    .X(_02805_));
 sky130_fd_sc_hd__buf_2 _18781_ (.A(_02686_),
    .X(_02806_));
 sky130_fd_sc_hd__or2_1 _18782_ (.A(\rbzero.spi_registers.buf_texadd1[11] ),
    .B(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__o211a_1 _18783_ (.A1(\rbzero.spi_registers.texadd1[11] ),
    .A2(_02805_),
    .B1(_02807_),
    .C1(_02799_),
    .X(_00719_));
 sky130_fd_sc_hd__or2_1 _18784_ (.A(\rbzero.spi_registers.buf_texadd1[12] ),
    .B(_02806_),
    .X(_02808_));
 sky130_fd_sc_hd__o211a_1 _18785_ (.A1(\rbzero.spi_registers.texadd1[12] ),
    .A2(_02805_),
    .B1(_02808_),
    .C1(_02799_),
    .X(_00720_));
 sky130_fd_sc_hd__or2_1 _18786_ (.A(\rbzero.spi_registers.buf_texadd1[13] ),
    .B(_02806_),
    .X(_02809_));
 sky130_fd_sc_hd__o211a_1 _18787_ (.A1(\rbzero.spi_registers.texadd1[13] ),
    .A2(_02805_),
    .B1(_02809_),
    .C1(_02799_),
    .X(_00721_));
 sky130_fd_sc_hd__or2_1 _18788_ (.A(\rbzero.spi_registers.buf_texadd1[14] ),
    .B(_02806_),
    .X(_02810_));
 sky130_fd_sc_hd__o211a_1 _18789_ (.A1(\rbzero.spi_registers.texadd1[14] ),
    .A2(_02805_),
    .B1(_02810_),
    .C1(_02799_),
    .X(_00722_));
 sky130_fd_sc_hd__or2_1 _18790_ (.A(\rbzero.spi_registers.buf_texadd1[15] ),
    .B(_02806_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_4 _18791_ (.A(_02693_),
    .X(_02812_));
 sky130_fd_sc_hd__o211a_1 _18792_ (.A1(\rbzero.spi_registers.texadd1[15] ),
    .A2(_02805_),
    .B1(_02811_),
    .C1(_02812_),
    .X(_00723_));
 sky130_fd_sc_hd__or2_1 _18793_ (.A(\rbzero.spi_registers.buf_texadd1[16] ),
    .B(_02806_),
    .X(_02813_));
 sky130_fd_sc_hd__o211a_1 _18794_ (.A1(\rbzero.spi_registers.texadd1[16] ),
    .A2(_02805_),
    .B1(_02813_),
    .C1(_02812_),
    .X(_00724_));
 sky130_fd_sc_hd__or2_1 _18795_ (.A(\rbzero.spi_registers.buf_texadd1[17] ),
    .B(_02806_),
    .X(_02814_));
 sky130_fd_sc_hd__o211a_1 _18796_ (.A1(\rbzero.spi_registers.texadd1[17] ),
    .A2(_02805_),
    .B1(_02814_),
    .C1(_02812_),
    .X(_00725_));
 sky130_fd_sc_hd__or2_1 _18797_ (.A(\rbzero.spi_registers.buf_texadd1[18] ),
    .B(_02806_),
    .X(_02815_));
 sky130_fd_sc_hd__o211a_1 _18798_ (.A1(\rbzero.spi_registers.texadd1[18] ),
    .A2(_02805_),
    .B1(_02815_),
    .C1(_02812_),
    .X(_00726_));
 sky130_fd_sc_hd__or2_1 _18799_ (.A(\rbzero.spi_registers.buf_texadd1[19] ),
    .B(_02806_),
    .X(_02816_));
 sky130_fd_sc_hd__o211a_1 _18800_ (.A1(\rbzero.spi_registers.texadd1[19] ),
    .A2(_02805_),
    .B1(_02816_),
    .C1(_02812_),
    .X(_00727_));
 sky130_fd_sc_hd__or2_1 _18801_ (.A(\rbzero.spi_registers.buf_texadd1[20] ),
    .B(_02806_),
    .X(_02817_));
 sky130_fd_sc_hd__o211a_1 _18802_ (.A1(\rbzero.spi_registers.texadd1[20] ),
    .A2(_02805_),
    .B1(_02817_),
    .C1(_02812_),
    .X(_00728_));
 sky130_fd_sc_hd__clkbuf_4 _18803_ (.A(_02682_),
    .X(_02818_));
 sky130_fd_sc_hd__buf_2 _18804_ (.A(_02732_),
    .X(_02819_));
 sky130_fd_sc_hd__or2_1 _18805_ (.A(\rbzero.spi_registers.buf_texadd1[21] ),
    .B(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__o211a_1 _18806_ (.A1(\rbzero.spi_registers.texadd1[21] ),
    .A2(_02818_),
    .B1(_02820_),
    .C1(_02812_),
    .X(_00729_));
 sky130_fd_sc_hd__or2_1 _18807_ (.A(\rbzero.spi_registers.buf_texadd1[22] ),
    .B(_02819_),
    .X(_02821_));
 sky130_fd_sc_hd__o211a_1 _18808_ (.A1(\rbzero.spi_registers.texadd1[22] ),
    .A2(_02818_),
    .B1(_02821_),
    .C1(_02812_),
    .X(_00730_));
 sky130_fd_sc_hd__or2_1 _18809_ (.A(\rbzero.spi_registers.buf_texadd1[23] ),
    .B(_02819_),
    .X(_02822_));
 sky130_fd_sc_hd__o211a_1 _18810_ (.A1(\rbzero.spi_registers.texadd1[23] ),
    .A2(_02818_),
    .B1(_02822_),
    .C1(_02812_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_1 _18811_ (.A(\rbzero.spi_registers.buf_texadd2[0] ),
    .B(_02819_),
    .X(_02823_));
 sky130_fd_sc_hd__o211a_1 _18812_ (.A1(\rbzero.spi_registers.texadd2[0] ),
    .A2(_02818_),
    .B1(_02823_),
    .C1(_02812_),
    .X(_00732_));
 sky130_fd_sc_hd__or2_1 _18813_ (.A(\rbzero.spi_registers.buf_texadd2[1] ),
    .B(_02819_),
    .X(_02824_));
 sky130_fd_sc_hd__clkbuf_4 _18814_ (.A(_02693_),
    .X(_02825_));
 sky130_fd_sc_hd__o211a_1 _18815_ (.A1(\rbzero.spi_registers.texadd2[1] ),
    .A2(_02818_),
    .B1(_02824_),
    .C1(_02825_),
    .X(_00733_));
 sky130_fd_sc_hd__or2_1 _18816_ (.A(\rbzero.spi_registers.buf_texadd2[2] ),
    .B(_02819_),
    .X(_02826_));
 sky130_fd_sc_hd__o211a_1 _18817_ (.A1(\rbzero.spi_registers.texadd2[2] ),
    .A2(_02818_),
    .B1(_02826_),
    .C1(_02825_),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _18818_ (.A(\rbzero.spi_registers.buf_texadd2[3] ),
    .B(_02819_),
    .X(_02827_));
 sky130_fd_sc_hd__o211a_1 _18819_ (.A1(\rbzero.spi_registers.texadd2[3] ),
    .A2(_02818_),
    .B1(_02827_),
    .C1(_02825_),
    .X(_00735_));
 sky130_fd_sc_hd__or2_1 _18820_ (.A(\rbzero.spi_registers.buf_texadd2[4] ),
    .B(_02819_),
    .X(_02828_));
 sky130_fd_sc_hd__o211a_1 _18821_ (.A1(\rbzero.spi_registers.texadd2[4] ),
    .A2(_02818_),
    .B1(_02828_),
    .C1(_02825_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _18822_ (.A(\rbzero.spi_registers.buf_texadd2[5] ),
    .B(_02819_),
    .X(_02829_));
 sky130_fd_sc_hd__o211a_1 _18823_ (.A1(\rbzero.spi_registers.texadd2[5] ),
    .A2(_02818_),
    .B1(_02829_),
    .C1(_02825_),
    .X(_00737_));
 sky130_fd_sc_hd__or2_1 _18824_ (.A(\rbzero.spi_registers.buf_texadd2[6] ),
    .B(_02819_),
    .X(_02830_));
 sky130_fd_sc_hd__o211a_1 _18825_ (.A1(\rbzero.spi_registers.texadd2[6] ),
    .A2(_02818_),
    .B1(_02830_),
    .C1(_02825_),
    .X(_00738_));
 sky130_fd_sc_hd__clkbuf_4 _18826_ (.A(_02682_),
    .X(_02831_));
 sky130_fd_sc_hd__buf_2 _18827_ (.A(_02732_),
    .X(_02832_));
 sky130_fd_sc_hd__or2_1 _18828_ (.A(\rbzero.spi_registers.buf_texadd2[7] ),
    .B(_02832_),
    .X(_02833_));
 sky130_fd_sc_hd__o211a_1 _18829_ (.A1(\rbzero.spi_registers.texadd2[7] ),
    .A2(_02831_),
    .B1(_02833_),
    .C1(_02825_),
    .X(_00739_));
 sky130_fd_sc_hd__or2_1 _18830_ (.A(\rbzero.spi_registers.buf_texadd2[8] ),
    .B(_02832_),
    .X(_02834_));
 sky130_fd_sc_hd__o211a_1 _18831_ (.A1(\rbzero.spi_registers.texadd2[8] ),
    .A2(_02831_),
    .B1(_02834_),
    .C1(_02825_),
    .X(_00740_));
 sky130_fd_sc_hd__or2_1 _18832_ (.A(\rbzero.spi_registers.buf_texadd2[9] ),
    .B(_02832_),
    .X(_02835_));
 sky130_fd_sc_hd__o211a_1 _18833_ (.A1(\rbzero.spi_registers.texadd2[9] ),
    .A2(_02831_),
    .B1(_02835_),
    .C1(_02825_),
    .X(_00741_));
 sky130_fd_sc_hd__or2_1 _18834_ (.A(\rbzero.spi_registers.buf_texadd2[10] ),
    .B(_02832_),
    .X(_02836_));
 sky130_fd_sc_hd__o211a_1 _18835_ (.A1(\rbzero.spi_registers.texadd2[10] ),
    .A2(_02831_),
    .B1(_02836_),
    .C1(_02825_),
    .X(_00742_));
 sky130_fd_sc_hd__or2_1 _18836_ (.A(\rbzero.spi_registers.buf_texadd2[11] ),
    .B(_02832_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_4 _18837_ (.A(_08091_),
    .X(_02838_));
 sky130_fd_sc_hd__buf_2 _18838_ (.A(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__o211a_1 _18839_ (.A1(\rbzero.spi_registers.texadd2[11] ),
    .A2(_02831_),
    .B1(_02837_),
    .C1(_02839_),
    .X(_00743_));
 sky130_fd_sc_hd__or2_1 _18840_ (.A(\rbzero.spi_registers.buf_texadd2[12] ),
    .B(_02832_),
    .X(_02840_));
 sky130_fd_sc_hd__o211a_1 _18841_ (.A1(\rbzero.spi_registers.texadd2[12] ),
    .A2(_02831_),
    .B1(_02840_),
    .C1(_02839_),
    .X(_00744_));
 sky130_fd_sc_hd__or2_1 _18842_ (.A(\rbzero.spi_registers.buf_texadd2[13] ),
    .B(_02832_),
    .X(_02841_));
 sky130_fd_sc_hd__o211a_1 _18843_ (.A1(\rbzero.spi_registers.texadd2[13] ),
    .A2(_02831_),
    .B1(_02841_),
    .C1(_02839_),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _18844_ (.A(\rbzero.spi_registers.buf_texadd2[14] ),
    .B(_02832_),
    .X(_02842_));
 sky130_fd_sc_hd__o211a_1 _18845_ (.A1(\rbzero.spi_registers.texadd2[14] ),
    .A2(_02831_),
    .B1(_02842_),
    .C1(_02839_),
    .X(_00746_));
 sky130_fd_sc_hd__or2_1 _18846_ (.A(\rbzero.spi_registers.buf_texadd2[15] ),
    .B(_02832_),
    .X(_02843_));
 sky130_fd_sc_hd__o211a_1 _18847_ (.A1(\rbzero.spi_registers.texadd2[15] ),
    .A2(_02831_),
    .B1(_02843_),
    .C1(_02839_),
    .X(_00747_));
 sky130_fd_sc_hd__or2_1 _18848_ (.A(\rbzero.spi_registers.buf_texadd2[16] ),
    .B(_02832_),
    .X(_02844_));
 sky130_fd_sc_hd__o211a_1 _18849_ (.A1(\rbzero.spi_registers.texadd2[16] ),
    .A2(_02831_),
    .B1(_02844_),
    .C1(_02839_),
    .X(_00748_));
 sky130_fd_sc_hd__buf_4 _18850_ (.A(_02682_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_4 _18851_ (.A(_02732_),
    .X(_02846_));
 sky130_fd_sc_hd__or2_1 _18852_ (.A(\rbzero.spi_registers.buf_texadd2[17] ),
    .B(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__o211a_1 _18853_ (.A1(\rbzero.spi_registers.texadd2[17] ),
    .A2(_02845_),
    .B1(_02847_),
    .C1(_02839_),
    .X(_00749_));
 sky130_fd_sc_hd__or2_1 _18854_ (.A(\rbzero.spi_registers.buf_texadd2[18] ),
    .B(_02846_),
    .X(_02848_));
 sky130_fd_sc_hd__o211a_1 _18855_ (.A1(\rbzero.spi_registers.texadd2[18] ),
    .A2(_02845_),
    .B1(_02848_),
    .C1(_02839_),
    .X(_00750_));
 sky130_fd_sc_hd__or2_1 _18856_ (.A(\rbzero.spi_registers.buf_texadd2[19] ),
    .B(_02846_),
    .X(_02849_));
 sky130_fd_sc_hd__o211a_1 _18857_ (.A1(\rbzero.spi_registers.texadd2[19] ),
    .A2(_02845_),
    .B1(_02849_),
    .C1(_02839_),
    .X(_00751_));
 sky130_fd_sc_hd__or2_1 _18858_ (.A(\rbzero.spi_registers.buf_texadd2[20] ),
    .B(_02846_),
    .X(_02850_));
 sky130_fd_sc_hd__o211a_1 _18859_ (.A1(\rbzero.spi_registers.texadd2[20] ),
    .A2(_02845_),
    .B1(_02850_),
    .C1(_02839_),
    .X(_00752_));
 sky130_fd_sc_hd__or2_1 _18860_ (.A(\rbzero.spi_registers.buf_texadd2[21] ),
    .B(_02846_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_4 _18861_ (.A(_02838_),
    .X(_02852_));
 sky130_fd_sc_hd__o211a_1 _18862_ (.A1(\rbzero.spi_registers.texadd2[21] ),
    .A2(_02845_),
    .B1(_02851_),
    .C1(_02852_),
    .X(_00753_));
 sky130_fd_sc_hd__or2_1 _18863_ (.A(\rbzero.spi_registers.buf_texadd2[22] ),
    .B(_02846_),
    .X(_02853_));
 sky130_fd_sc_hd__o211a_1 _18864_ (.A1(\rbzero.spi_registers.texadd2[22] ),
    .A2(_02845_),
    .B1(_02853_),
    .C1(_02852_),
    .X(_00754_));
 sky130_fd_sc_hd__or2_1 _18865_ (.A(\rbzero.spi_registers.buf_texadd2[23] ),
    .B(_02846_),
    .X(_02854_));
 sky130_fd_sc_hd__o211a_1 _18866_ (.A1(\rbzero.spi_registers.texadd2[23] ),
    .A2(_02845_),
    .B1(_02854_),
    .C1(_02852_),
    .X(_00755_));
 sky130_fd_sc_hd__or2_1 _18867_ (.A(\rbzero.spi_registers.buf_texadd3[0] ),
    .B(_02846_),
    .X(_02855_));
 sky130_fd_sc_hd__o211a_1 _18868_ (.A1(\rbzero.spi_registers.texadd3[0] ),
    .A2(_02845_),
    .B1(_02855_),
    .C1(_02852_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _18869_ (.A(\rbzero.spi_registers.buf_texadd3[1] ),
    .B(_02846_),
    .X(_02856_));
 sky130_fd_sc_hd__o211a_1 _18870_ (.A1(\rbzero.spi_registers.texadd3[1] ),
    .A2(_02845_),
    .B1(_02856_),
    .C1(_02852_),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _18871_ (.A(\rbzero.spi_registers.buf_texadd3[2] ),
    .B(_02846_),
    .X(_02857_));
 sky130_fd_sc_hd__o211a_1 _18872_ (.A1(\rbzero.spi_registers.texadd3[2] ),
    .A2(_02845_),
    .B1(_02857_),
    .C1(_02852_),
    .X(_00758_));
 sky130_fd_sc_hd__clkbuf_4 _18873_ (.A(_02682_),
    .X(_02858_));
 sky130_fd_sc_hd__buf_2 _18874_ (.A(_02732_),
    .X(_02859_));
 sky130_fd_sc_hd__or2_1 _18875_ (.A(\rbzero.spi_registers.buf_texadd3[3] ),
    .B(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__o211a_1 _18876_ (.A1(\rbzero.spi_registers.texadd3[3] ),
    .A2(_02858_),
    .B1(_02860_),
    .C1(_02852_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _18877_ (.A(\rbzero.spi_registers.buf_texadd3[4] ),
    .B(_02859_),
    .X(_02861_));
 sky130_fd_sc_hd__o211a_1 _18878_ (.A1(\rbzero.spi_registers.texadd3[4] ),
    .A2(_02858_),
    .B1(_02861_),
    .C1(_02852_),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _18879_ (.A(\rbzero.spi_registers.buf_texadd3[5] ),
    .B(_02859_),
    .X(_02862_));
 sky130_fd_sc_hd__o211a_1 _18880_ (.A1(\rbzero.spi_registers.texadd3[5] ),
    .A2(_02858_),
    .B1(_02862_),
    .C1(_02852_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _18881_ (.A(\rbzero.spi_registers.buf_texadd3[6] ),
    .B(_02859_),
    .X(_02863_));
 sky130_fd_sc_hd__o211a_1 _18882_ (.A1(\rbzero.spi_registers.texadd3[6] ),
    .A2(_02858_),
    .B1(_02863_),
    .C1(_02852_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _18883_ (.A(\rbzero.spi_registers.buf_texadd3[7] ),
    .B(_02859_),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_4 _18884_ (.A(_02838_),
    .X(_02865_));
 sky130_fd_sc_hd__o211a_1 _18885_ (.A1(\rbzero.spi_registers.texadd3[7] ),
    .A2(_02858_),
    .B1(_02864_),
    .C1(_02865_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _18886_ (.A(\rbzero.spi_registers.buf_texadd3[8] ),
    .B(_02859_),
    .X(_02866_));
 sky130_fd_sc_hd__o211a_1 _18887_ (.A1(\rbzero.spi_registers.texadd3[8] ),
    .A2(_02858_),
    .B1(_02866_),
    .C1(_02865_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _18888_ (.A(\rbzero.spi_registers.buf_texadd3[9] ),
    .B(_02859_),
    .X(_02867_));
 sky130_fd_sc_hd__o211a_1 _18889_ (.A1(\rbzero.spi_registers.texadd3[9] ),
    .A2(_02858_),
    .B1(_02867_),
    .C1(_02865_),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _18890_ (.A(\rbzero.spi_registers.buf_texadd3[10] ),
    .B(_02859_),
    .X(_02868_));
 sky130_fd_sc_hd__o211a_1 _18891_ (.A1(\rbzero.spi_registers.texadd3[10] ),
    .A2(_02858_),
    .B1(_02868_),
    .C1(_02865_),
    .X(_00766_));
 sky130_fd_sc_hd__or2_1 _18892_ (.A(\rbzero.spi_registers.buf_texadd3[11] ),
    .B(_02859_),
    .X(_02869_));
 sky130_fd_sc_hd__o211a_1 _18893_ (.A1(\rbzero.spi_registers.texadd3[11] ),
    .A2(_02858_),
    .B1(_02869_),
    .C1(_02865_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _18894_ (.A(\rbzero.spi_registers.buf_texadd3[12] ),
    .B(_02859_),
    .X(_02870_));
 sky130_fd_sc_hd__o211a_1 _18895_ (.A1(\rbzero.spi_registers.texadd3[12] ),
    .A2(_02858_),
    .B1(_02870_),
    .C1(_02865_),
    .X(_00768_));
 sky130_fd_sc_hd__buf_2 _18896_ (.A(_02682_),
    .X(_02871_));
 sky130_fd_sc_hd__clkbuf_2 _18897_ (.A(_02732_),
    .X(_02872_));
 sky130_fd_sc_hd__or2_1 _18898_ (.A(\rbzero.spi_registers.buf_texadd3[13] ),
    .B(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__o211a_1 _18899_ (.A1(\rbzero.spi_registers.texadd3[13] ),
    .A2(_02871_),
    .B1(_02873_),
    .C1(_02865_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _18900_ (.A(\rbzero.spi_registers.buf_texadd3[14] ),
    .B(_02872_),
    .X(_02874_));
 sky130_fd_sc_hd__o211a_1 _18901_ (.A1(\rbzero.spi_registers.texadd3[14] ),
    .A2(_02871_),
    .B1(_02874_),
    .C1(_02865_),
    .X(_00770_));
 sky130_fd_sc_hd__or2_1 _18902_ (.A(\rbzero.spi_registers.buf_texadd3[15] ),
    .B(_02872_),
    .X(_02875_));
 sky130_fd_sc_hd__o211a_1 _18903_ (.A1(\rbzero.spi_registers.texadd3[15] ),
    .A2(_02871_),
    .B1(_02875_),
    .C1(_02865_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _18904_ (.A(\rbzero.spi_registers.buf_texadd3[16] ),
    .B(_02872_),
    .X(_02876_));
 sky130_fd_sc_hd__o211a_1 _18905_ (.A1(\rbzero.spi_registers.texadd3[16] ),
    .A2(_02871_),
    .B1(_02876_),
    .C1(_02865_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _18906_ (.A(\rbzero.spi_registers.buf_texadd3[17] ),
    .B(_02872_),
    .X(_02877_));
 sky130_fd_sc_hd__clkbuf_4 _18907_ (.A(_02838_),
    .X(_02878_));
 sky130_fd_sc_hd__o211a_1 _18908_ (.A1(\rbzero.spi_registers.texadd3[17] ),
    .A2(_02871_),
    .B1(_02877_),
    .C1(_02878_),
    .X(_00773_));
 sky130_fd_sc_hd__or2_1 _18909_ (.A(\rbzero.spi_registers.buf_texadd3[18] ),
    .B(_02872_),
    .X(_02879_));
 sky130_fd_sc_hd__o211a_1 _18910_ (.A1(\rbzero.spi_registers.texadd3[18] ),
    .A2(_02871_),
    .B1(_02879_),
    .C1(_02878_),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _18911_ (.A(\rbzero.spi_registers.buf_texadd3[19] ),
    .B(_02872_),
    .X(_02880_));
 sky130_fd_sc_hd__o211a_1 _18912_ (.A1(\rbzero.spi_registers.texadd3[19] ),
    .A2(_02871_),
    .B1(_02880_),
    .C1(_02878_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _18913_ (.A(\rbzero.spi_registers.buf_texadd3[20] ),
    .B(_02872_),
    .X(_02881_));
 sky130_fd_sc_hd__o211a_1 _18914_ (.A1(\rbzero.spi_registers.texadd3[20] ),
    .A2(_02871_),
    .B1(_02881_),
    .C1(_02878_),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _18915_ (.A(\rbzero.spi_registers.buf_texadd3[21] ),
    .B(_02872_),
    .X(_02882_));
 sky130_fd_sc_hd__o211a_1 _18916_ (.A1(\rbzero.spi_registers.texadd3[21] ),
    .A2(_02871_),
    .B1(_02882_),
    .C1(_02878_),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _18917_ (.A(\rbzero.spi_registers.buf_texadd3[22] ),
    .B(_02872_),
    .X(_02883_));
 sky130_fd_sc_hd__o211a_1 _18918_ (.A1(\rbzero.spi_registers.texadd3[22] ),
    .A2(_02871_),
    .B1(_02883_),
    .C1(_02878_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _18919_ (.A(\rbzero.spi_registers.buf_texadd3[23] ),
    .B(_02686_),
    .X(_02884_));
 sky130_fd_sc_hd__o211a_1 _18920_ (.A1(\rbzero.spi_registers.texadd3[23] ),
    .A2(_02683_),
    .B1(_02884_),
    .C1(_02878_),
    .X(_00779_));
 sky130_fd_sc_hd__nand2_1 _18921_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02386_),
    .Y(_02885_));
 sky130_fd_sc_hd__or3_1 _18922_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .C(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__clkbuf_2 _18923_ (.A(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__mux2_1 _18924_ (.A0(\rbzero.spi_registers.spi_buffer[0] ),
    .A1(\rbzero.spi_registers.buf_sky[0] ),
    .S(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__or2_1 _18925_ (.A(_02731_),
    .B(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__clkbuf_1 _18926_ (.A(_02889_),
    .X(_00780_));
 sky130_fd_sc_hd__a31o_1 _18927_ (.A1(_02374_),
    .A2(_02384_),
    .A3(_02386_),
    .B1(\rbzero.spi_registers.buf_sky[1] ),
    .X(_02890_));
 sky130_fd_sc_hd__o211a_1 _18928_ (.A1(_02640_),
    .A2(_02887_),
    .B1(_02890_),
    .C1(_02878_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _18929_ (.A0(\rbzero.spi_registers.spi_buffer[2] ),
    .A1(\rbzero.spi_registers.buf_sky[2] ),
    .S(_02887_),
    .X(_02891_));
 sky130_fd_sc_hd__or2_1 _18930_ (.A(_04450_),
    .B(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__clkbuf_1 _18931_ (.A(_02892_),
    .X(_00782_));
 sky130_fd_sc_hd__a31o_1 _18932_ (.A1(_02374_),
    .A2(_02384_),
    .A3(_02386_),
    .B1(\rbzero.spi_registers.buf_sky[3] ),
    .X(_02893_));
 sky130_fd_sc_hd__o211a_1 _18933_ (.A1(_02644_),
    .A2(_02887_),
    .B1(_02893_),
    .C1(_02878_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _18934_ (.A0(\rbzero.spi_registers.spi_buffer[4] ),
    .A1(\rbzero.spi_registers.buf_sky[4] ),
    .S(_02887_),
    .X(_02894_));
 sky130_fd_sc_hd__or2_1 _18935_ (.A(_04450_),
    .B(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _18936_ (.A(_02895_),
    .X(_00784_));
 sky130_fd_sc_hd__a31o_1 _18937_ (.A1(_02374_),
    .A2(_02384_),
    .A3(_02386_),
    .B1(\rbzero.spi_registers.buf_sky[5] ),
    .X(_02896_));
 sky130_fd_sc_hd__o211a_1 _18938_ (.A1(_02648_),
    .A2(_02887_),
    .B1(_02896_),
    .C1(_02878_),
    .X(_00785_));
 sky130_fd_sc_hd__and2b_1 _18939_ (.A_N(\rbzero.spi_registers.spi_cmd[1] ),
    .B(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_02897_));
 sky130_fd_sc_hd__nand2_2 _18940_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__nor2_2 _18941_ (.A(_02395_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__or2_1 _18942_ (.A(\rbzero.spi_registers.buf_floor[0] ),
    .B(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__buf_4 _18943_ (.A(_08092_),
    .X(_02901_));
 sky130_fd_sc_hd__o311a_1 _18944_ (.A1(_02632_),
    .A2(_02395_),
    .A3(_02898_),
    .B1(_02900_),
    .C1(_02901_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _18945_ (.A0(\rbzero.spi_registers.buf_floor[1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_02899_),
    .X(_02902_));
 sky130_fd_sc_hd__or2_1 _18946_ (.A(_04450_),
    .B(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__clkbuf_1 _18947_ (.A(_02903_),
    .X(_00787_));
 sky130_fd_sc_hd__or2_1 _18948_ (.A(\rbzero.spi_registers.buf_floor[2] ),
    .B(_02899_),
    .X(_02904_));
 sky130_fd_sc_hd__o311a_1 _18949_ (.A1(_02642_),
    .A2(_02395_),
    .A3(_02898_),
    .B1(_02904_),
    .C1(_02901_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _18950_ (.A0(\rbzero.spi_registers.buf_floor[3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_02899_),
    .X(_02905_));
 sky130_fd_sc_hd__or2_1 _18951_ (.A(_04450_),
    .B(_02905_),
    .X(_02906_));
 sky130_fd_sc_hd__clkbuf_1 _18952_ (.A(_02906_),
    .X(_00789_));
 sky130_fd_sc_hd__or2_1 _18953_ (.A(\rbzero.spi_registers.buf_floor[4] ),
    .B(_02899_),
    .X(_02907_));
 sky130_fd_sc_hd__o311a_1 _18954_ (.A1(_02646_),
    .A2(_02395_),
    .A3(_02898_),
    .B1(_02907_),
    .C1(_02901_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _18955_ (.A0(\rbzero.spi_registers.buf_floor[5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_02899_),
    .X(_02908_));
 sky130_fd_sc_hd__or2_1 _18956_ (.A(_04450_),
    .B(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__clkbuf_1 _18957_ (.A(_02909_),
    .X(_00791_));
 sky130_fd_sc_hd__or3b_2 _18958_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02885_),
    .C_N(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02910_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18959_ (.A(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__and3_1 _18960_ (.A(_02374_),
    .B(_02386_),
    .C(_02376_),
    .X(_02912_));
 sky130_fd_sc_hd__or2_1 _18961_ (.A(\rbzero.spi_registers.buf_leak[0] ),
    .B(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_4 _18962_ (.A(_02838_),
    .X(_02914_));
 sky130_fd_sc_hd__o211a_1 _18963_ (.A1(_02632_),
    .A2(_02911_),
    .B1(_02913_),
    .C1(_02914_),
    .X(_00792_));
 sky130_fd_sc_hd__or2_1 _18964_ (.A(\rbzero.spi_registers.buf_leak[1] ),
    .B(_02912_),
    .X(_02915_));
 sky130_fd_sc_hd__o211a_1 _18965_ (.A1(_02640_),
    .A2(_02911_),
    .B1(_02915_),
    .C1(_02914_),
    .X(_00793_));
 sky130_fd_sc_hd__or2_1 _18966_ (.A(\rbzero.spi_registers.buf_leak[2] ),
    .B(_02912_),
    .X(_02916_));
 sky130_fd_sc_hd__o211a_1 _18967_ (.A1(_02642_),
    .A2(_02911_),
    .B1(_02916_),
    .C1(_02914_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _18968_ (.A(\rbzero.spi_registers.buf_leak[3] ),
    .B(_02912_),
    .X(_02917_));
 sky130_fd_sc_hd__o211a_1 _18969_ (.A1(_02644_),
    .A2(_02911_),
    .B1(_02917_),
    .C1(_02914_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _18970_ (.A(\rbzero.spi_registers.buf_leak[4] ),
    .B(_02912_),
    .X(_02918_));
 sky130_fd_sc_hd__o211a_1 _18971_ (.A1(_02646_),
    .A2(_02911_),
    .B1(_02918_),
    .C1(_02914_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _18972_ (.A(\rbzero.spi_registers.buf_leak[5] ),
    .B(_02912_),
    .X(_02919_));
 sky130_fd_sc_hd__o211a_1 _18973_ (.A1(_02648_),
    .A2(_02911_),
    .B1(_02919_),
    .C1(_02914_),
    .X(_00797_));
 sky130_fd_sc_hd__nor2_4 _18974_ (.A(_02380_),
    .B(_02885_),
    .Y(_02920_));
 sky130_fd_sc_hd__or2_2 _18975_ (.A(_02380_),
    .B(_02885_),
    .X(_02921_));
 sky130_fd_sc_hd__or2_1 _18976_ (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .B(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__o211a_1 _18977_ (.A1(\rbzero.spi_registers.buf_otherx[0] ),
    .A2(_02920_),
    .B1(_02922_),
    .C1(_02914_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _18978_ (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .B(_02921_),
    .X(_02923_));
 sky130_fd_sc_hd__o211a_1 _18979_ (.A1(\rbzero.spi_registers.buf_otherx[1] ),
    .A2(_02920_),
    .B1(_02923_),
    .C1(_02914_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _18980_ (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .B(_02921_),
    .X(_02924_));
 sky130_fd_sc_hd__o211a_1 _18981_ (.A1(\rbzero.spi_registers.buf_otherx[2] ),
    .A2(_02920_),
    .B1(_02924_),
    .C1(_02914_),
    .X(_00800_));
 sky130_fd_sc_hd__or2_1 _18982_ (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .B(_02921_),
    .X(_02925_));
 sky130_fd_sc_hd__o211a_1 _18983_ (.A1(\rbzero.spi_registers.buf_otherx[3] ),
    .A2(_02920_),
    .B1(_02925_),
    .C1(_02914_),
    .X(_00801_));
 sky130_fd_sc_hd__or2_1 _18984_ (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .B(_02921_),
    .X(_02926_));
 sky130_fd_sc_hd__buf_4 _18985_ (.A(_02838_),
    .X(_02927_));
 sky130_fd_sc_hd__o211a_1 _18986_ (.A1(\rbzero.spi_registers.buf_otherx[4] ),
    .A2(_02920_),
    .B1(_02926_),
    .C1(_02927_),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _18987_ (.A(_02632_),
    .B(_02921_),
    .X(_02928_));
 sky130_fd_sc_hd__o211a_1 _18988_ (.A1(\rbzero.spi_registers.buf_othery[0] ),
    .A2(_02920_),
    .B1(_02928_),
    .C1(_02927_),
    .X(_00803_));
 sky130_fd_sc_hd__or2_1 _18989_ (.A(_02640_),
    .B(_02921_),
    .X(_02929_));
 sky130_fd_sc_hd__o211a_1 _18990_ (.A1(\rbzero.spi_registers.buf_othery[1] ),
    .A2(_02920_),
    .B1(_02929_),
    .C1(_02927_),
    .X(_00804_));
 sky130_fd_sc_hd__or2_1 _18991_ (.A(_02642_),
    .B(_02921_),
    .X(_02930_));
 sky130_fd_sc_hd__o211a_1 _18992_ (.A1(\rbzero.spi_registers.buf_othery[2] ),
    .A2(_02920_),
    .B1(_02930_),
    .C1(_02927_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _18993_ (.A(_02644_),
    .B(_02921_),
    .X(_02931_));
 sky130_fd_sc_hd__o211a_1 _18994_ (.A1(\rbzero.spi_registers.buf_othery[3] ),
    .A2(_02920_),
    .B1(_02931_),
    .C1(_02927_),
    .X(_00806_));
 sky130_fd_sc_hd__or2_1 _18995_ (.A(_02646_),
    .B(_02921_),
    .X(_02932_));
 sky130_fd_sc_hd__o211a_1 _18996_ (.A1(\rbzero.spi_registers.buf_othery[4] ),
    .A2(_02920_),
    .B1(_02932_),
    .C1(_02927_),
    .X(_00807_));
 sky130_fd_sc_hd__nand2_2 _18997_ (.A(_02374_),
    .B(_02385_),
    .Y(_02933_));
 sky130_fd_sc_hd__and3_2 _18998_ (.A(_02374_),
    .B(_02375_),
    .C(_02384_),
    .X(_02934_));
 sky130_fd_sc_hd__or2_1 _18999_ (.A(\rbzero.spi_registers.buf_vshift[0] ),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__o211a_1 _19000_ (.A1(_02632_),
    .A2(_02933_),
    .B1(_02935_),
    .C1(_02927_),
    .X(_00808_));
 sky130_fd_sc_hd__or2_1 _19001_ (.A(\rbzero.spi_registers.buf_vshift[1] ),
    .B(_02934_),
    .X(_02936_));
 sky130_fd_sc_hd__o211a_1 _19002_ (.A1(_02640_),
    .A2(_02933_),
    .B1(_02936_),
    .C1(_02927_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _19003_ (.A(\rbzero.spi_registers.buf_vshift[2] ),
    .B(_02934_),
    .X(_02937_));
 sky130_fd_sc_hd__o211a_1 _19004_ (.A1(_02642_),
    .A2(_02933_),
    .B1(_02937_),
    .C1(_02927_),
    .X(_00810_));
 sky130_fd_sc_hd__or2_1 _19005_ (.A(\rbzero.spi_registers.buf_vshift[3] ),
    .B(_02934_),
    .X(_02938_));
 sky130_fd_sc_hd__o211a_1 _19006_ (.A1(_02644_),
    .A2(_02933_),
    .B1(_02938_),
    .C1(_02927_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _19007_ (.A(\rbzero.spi_registers.buf_vshift[4] ),
    .B(_02934_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_4 _19008_ (.A(_02838_),
    .X(_02940_));
 sky130_fd_sc_hd__o211a_1 _19009_ (.A1(_02646_),
    .A2(_02933_),
    .B1(_02939_),
    .C1(_02940_),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _19010_ (.A(\rbzero.spi_registers.buf_vshift[5] ),
    .B(_02934_),
    .X(_02941_));
 sky130_fd_sc_hd__o211a_1 _19011_ (.A1(_02648_),
    .A2(_02933_),
    .B1(_02941_),
    .C1(_02940_),
    .X(_00813_));
 sky130_fd_sc_hd__a31o_1 _19012_ (.A1(_02374_),
    .A2(_02375_),
    .A3(_02897_),
    .B1(\rbzero.spi_registers.buf_vinf ),
    .X(_02942_));
 sky130_fd_sc_hd__o311a_1 _19013_ (.A1(_02632_),
    .A2(_02377_),
    .A3(_02898_),
    .B1(_02942_),
    .C1(_02901_),
    .X(_00814_));
 sky130_fd_sc_hd__nand2_1 _19014_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02375_),
    .Y(_02943_));
 sky130_fd_sc_hd__or3b_1 _19015_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02943_),
    .C_N(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_2 _19016_ (.A(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__buf_2 _19017_ (.A(_02945_),
    .X(_02946_));
 sky130_fd_sc_hd__and3_1 _19018_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02375_),
    .C(_02376_),
    .X(_02947_));
 sky130_fd_sc_hd__clkbuf_2 _19019_ (.A(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__or2_1 _19020_ (.A(\rbzero.spi_registers.buf_mapdx[0] ),
    .B(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__o211a_1 _19021_ (.A1(\rbzero.spi_registers.spi_buffer[10] ),
    .A2(_02946_),
    .B1(_02949_),
    .C1(_02940_),
    .X(_00815_));
 sky130_fd_sc_hd__or2_1 _19022_ (.A(\rbzero.spi_registers.buf_mapdx[1] ),
    .B(_02948_),
    .X(_02950_));
 sky130_fd_sc_hd__o211a_1 _19023_ (.A1(\rbzero.spi_registers.spi_buffer[11] ),
    .A2(_02946_),
    .B1(_02950_),
    .C1(_02940_),
    .X(_00816_));
 sky130_fd_sc_hd__or2_1 _19024_ (.A(\rbzero.spi_registers.buf_mapdx[2] ),
    .B(_02948_),
    .X(_02951_));
 sky130_fd_sc_hd__o211a_1 _19025_ (.A1(\rbzero.spi_registers.spi_buffer[12] ),
    .A2(_02946_),
    .B1(_02951_),
    .C1(_02940_),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _19026_ (.A(\rbzero.spi_registers.buf_mapdx[3] ),
    .B(_02948_),
    .X(_02952_));
 sky130_fd_sc_hd__o211a_1 _19027_ (.A1(\rbzero.spi_registers.spi_buffer[13] ),
    .A2(_02946_),
    .B1(_02952_),
    .C1(_02940_),
    .X(_00818_));
 sky130_fd_sc_hd__or2_1 _19028_ (.A(\rbzero.spi_registers.buf_mapdx[4] ),
    .B(_02948_),
    .X(_02953_));
 sky130_fd_sc_hd__o211a_1 _19029_ (.A1(\rbzero.spi_registers.spi_buffer[14] ),
    .A2(_02946_),
    .B1(_02953_),
    .C1(_02940_),
    .X(_00819_));
 sky130_fd_sc_hd__or2_1 _19030_ (.A(\rbzero.spi_registers.buf_mapdx[5] ),
    .B(_02948_),
    .X(_02954_));
 sky130_fd_sc_hd__o211a_1 _19031_ (.A1(\rbzero.spi_registers.spi_buffer[15] ),
    .A2(_02946_),
    .B1(_02954_),
    .C1(_02940_),
    .X(_00820_));
 sky130_fd_sc_hd__or2_1 _19032_ (.A(\rbzero.spi_registers.buf_mapdy[0] ),
    .B(_02948_),
    .X(_02955_));
 sky130_fd_sc_hd__o211a_1 _19033_ (.A1(_02646_),
    .A2(_02946_),
    .B1(_02955_),
    .C1(_02940_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _19034_ (.A(\rbzero.spi_registers.buf_mapdy[1] ),
    .B(_02948_),
    .X(_02956_));
 sky130_fd_sc_hd__o211a_1 _19035_ (.A1(_02648_),
    .A2(_02946_),
    .B1(_02956_),
    .C1(_02940_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _19036_ (.A(\rbzero.spi_registers.buf_mapdy[2] ),
    .B(_02948_),
    .X(_02957_));
 sky130_fd_sc_hd__clkbuf_4 _19037_ (.A(_02838_),
    .X(_02958_));
 sky130_fd_sc_hd__o211a_1 _19038_ (.A1(\rbzero.spi_registers.spi_buffer[6] ),
    .A2(_02946_),
    .B1(_02957_),
    .C1(_02958_),
    .X(_00823_));
 sky130_fd_sc_hd__or2_1 _19039_ (.A(\rbzero.spi_registers.buf_mapdy[3] ),
    .B(_02948_),
    .X(_02959_));
 sky130_fd_sc_hd__o211a_1 _19040_ (.A1(\rbzero.spi_registers.spi_buffer[7] ),
    .A2(_02946_),
    .B1(_02959_),
    .C1(_02958_),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _19041_ (.A(\rbzero.spi_registers.buf_mapdy[4] ),
    .B(_02947_),
    .X(_02960_));
 sky130_fd_sc_hd__o211a_1 _19042_ (.A1(\rbzero.spi_registers.spi_buffer[8] ),
    .A2(_02945_),
    .B1(_02960_),
    .C1(_02958_),
    .X(_00825_));
 sky130_fd_sc_hd__or2_1 _19043_ (.A(\rbzero.spi_registers.buf_mapdy[5] ),
    .B(_02947_),
    .X(_02961_));
 sky130_fd_sc_hd__o211a_1 _19044_ (.A1(\rbzero.spi_registers.spi_buffer[9] ),
    .A2(_02945_),
    .B1(_02961_),
    .C1(_02958_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _19045_ (.A(\rbzero.spi_registers.buf_mapdxw[0] ),
    .B(_02947_),
    .X(_02962_));
 sky130_fd_sc_hd__o211a_1 _19046_ (.A1(_02642_),
    .A2(_02945_),
    .B1(_02962_),
    .C1(_02958_),
    .X(_00827_));
 sky130_fd_sc_hd__or2_1 _19047_ (.A(\rbzero.spi_registers.buf_mapdxw[1] ),
    .B(_02947_),
    .X(_02963_));
 sky130_fd_sc_hd__o211a_1 _19048_ (.A1(_02644_),
    .A2(_02945_),
    .B1(_02963_),
    .C1(_02958_),
    .X(_00828_));
 sky130_fd_sc_hd__or2_1 _19049_ (.A(\rbzero.spi_registers.buf_mapdyw[0] ),
    .B(_02947_),
    .X(_02964_));
 sky130_fd_sc_hd__o211a_1 _19050_ (.A1(_02632_),
    .A2(_02945_),
    .B1(_02964_),
    .C1(_02958_),
    .X(_00829_));
 sky130_fd_sc_hd__or2_1 _19051_ (.A(\rbzero.spi_registers.buf_mapdyw[1] ),
    .B(_02947_),
    .X(_02965_));
 sky130_fd_sc_hd__o211a_1 _19052_ (.A1(_02640_),
    .A2(_02945_),
    .B1(_02965_),
    .C1(_02958_),
    .X(_00830_));
 sky130_fd_sc_hd__nor2_2 _19053_ (.A(_02380_),
    .B(_02943_),
    .Y(_02966_));
 sky130_fd_sc_hd__clkbuf_4 _19054_ (.A(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__or2_2 _19055_ (.A(_02380_),
    .B(_02943_),
    .X(_02968_));
 sky130_fd_sc_hd__buf_2 _19056_ (.A(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__or2_1 _19057_ (.A(_02632_),
    .B(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__o211a_1 _19058_ (.A1(\rbzero.spi_registers.buf_texadd0[0] ),
    .A2(_02967_),
    .B1(_02970_),
    .C1(_02958_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _19059_ (.A(_02640_),
    .B(_02969_),
    .X(_02971_));
 sky130_fd_sc_hd__o211a_1 _19060_ (.A1(\rbzero.spi_registers.buf_texadd0[1] ),
    .A2(_02967_),
    .B1(_02971_),
    .C1(_02958_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _19061_ (.A(_02642_),
    .B(_02969_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_4 _19062_ (.A(_02838_),
    .X(_02973_));
 sky130_fd_sc_hd__o211a_1 _19063_ (.A1(\rbzero.spi_registers.buf_texadd0[2] ),
    .A2(_02967_),
    .B1(_02972_),
    .C1(_02973_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_1 _19064_ (.A(_02644_),
    .B(_02969_),
    .X(_02974_));
 sky130_fd_sc_hd__o211a_1 _19065_ (.A1(\rbzero.spi_registers.buf_texadd0[3] ),
    .A2(_02967_),
    .B1(_02974_),
    .C1(_02973_),
    .X(_00834_));
 sky130_fd_sc_hd__or2_1 _19066_ (.A(_02646_),
    .B(_02969_),
    .X(_02975_));
 sky130_fd_sc_hd__o211a_1 _19067_ (.A1(\rbzero.spi_registers.buf_texadd0[4] ),
    .A2(_02967_),
    .B1(_02975_),
    .C1(_02973_),
    .X(_00835_));
 sky130_fd_sc_hd__or2_1 _19068_ (.A(_02648_),
    .B(_02969_),
    .X(_02976_));
 sky130_fd_sc_hd__o211a_1 _19069_ (.A1(\rbzero.spi_registers.buf_texadd0[5] ),
    .A2(_02967_),
    .B1(_02976_),
    .C1(_02973_),
    .X(_00836_));
 sky130_fd_sc_hd__or2_1 _19070_ (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .B(_02969_),
    .X(_02977_));
 sky130_fd_sc_hd__o211a_1 _19071_ (.A1(\rbzero.spi_registers.buf_texadd0[6] ),
    .A2(_02967_),
    .B1(_02977_),
    .C1(_02973_),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _19072_ (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .B(_02969_),
    .X(_02978_));
 sky130_fd_sc_hd__o211a_1 _19073_ (.A1(\rbzero.spi_registers.buf_texadd0[7] ),
    .A2(_02967_),
    .B1(_02978_),
    .C1(_02973_),
    .X(_00838_));
 sky130_fd_sc_hd__or2_1 _19074_ (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .B(_02969_),
    .X(_02979_));
 sky130_fd_sc_hd__o211a_1 _19075_ (.A1(\rbzero.spi_registers.buf_texadd0[8] ),
    .A2(_02967_),
    .B1(_02979_),
    .C1(_02973_),
    .X(_00839_));
 sky130_fd_sc_hd__or2_1 _19076_ (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .B(_02969_),
    .X(_02980_));
 sky130_fd_sc_hd__o211a_1 _19077_ (.A1(\rbzero.spi_registers.buf_texadd0[9] ),
    .A2(_02967_),
    .B1(_02980_),
    .C1(_02973_),
    .X(_00840_));
 sky130_fd_sc_hd__buf_2 _19078_ (.A(_02966_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_2 _19079_ (.A(_02968_),
    .X(_02982_));
 sky130_fd_sc_hd__or2_1 _19080_ (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .B(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__o211a_1 _19081_ (.A1(\rbzero.spi_registers.buf_texadd0[10] ),
    .A2(_02981_),
    .B1(_02983_),
    .C1(_02973_),
    .X(_00841_));
 sky130_fd_sc_hd__or2_1 _19082_ (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .B(_02982_),
    .X(_02984_));
 sky130_fd_sc_hd__o211a_1 _19083_ (.A1(\rbzero.spi_registers.buf_texadd0[11] ),
    .A2(_02981_),
    .B1(_02984_),
    .C1(_02973_),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _19084_ (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .B(_02982_),
    .X(_02985_));
 sky130_fd_sc_hd__buf_2 _19085_ (.A(_02838_),
    .X(_02986_));
 sky130_fd_sc_hd__o211a_1 _19086_ (.A1(\rbzero.spi_registers.buf_texadd0[12] ),
    .A2(_02981_),
    .B1(_02985_),
    .C1(_02986_),
    .X(_00843_));
 sky130_fd_sc_hd__or2_1 _19087_ (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .B(_02982_),
    .X(_02987_));
 sky130_fd_sc_hd__o211a_1 _19088_ (.A1(\rbzero.spi_registers.buf_texadd0[13] ),
    .A2(_02981_),
    .B1(_02987_),
    .C1(_02986_),
    .X(_00844_));
 sky130_fd_sc_hd__or2_1 _19089_ (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .B(_02982_),
    .X(_02988_));
 sky130_fd_sc_hd__o211a_1 _19090_ (.A1(\rbzero.spi_registers.buf_texadd0[14] ),
    .A2(_02981_),
    .B1(_02988_),
    .C1(_02986_),
    .X(_00845_));
 sky130_fd_sc_hd__or2_1 _19091_ (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .B(_02982_),
    .X(_02989_));
 sky130_fd_sc_hd__o211a_1 _19092_ (.A1(\rbzero.spi_registers.buf_texadd0[15] ),
    .A2(_02981_),
    .B1(_02989_),
    .C1(_02986_),
    .X(_00846_));
 sky130_fd_sc_hd__or2_1 _19093_ (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .B(_02982_),
    .X(_02990_));
 sky130_fd_sc_hd__o211a_1 _19094_ (.A1(\rbzero.spi_registers.buf_texadd0[16] ),
    .A2(_02981_),
    .B1(_02990_),
    .C1(_02986_),
    .X(_00847_));
 sky130_fd_sc_hd__or2_1 _19095_ (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .B(_02982_),
    .X(_02991_));
 sky130_fd_sc_hd__o211a_1 _19096_ (.A1(\rbzero.spi_registers.buf_texadd0[17] ),
    .A2(_02981_),
    .B1(_02991_),
    .C1(_02986_),
    .X(_00848_));
 sky130_fd_sc_hd__or2_1 _19097_ (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .B(_02982_),
    .X(_02992_));
 sky130_fd_sc_hd__o211a_1 _19098_ (.A1(\rbzero.spi_registers.buf_texadd0[18] ),
    .A2(_02981_),
    .B1(_02992_),
    .C1(_02986_),
    .X(_00849_));
 sky130_fd_sc_hd__or2_1 _19099_ (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .B(_02982_),
    .X(_02993_));
 sky130_fd_sc_hd__o211a_1 _19100_ (.A1(\rbzero.spi_registers.buf_texadd0[19] ),
    .A2(_02981_),
    .B1(_02993_),
    .C1(_02986_),
    .X(_00850_));
 sky130_fd_sc_hd__or2_1 _19101_ (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .B(_02968_),
    .X(_02994_));
 sky130_fd_sc_hd__o211a_1 _19102_ (.A1(\rbzero.spi_registers.buf_texadd0[20] ),
    .A2(_02966_),
    .B1(_02994_),
    .C1(_02986_),
    .X(_00851_));
 sky130_fd_sc_hd__or2_1 _19103_ (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .B(_02968_),
    .X(_02995_));
 sky130_fd_sc_hd__o211a_1 _19104_ (.A1(\rbzero.spi_registers.buf_texadd0[21] ),
    .A2(_02966_),
    .B1(_02995_),
    .C1(_02986_),
    .X(_00852_));
 sky130_fd_sc_hd__or2_1 _19105_ (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .B(_02968_),
    .X(_02996_));
 sky130_fd_sc_hd__buf_4 _19106_ (.A(_08091_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_4 _19107_ (.A(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__o211a_1 _19108_ (.A1(\rbzero.spi_registers.buf_texadd0[22] ),
    .A2(_02966_),
    .B1(_02996_),
    .C1(_02998_),
    .X(_00853_));
 sky130_fd_sc_hd__or2_1 _19109_ (.A(\rbzero.spi_registers.spi_buffer[23] ),
    .B(_02968_),
    .X(_02999_));
 sky130_fd_sc_hd__o211a_1 _19110_ (.A1(\rbzero.spi_registers.buf_texadd0[23] ),
    .A2(_02966_),
    .B1(_02999_),
    .C1(_02998_),
    .X(_00854_));
 sky130_fd_sc_hd__and3_1 _19111_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02384_),
    .C(_02378_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_2 _19112_ (.A(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_4 _19113_ (.A(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__nand3_2 _19114_ (.A(_02374_),
    .B(_02384_),
    .C(_02378_),
    .Y(_03003_));
 sky130_fd_sc_hd__buf_2 _19115_ (.A(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__or2_1 _19116_ (.A(_02632_),
    .B(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__o211a_1 _19117_ (.A1(\rbzero.spi_registers.buf_texadd1[0] ),
    .A2(_03002_),
    .B1(_03005_),
    .C1(_02998_),
    .X(_00855_));
 sky130_fd_sc_hd__or2_1 _19118_ (.A(_02640_),
    .B(_03004_),
    .X(_03006_));
 sky130_fd_sc_hd__o211a_1 _19119_ (.A1(\rbzero.spi_registers.buf_texadd1[1] ),
    .A2(_03002_),
    .B1(_03006_),
    .C1(_02998_),
    .X(_00856_));
 sky130_fd_sc_hd__or2_1 _19120_ (.A(_02642_),
    .B(_03004_),
    .X(_03007_));
 sky130_fd_sc_hd__o211a_1 _19121_ (.A1(\rbzero.spi_registers.buf_texadd1[2] ),
    .A2(_03002_),
    .B1(_03007_),
    .C1(_02998_),
    .X(_00857_));
 sky130_fd_sc_hd__or2_1 _19122_ (.A(_02644_),
    .B(_03004_),
    .X(_03008_));
 sky130_fd_sc_hd__o211a_1 _19123_ (.A1(\rbzero.spi_registers.buf_texadd1[3] ),
    .A2(_03002_),
    .B1(_03008_),
    .C1(_02998_),
    .X(_00858_));
 sky130_fd_sc_hd__or2_1 _19124_ (.A(_02646_),
    .B(_03004_),
    .X(_03009_));
 sky130_fd_sc_hd__o211a_1 _19125_ (.A1(\rbzero.spi_registers.buf_texadd1[4] ),
    .A2(_03002_),
    .B1(_03009_),
    .C1(_02998_),
    .X(_00859_));
 sky130_fd_sc_hd__or2_1 _19126_ (.A(_02648_),
    .B(_03004_),
    .X(_03010_));
 sky130_fd_sc_hd__o211a_1 _19127_ (.A1(\rbzero.spi_registers.buf_texadd1[5] ),
    .A2(_03002_),
    .B1(_03010_),
    .C1(_02998_),
    .X(_00860_));
 sky130_fd_sc_hd__or2_1 _19128_ (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .B(_03004_),
    .X(_03011_));
 sky130_fd_sc_hd__o211a_1 _19129_ (.A1(\rbzero.spi_registers.buf_texadd1[6] ),
    .A2(_03002_),
    .B1(_03011_),
    .C1(_02998_),
    .X(_00861_));
 sky130_fd_sc_hd__or2_1 _19130_ (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .B(_03004_),
    .X(_03012_));
 sky130_fd_sc_hd__o211a_1 _19131_ (.A1(\rbzero.spi_registers.buf_texadd1[7] ),
    .A2(_03002_),
    .B1(_03012_),
    .C1(_02998_),
    .X(_00862_));
 sky130_fd_sc_hd__or2_1 _19132_ (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .B(_03004_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_4 _19133_ (.A(_02997_),
    .X(_03014_));
 sky130_fd_sc_hd__o211a_1 _19134_ (.A1(\rbzero.spi_registers.buf_texadd1[8] ),
    .A2(_03002_),
    .B1(_03013_),
    .C1(_03014_),
    .X(_00863_));
 sky130_fd_sc_hd__or2_1 _19135_ (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .B(_03004_),
    .X(_03015_));
 sky130_fd_sc_hd__o211a_1 _19136_ (.A1(\rbzero.spi_registers.buf_texadd1[9] ),
    .A2(_03002_),
    .B1(_03015_),
    .C1(_03014_),
    .X(_00864_));
 sky130_fd_sc_hd__buf_2 _19137_ (.A(_03001_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_2 _19138_ (.A(_03003_),
    .X(_03017_));
 sky130_fd_sc_hd__or2_1 _19139_ (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .B(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__o211a_1 _19140_ (.A1(\rbzero.spi_registers.buf_texadd1[10] ),
    .A2(_03016_),
    .B1(_03018_),
    .C1(_03014_),
    .X(_00865_));
 sky130_fd_sc_hd__or2_1 _19141_ (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .B(_03017_),
    .X(_03019_));
 sky130_fd_sc_hd__o211a_1 _19142_ (.A1(\rbzero.spi_registers.buf_texadd1[11] ),
    .A2(_03016_),
    .B1(_03019_),
    .C1(_03014_),
    .X(_00866_));
 sky130_fd_sc_hd__or2_1 _19143_ (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .B(_03017_),
    .X(_03020_));
 sky130_fd_sc_hd__o211a_1 _19144_ (.A1(\rbzero.spi_registers.buf_texadd1[12] ),
    .A2(_03016_),
    .B1(_03020_),
    .C1(_03014_),
    .X(_00867_));
 sky130_fd_sc_hd__or2_1 _19145_ (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .B(_03017_),
    .X(_03021_));
 sky130_fd_sc_hd__o211a_1 _19146_ (.A1(\rbzero.spi_registers.buf_texadd1[13] ),
    .A2(_03016_),
    .B1(_03021_),
    .C1(_03014_),
    .X(_00868_));
 sky130_fd_sc_hd__or2_1 _19147_ (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .B(_03017_),
    .X(_03022_));
 sky130_fd_sc_hd__o211a_1 _19148_ (.A1(\rbzero.spi_registers.buf_texadd1[14] ),
    .A2(_03016_),
    .B1(_03022_),
    .C1(_03014_),
    .X(_00869_));
 sky130_fd_sc_hd__or2_1 _19149_ (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .B(_03017_),
    .X(_03023_));
 sky130_fd_sc_hd__o211a_1 _19150_ (.A1(\rbzero.spi_registers.buf_texadd1[15] ),
    .A2(_03016_),
    .B1(_03023_),
    .C1(_03014_),
    .X(_00870_));
 sky130_fd_sc_hd__or2_1 _19151_ (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .B(_03017_),
    .X(_03024_));
 sky130_fd_sc_hd__o211a_1 _19152_ (.A1(\rbzero.spi_registers.buf_texadd1[16] ),
    .A2(_03016_),
    .B1(_03024_),
    .C1(_03014_),
    .X(_00871_));
 sky130_fd_sc_hd__or2_1 _19153_ (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .B(_03017_),
    .X(_03025_));
 sky130_fd_sc_hd__o211a_1 _19154_ (.A1(\rbzero.spi_registers.buf_texadd1[17] ),
    .A2(_03016_),
    .B1(_03025_),
    .C1(_03014_),
    .X(_00872_));
 sky130_fd_sc_hd__or2_1 _19155_ (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .B(_03017_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_4 _19156_ (.A(_02997_),
    .X(_03027_));
 sky130_fd_sc_hd__o211a_1 _19157_ (.A1(\rbzero.spi_registers.buf_texadd1[18] ),
    .A2(_03016_),
    .B1(_03026_),
    .C1(_03027_),
    .X(_00873_));
 sky130_fd_sc_hd__or2_1 _19158_ (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .B(_03017_),
    .X(_03028_));
 sky130_fd_sc_hd__o211a_1 _19159_ (.A1(\rbzero.spi_registers.buf_texadd1[19] ),
    .A2(_03016_),
    .B1(_03028_),
    .C1(_03027_),
    .X(_00874_));
 sky130_fd_sc_hd__or2_1 _19160_ (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .B(_03003_),
    .X(_03029_));
 sky130_fd_sc_hd__o211a_1 _19161_ (.A1(\rbzero.spi_registers.buf_texadd1[20] ),
    .A2(_03001_),
    .B1(_03029_),
    .C1(_03027_),
    .X(_00875_));
 sky130_fd_sc_hd__or2_1 _19162_ (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .B(_03003_),
    .X(_03030_));
 sky130_fd_sc_hd__o211a_1 _19163_ (.A1(\rbzero.spi_registers.buf_texadd1[21] ),
    .A2(_03001_),
    .B1(_03030_),
    .C1(_03027_),
    .X(_00876_));
 sky130_fd_sc_hd__or2_1 _19164_ (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .B(_03003_),
    .X(_03031_));
 sky130_fd_sc_hd__o211a_1 _19165_ (.A1(\rbzero.spi_registers.buf_texadd1[22] ),
    .A2(_03001_),
    .B1(_03031_),
    .C1(_03027_),
    .X(_00877_));
 sky130_fd_sc_hd__or2_1 _19166_ (.A(\rbzero.spi_registers.spi_buffer[23] ),
    .B(_03003_),
    .X(_03032_));
 sky130_fd_sc_hd__o211a_1 _19167_ (.A1(\rbzero.spi_registers.buf_texadd1[23] ),
    .A2(_03001_),
    .B1(_03032_),
    .C1(_03027_),
    .X(_00878_));
 sky130_fd_sc_hd__and3_1 _19168_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02378_),
    .C(_02897_),
    .X(_03033_));
 sky130_fd_sc_hd__buf_2 _19169_ (.A(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__buf_2 _19170_ (.A(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__nand3_4 _19171_ (.A(_02374_),
    .B(_02378_),
    .C(_02897_),
    .Y(_03036_));
 sky130_fd_sc_hd__clkbuf_2 _19172_ (.A(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__or2_1 _19173_ (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .B(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__o211a_1 _19174_ (.A1(\rbzero.spi_registers.buf_texadd2[0] ),
    .A2(_03035_),
    .B1(_03038_),
    .C1(_03027_),
    .X(_00879_));
 sky130_fd_sc_hd__or2_1 _19175_ (.A(_02640_),
    .B(_03037_),
    .X(_03039_));
 sky130_fd_sc_hd__o211a_1 _19176_ (.A1(\rbzero.spi_registers.buf_texadd2[1] ),
    .A2(_03035_),
    .B1(_03039_),
    .C1(_03027_),
    .X(_00880_));
 sky130_fd_sc_hd__or2_1 _19177_ (.A(_02642_),
    .B(_03037_),
    .X(_03040_));
 sky130_fd_sc_hd__o211a_1 _19178_ (.A1(\rbzero.spi_registers.buf_texadd2[2] ),
    .A2(_03035_),
    .B1(_03040_),
    .C1(_03027_),
    .X(_00881_));
 sky130_fd_sc_hd__or2_1 _19179_ (.A(_02644_),
    .B(_03037_),
    .X(_03041_));
 sky130_fd_sc_hd__o211a_1 _19180_ (.A1(\rbzero.spi_registers.buf_texadd2[3] ),
    .A2(_03035_),
    .B1(_03041_),
    .C1(_03027_),
    .X(_00882_));
 sky130_fd_sc_hd__or2_1 _19181_ (.A(_02646_),
    .B(_03037_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_4 _19182_ (.A(_02997_),
    .X(_03043_));
 sky130_fd_sc_hd__o211a_1 _19183_ (.A1(\rbzero.spi_registers.buf_texadd2[4] ),
    .A2(_03035_),
    .B1(_03042_),
    .C1(_03043_),
    .X(_00883_));
 sky130_fd_sc_hd__or2_1 _19184_ (.A(_02648_),
    .B(_03037_),
    .X(_03044_));
 sky130_fd_sc_hd__o211a_1 _19185_ (.A1(\rbzero.spi_registers.buf_texadd2[5] ),
    .A2(_03035_),
    .B1(_03044_),
    .C1(_03043_),
    .X(_00884_));
 sky130_fd_sc_hd__or2_1 _19186_ (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .B(_03037_),
    .X(_03045_));
 sky130_fd_sc_hd__o211a_1 _19187_ (.A1(\rbzero.spi_registers.buf_texadd2[6] ),
    .A2(_03035_),
    .B1(_03045_),
    .C1(_03043_),
    .X(_00885_));
 sky130_fd_sc_hd__or2_1 _19188_ (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .B(_03037_),
    .X(_03046_));
 sky130_fd_sc_hd__o211a_1 _19189_ (.A1(\rbzero.spi_registers.buf_texadd2[7] ),
    .A2(_03035_),
    .B1(_03046_),
    .C1(_03043_),
    .X(_00886_));
 sky130_fd_sc_hd__or2_1 _19190_ (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .B(_03037_),
    .X(_03047_));
 sky130_fd_sc_hd__o211a_1 _19191_ (.A1(\rbzero.spi_registers.buf_texadd2[8] ),
    .A2(_03035_),
    .B1(_03047_),
    .C1(_03043_),
    .X(_00887_));
 sky130_fd_sc_hd__or2_1 _19192_ (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .B(_03037_),
    .X(_03048_));
 sky130_fd_sc_hd__o211a_1 _19193_ (.A1(\rbzero.spi_registers.buf_texadd2[9] ),
    .A2(_03035_),
    .B1(_03048_),
    .C1(_03043_),
    .X(_00888_));
 sky130_fd_sc_hd__clkbuf_4 _19194_ (.A(_03034_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_2 _19195_ (.A(_03036_),
    .X(_03050_));
 sky130_fd_sc_hd__or2_1 _19196_ (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .B(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__o211a_1 _19197_ (.A1(\rbzero.spi_registers.buf_texadd2[10] ),
    .A2(_03049_),
    .B1(_03051_),
    .C1(_03043_),
    .X(_00889_));
 sky130_fd_sc_hd__or2_1 _19198_ (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .B(_03050_),
    .X(_03052_));
 sky130_fd_sc_hd__o211a_1 _19199_ (.A1(\rbzero.spi_registers.buf_texadd2[11] ),
    .A2(_03049_),
    .B1(_03052_),
    .C1(_03043_),
    .X(_00890_));
 sky130_fd_sc_hd__or2_1 _19200_ (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .B(_03050_),
    .X(_03053_));
 sky130_fd_sc_hd__o211a_1 _19201_ (.A1(\rbzero.spi_registers.buf_texadd2[12] ),
    .A2(_03049_),
    .B1(_03053_),
    .C1(_03043_),
    .X(_00891_));
 sky130_fd_sc_hd__or2_1 _19202_ (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .B(_03050_),
    .X(_03054_));
 sky130_fd_sc_hd__o211a_1 _19203_ (.A1(\rbzero.spi_registers.buf_texadd2[13] ),
    .A2(_03049_),
    .B1(_03054_),
    .C1(_03043_),
    .X(_00892_));
 sky130_fd_sc_hd__or2_1 _19204_ (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .B(_03050_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_4 _19205_ (.A(_02997_),
    .X(_03056_));
 sky130_fd_sc_hd__o211a_1 _19206_ (.A1(\rbzero.spi_registers.buf_texadd2[14] ),
    .A2(_03049_),
    .B1(_03055_),
    .C1(_03056_),
    .X(_00893_));
 sky130_fd_sc_hd__or2_1 _19207_ (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .B(_03050_),
    .X(_03057_));
 sky130_fd_sc_hd__o211a_1 _19208_ (.A1(\rbzero.spi_registers.buf_texadd2[15] ),
    .A2(_03049_),
    .B1(_03057_),
    .C1(_03056_),
    .X(_00894_));
 sky130_fd_sc_hd__or2_1 _19209_ (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .B(_03050_),
    .X(_03058_));
 sky130_fd_sc_hd__o211a_1 _19210_ (.A1(\rbzero.spi_registers.buf_texadd2[16] ),
    .A2(_03049_),
    .B1(_03058_),
    .C1(_03056_),
    .X(_00895_));
 sky130_fd_sc_hd__or2_1 _19211_ (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .B(_03050_),
    .X(_03059_));
 sky130_fd_sc_hd__o211a_1 _19212_ (.A1(\rbzero.spi_registers.buf_texadd2[17] ),
    .A2(_03049_),
    .B1(_03059_),
    .C1(_03056_),
    .X(_00896_));
 sky130_fd_sc_hd__or2_1 _19213_ (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .B(_03050_),
    .X(_03060_));
 sky130_fd_sc_hd__o211a_1 _19214_ (.A1(\rbzero.spi_registers.buf_texadd2[18] ),
    .A2(_03049_),
    .B1(_03060_),
    .C1(_03056_),
    .X(_00897_));
 sky130_fd_sc_hd__or2_1 _19215_ (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .B(_03050_),
    .X(_03061_));
 sky130_fd_sc_hd__o211a_1 _19216_ (.A1(\rbzero.spi_registers.buf_texadd2[19] ),
    .A2(_03049_),
    .B1(_03061_),
    .C1(_03056_),
    .X(_00898_));
 sky130_fd_sc_hd__or2_1 _19217_ (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .B(_03036_),
    .X(_03062_));
 sky130_fd_sc_hd__o211a_1 _19218_ (.A1(\rbzero.spi_registers.buf_texadd2[20] ),
    .A2(_03034_),
    .B1(_03062_),
    .C1(_03056_),
    .X(_00899_));
 sky130_fd_sc_hd__or2_1 _19219_ (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .B(_03036_),
    .X(_03063_));
 sky130_fd_sc_hd__o211a_1 _19220_ (.A1(\rbzero.spi_registers.buf_texadd2[21] ),
    .A2(_03034_),
    .B1(_03063_),
    .C1(_03056_),
    .X(_00900_));
 sky130_fd_sc_hd__or2_1 _19221_ (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .B(_03036_),
    .X(_03064_));
 sky130_fd_sc_hd__o211a_1 _19222_ (.A1(\rbzero.spi_registers.buf_texadd2[22] ),
    .A2(_03034_),
    .B1(_03064_),
    .C1(_03056_),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _19223_ (.A(\rbzero.spi_registers.spi_buffer[23] ),
    .B(_03036_),
    .X(_03065_));
 sky130_fd_sc_hd__o211a_1 _19224_ (.A1(\rbzero.spi_registers.buf_texadd2[23] ),
    .A2(_03034_),
    .B1(_03065_),
    .C1(_03056_),
    .X(_00902_));
 sky130_fd_sc_hd__and3_1 _19225_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02376_),
    .C(_02378_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_2 _19226_ (.A(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_4 _19227_ (.A(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__nand3_2 _19228_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02376_),
    .C(_02378_),
    .Y(_03069_));
 sky130_fd_sc_hd__buf_2 _19229_ (.A(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__or2_1 _19230_ (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .B(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__buf_2 _19231_ (.A(_02997_),
    .X(_03072_));
 sky130_fd_sc_hd__o211a_1 _19232_ (.A1(\rbzero.spi_registers.buf_texadd3[0] ),
    .A2(_03068_),
    .B1(_03071_),
    .C1(_03072_),
    .X(_00903_));
 sky130_fd_sc_hd__or2_1 _19233_ (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .B(_03070_),
    .X(_03073_));
 sky130_fd_sc_hd__o211a_1 _19234_ (.A1(\rbzero.spi_registers.buf_texadd3[1] ),
    .A2(_03068_),
    .B1(_03073_),
    .C1(_03072_),
    .X(_00904_));
 sky130_fd_sc_hd__or2_1 _19235_ (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .B(_03070_),
    .X(_03074_));
 sky130_fd_sc_hd__o211a_1 _19236_ (.A1(\rbzero.spi_registers.buf_texadd3[2] ),
    .A2(_03068_),
    .B1(_03074_),
    .C1(_03072_),
    .X(_00905_));
 sky130_fd_sc_hd__or2_1 _19237_ (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .B(_03070_),
    .X(_03075_));
 sky130_fd_sc_hd__o211a_1 _19238_ (.A1(\rbzero.spi_registers.buf_texadd3[3] ),
    .A2(_03068_),
    .B1(_03075_),
    .C1(_03072_),
    .X(_00906_));
 sky130_fd_sc_hd__or2_1 _19239_ (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .B(_03070_),
    .X(_03076_));
 sky130_fd_sc_hd__o211a_1 _19240_ (.A1(\rbzero.spi_registers.buf_texadd3[4] ),
    .A2(_03068_),
    .B1(_03076_),
    .C1(_03072_),
    .X(_00907_));
 sky130_fd_sc_hd__or2_1 _19241_ (.A(_02648_),
    .B(_03070_),
    .X(_03077_));
 sky130_fd_sc_hd__o211a_1 _19242_ (.A1(\rbzero.spi_registers.buf_texadd3[5] ),
    .A2(_03068_),
    .B1(_03077_),
    .C1(_03072_),
    .X(_00908_));
 sky130_fd_sc_hd__or2_1 _19243_ (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .B(_03070_),
    .X(_03078_));
 sky130_fd_sc_hd__o211a_1 _19244_ (.A1(\rbzero.spi_registers.buf_texadd3[6] ),
    .A2(_03068_),
    .B1(_03078_),
    .C1(_03072_),
    .X(_00909_));
 sky130_fd_sc_hd__or2_1 _19245_ (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .B(_03070_),
    .X(_03079_));
 sky130_fd_sc_hd__o211a_1 _19246_ (.A1(\rbzero.spi_registers.buf_texadd3[7] ),
    .A2(_03068_),
    .B1(_03079_),
    .C1(_03072_),
    .X(_00910_));
 sky130_fd_sc_hd__or2_1 _19247_ (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .B(_03070_),
    .X(_03080_));
 sky130_fd_sc_hd__o211a_1 _19248_ (.A1(\rbzero.spi_registers.buf_texadd3[8] ),
    .A2(_03068_),
    .B1(_03080_),
    .C1(_03072_),
    .X(_00911_));
 sky130_fd_sc_hd__or2_1 _19249_ (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .B(_03070_),
    .X(_03081_));
 sky130_fd_sc_hd__o211a_1 _19250_ (.A1(\rbzero.spi_registers.buf_texadd3[9] ),
    .A2(_03068_),
    .B1(_03081_),
    .C1(_03072_),
    .X(_00912_));
 sky130_fd_sc_hd__buf_2 _19251_ (.A(_03067_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_2 _19252_ (.A(_03069_),
    .X(_03083_));
 sky130_fd_sc_hd__or2_1 _19253_ (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .B(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__buf_2 _19254_ (.A(_02997_),
    .X(_03085_));
 sky130_fd_sc_hd__o211a_1 _19255_ (.A1(\rbzero.spi_registers.buf_texadd3[10] ),
    .A2(_03082_),
    .B1(_03084_),
    .C1(_03085_),
    .X(_00913_));
 sky130_fd_sc_hd__or2_1 _19256_ (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .B(_03083_),
    .X(_03086_));
 sky130_fd_sc_hd__o211a_1 _19257_ (.A1(\rbzero.spi_registers.buf_texadd3[11] ),
    .A2(_03082_),
    .B1(_03086_),
    .C1(_03085_),
    .X(_00914_));
 sky130_fd_sc_hd__or2_1 _19258_ (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .B(_03083_),
    .X(_03087_));
 sky130_fd_sc_hd__o211a_1 _19259_ (.A1(\rbzero.spi_registers.buf_texadd3[12] ),
    .A2(_03082_),
    .B1(_03087_),
    .C1(_03085_),
    .X(_00915_));
 sky130_fd_sc_hd__or2_1 _19260_ (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .B(_03083_),
    .X(_03088_));
 sky130_fd_sc_hd__o211a_1 _19261_ (.A1(\rbzero.spi_registers.buf_texadd3[13] ),
    .A2(_03082_),
    .B1(_03088_),
    .C1(_03085_),
    .X(_00916_));
 sky130_fd_sc_hd__or2_1 _19262_ (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .B(_03083_),
    .X(_03089_));
 sky130_fd_sc_hd__o211a_1 _19263_ (.A1(\rbzero.spi_registers.buf_texadd3[14] ),
    .A2(_03082_),
    .B1(_03089_),
    .C1(_03085_),
    .X(_00917_));
 sky130_fd_sc_hd__or2_1 _19264_ (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .B(_03083_),
    .X(_03090_));
 sky130_fd_sc_hd__o211a_1 _19265_ (.A1(\rbzero.spi_registers.buf_texadd3[15] ),
    .A2(_03082_),
    .B1(_03090_),
    .C1(_03085_),
    .X(_00918_));
 sky130_fd_sc_hd__or2_1 _19266_ (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .B(_03083_),
    .X(_03091_));
 sky130_fd_sc_hd__o211a_1 _19267_ (.A1(\rbzero.spi_registers.buf_texadd3[16] ),
    .A2(_03082_),
    .B1(_03091_),
    .C1(_03085_),
    .X(_00919_));
 sky130_fd_sc_hd__or2_1 _19268_ (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .B(_03083_),
    .X(_03092_));
 sky130_fd_sc_hd__o211a_1 _19269_ (.A1(\rbzero.spi_registers.buf_texadd3[17] ),
    .A2(_03082_),
    .B1(_03092_),
    .C1(_03085_),
    .X(_00920_));
 sky130_fd_sc_hd__or2_1 _19270_ (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .B(_03083_),
    .X(_03093_));
 sky130_fd_sc_hd__o211a_1 _19271_ (.A1(\rbzero.spi_registers.buf_texadd3[18] ),
    .A2(_03082_),
    .B1(_03093_),
    .C1(_03085_),
    .X(_00921_));
 sky130_fd_sc_hd__or2_1 _19272_ (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .B(_03083_),
    .X(_03094_));
 sky130_fd_sc_hd__o211a_1 _19273_ (.A1(\rbzero.spi_registers.buf_texadd3[19] ),
    .A2(_03082_),
    .B1(_03094_),
    .C1(_03085_),
    .X(_00922_));
 sky130_fd_sc_hd__or2_1 _19274_ (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .B(_03069_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_4 _19275_ (.A(_02997_),
    .X(_03096_));
 sky130_fd_sc_hd__o211a_1 _19276_ (.A1(\rbzero.spi_registers.buf_texadd3[20] ),
    .A2(_03067_),
    .B1(_03095_),
    .C1(_03096_),
    .X(_00923_));
 sky130_fd_sc_hd__or2_1 _19277_ (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .B(_03069_),
    .X(_03097_));
 sky130_fd_sc_hd__o211a_1 _19278_ (.A1(\rbzero.spi_registers.buf_texadd3[21] ),
    .A2(_03067_),
    .B1(_03097_),
    .C1(_03096_),
    .X(_00924_));
 sky130_fd_sc_hd__or2_1 _19279_ (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .B(_03069_),
    .X(_03098_));
 sky130_fd_sc_hd__o211a_1 _19280_ (.A1(\rbzero.spi_registers.buf_texadd3[22] ),
    .A2(_03067_),
    .B1(_03098_),
    .C1(_03096_),
    .X(_00925_));
 sky130_fd_sc_hd__or2_1 _19281_ (.A(\rbzero.spi_registers.spi_buffer[23] ),
    .B(_03069_),
    .X(_03099_));
 sky130_fd_sc_hd__o211a_1 _19282_ (.A1(\rbzero.spi_registers.buf_texadd3[23] ),
    .A2(_03067_),
    .B1(_03099_),
    .C1(_03096_),
    .X(_00926_));
 sky130_fd_sc_hd__nand2_2 _19283_ (.A(_02390_),
    .B(_02400_),
    .Y(_03100_));
 sky130_fd_sc_hd__mux2_1 _19284_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.spi_cmd[0] ),
    .S(_03100_),
    .X(_03101_));
 sky130_fd_sc_hd__and2_1 _19285_ (.A(_02621_),
    .B(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _19286_ (.A(_03102_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19287_ (.A0(\rbzero.spi_registers.spi_cmd[0] ),
    .A1(\rbzero.spi_registers.spi_cmd[1] ),
    .S(_03100_),
    .X(_03103_));
 sky130_fd_sc_hd__and2_1 _19288_ (.A(_02621_),
    .B(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _19289_ (.A(_03104_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _19290_ (.A0(\rbzero.spi_registers.spi_cmd[1] ),
    .A1(\rbzero.spi_registers.spi_cmd[2] ),
    .S(_03100_),
    .X(_03105_));
 sky130_fd_sc_hd__and2_1 _19291_ (.A(_02621_),
    .B(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _19292_ (.A(_03106_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19293_ (.A0(\rbzero.spi_registers.spi_cmd[2] ),
    .A1(\rbzero.spi_registers.spi_cmd[3] ),
    .S(_03100_),
    .X(_03107_));
 sky130_fd_sc_hd__and2_1 _19294_ (.A(_02621_),
    .B(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _19295_ (.A(_03108_),
    .X(_00930_));
 sky130_fd_sc_hd__and2_1 _19296_ (.A(net55),
    .B(_09712_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _19297_ (.A(_03109_),
    .X(_00931_));
 sky130_fd_sc_hd__and2_1 _19298_ (.A(\rbzero.pov.ss_buffer[0] ),
    .B(_09712_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _19299_ (.A(_03110_),
    .X(_00932_));
 sky130_fd_sc_hd__clkbuf_4 _19300_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_03111_));
 sky130_fd_sc_hd__nor2_1 _19301_ (.A(_03111_),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2_1 _19302_ (.A(_03111_),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_03113_));
 sky130_fd_sc_hd__or2b_1 _19303_ (.A(_03112_),
    .B_N(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__or2_1 _19304_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .X(_03115_));
 sky130_fd_sc_hd__nor2_1 _19305_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_03116_));
 sky130_fd_sc_hd__nand2_1 _19306_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_03117_));
 sky130_fd_sc_hd__or2_1 _19307_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_03118_));
 sky130_fd_sc_hd__nand4_1 _19308_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .C(_03117_),
    .D(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__and2_1 _19309_ (.A(_03117_),
    .B(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__nand2_1 _19310_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_03121_));
 sky130_fd_sc_hd__o21ai_1 _19311_ (.A1(_03116_),
    .A2(_03120_),
    .B1(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_1 _19312_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .Y(_03123_));
 sky130_fd_sc_hd__a21boi_1 _19313_ (.A1(_03115_),
    .A2(_03122_),
    .B1_N(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__xnor2_1 _19314_ (.A(_03114_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__nor2_1 _19315_ (.A(_09731_),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__a221o_1 _19316_ (.A1(_05282_),
    .A2(_08113_),
    .B1(_02406_),
    .B2(\rbzero.wall_tracer.rayAddendY[-5] ),
    .C1(_03126_),
    .X(_00933_));
 sky130_fd_sc_hd__clkbuf_4 _19317_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_03127_));
 sky130_fd_sc_hd__or2_1 _19318_ (.A(_03127_),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_03128_));
 sky130_fd_sc_hd__nand2_1 _19319_ (.A(_03127_),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .Y(_03129_));
 sky130_fd_sc_hd__o21ai_1 _19320_ (.A1(_03112_),
    .A2(_03124_),
    .B1(_03113_),
    .Y(_03130_));
 sky130_fd_sc_hd__and3_1 _19321_ (.A(_03128_),
    .B(_03129_),
    .C(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__a21oi_1 _19322_ (.A1(_03128_),
    .A2(_03129_),
    .B1(_03130_),
    .Y(_03132_));
 sky130_fd_sc_hd__o21ai_1 _19323_ (.A1(_03131_),
    .A2(_03132_),
    .B1(_04478_),
    .Y(_03133_));
 sky130_fd_sc_hd__nand2_1 _19324_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_05282_),
    .Y(_03134_));
 sky130_fd_sc_hd__or2_1 _19325_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_05282_),
    .X(_03135_));
 sky130_fd_sc_hd__a31o_1 _19326_ (.A1(_02425_),
    .A2(_03134_),
    .A3(_03135_),
    .B1(_09727_),
    .X(_03136_));
 sky130_fd_sc_hd__a22o_1 _19327_ (.A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_09738_),
    .B1(_03133_),
    .B2(_03136_),
    .X(_00934_));
 sky130_fd_sc_hd__nor2_1 _19328_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_03137_));
 sky130_fd_sc_hd__and2_1 _19329_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .X(_03138_));
 sky130_fd_sc_hd__a21o_1 _19330_ (.A1(_03127_),
    .A2(\rbzero.wall_tracer.rayAddendY[-4] ),
    .B1(_03130_),
    .X(_03139_));
 sky130_fd_sc_hd__o21ai_1 _19331_ (.A1(_03127_),
    .A2(\rbzero.wall_tracer.rayAddendY[-4] ),
    .B1(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__o21ai_1 _19332_ (.A1(_03137_),
    .A2(_03138_),
    .B1(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__o311a_1 _19333_ (.A1(_03137_),
    .A2(_03138_),
    .A3(_03140_),
    .B1(_03141_),
    .C1(_04469_),
    .X(_03142_));
 sky130_fd_sc_hd__or2_1 _19334_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03135_),
    .X(_03143_));
 sky130_fd_sc_hd__nand2_1 _19335_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03135_),
    .Y(_03144_));
 sky130_fd_sc_hd__a31o_1 _19336_ (.A1(_02439_),
    .A2(_03143_),
    .A3(_03144_),
    .B1(_09724_),
    .X(_03145_));
 sky130_fd_sc_hd__o22a_1 _19337_ (.A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A2(_02432_),
    .B1(_03142_),
    .B2(_03145_),
    .X(_00935_));
 sky130_fd_sc_hd__nor2_1 _19338_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_03146_));
 sky130_fd_sc_hd__and2_1 _19339_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_03147_));
 sky130_fd_sc_hd__nand2_1 _19340_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_03148_));
 sky130_fd_sc_hd__o21ai_1 _19341_ (.A1(_03137_),
    .A2(_03140_),
    .B1(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__or3_1 _19342_ (.A(_03146_),
    .B(_03147_),
    .C(_03149_),
    .X(_03150_));
 sky130_fd_sc_hd__o21ai_1 _19343_ (.A1(_03146_),
    .A2(_03147_),
    .B1(_03149_),
    .Y(_03151_));
 sky130_fd_sc_hd__a21oi_1 _19344_ (.A1(_03150_),
    .A2(_03151_),
    .B1(_08113_),
    .Y(_03152_));
 sky130_fd_sc_hd__nand2_1 _19345_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_03143_),
    .Y(_03153_));
 sky130_fd_sc_hd__or2_1 _19346_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .B(_03143_),
    .X(_03154_));
 sky130_fd_sc_hd__a31o_1 _19347_ (.A1(_02439_),
    .A2(_03153_),
    .A3(_03154_),
    .B1(_02405_),
    .X(_03155_));
 sky130_fd_sc_hd__o22a_1 _19348_ (.A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A2(_02432_),
    .B1(_03152_),
    .B2(_03155_),
    .X(_00936_));
 sky130_fd_sc_hd__or2_1 _19349_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_03156_));
 sky130_fd_sc_hd__nand2_1 _19350_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_03157_));
 sky130_fd_sc_hd__nor2_1 _19351_ (.A(_03147_),
    .B(_03149_),
    .Y(_03158_));
 sky130_fd_sc_hd__nor2_1 _19352_ (.A(_03146_),
    .B(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__a21oi_1 _19353_ (.A1(_03156_),
    .A2(_03157_),
    .B1(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__a31o_1 _19354_ (.A1(_03156_),
    .A2(_03157_),
    .A3(_03159_),
    .B1(_09730_),
    .X(_03161_));
 sky130_fd_sc_hd__inv_2 _19355_ (.A(_05282_),
    .Y(_03162_));
 sky130_fd_sc_hd__o31a_1 _19356_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(\rbzero.debug_overlay.vplaneY[-7] ),
    .A3(\rbzero.debug_overlay.vplaneY[-8] ),
    .B1(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__xnor2_1 _19357_ (.A(_03111_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__o2bb2a_1 _19358_ (.A1_N(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A2_N(_02405_),
    .B1(_03164_),
    .B2(_04469_),
    .X(_03165_));
 sky130_fd_sc_hd__o21ai_1 _19359_ (.A1(_03160_),
    .A2(_03161_),
    .B1(_03165_),
    .Y(_00937_));
 sky130_fd_sc_hd__a21bo_1 _19360_ (.A1(_03156_),
    .A2(_03159_),
    .B1_N(_03157_),
    .X(_03166_));
 sky130_fd_sc_hd__clkbuf_4 _19361_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_03167_));
 sky130_fd_sc_hd__nor2_1 _19362_ (.A(_03167_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_03168_));
 sky130_fd_sc_hd__and2_1 _19363_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_03169_));
 sky130_fd_sc_hd__or2_1 _19364_ (.A(_03168_),
    .B(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__xnor2_1 _19365_ (.A(_03166_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__or2_1 _19366_ (.A(_03127_),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_03172_));
 sky130_fd_sc_hd__nand2_1 _19367_ (.A(_03127_),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_03173_));
 sky130_fd_sc_hd__nand2_1 _19368_ (.A(_03172_),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__nor2_1 _19369_ (.A(_03111_),
    .B(_03154_),
    .Y(_03175_));
 sky130_fd_sc_hd__a21oi_1 _19370_ (.A1(_03111_),
    .A2(_05282_),
    .B1(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__xnor2_1 _19371_ (.A(_03174_),
    .B(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__mux2_1 _19372_ (.A0(_03171_),
    .A1(_03177_),
    .S(_08112_),
    .X(_03178_));
 sky130_fd_sc_hd__mux2_1 _19373_ (.A0(\rbzero.wall_tracer.rayAddendY[0] ),
    .A1(_03178_),
    .S(_02431_),
    .X(_03179_));
 sky130_fd_sc_hd__clkbuf_1 _19374_ (.A(_03179_),
    .X(_00938_));
 sky130_fd_sc_hd__nand2_1 _19375_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_03180_));
 sky130_fd_sc_hd__or2_1 _19376_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_03181_));
 sky130_fd_sc_hd__o21a_1 _19377_ (.A1(_03167_),
    .A2(\rbzero.wall_tracer.rayAddendY[0] ),
    .B1(_03166_),
    .X(_03182_));
 sky130_fd_sc_hd__a211o_1 _19378_ (.A1(_03180_),
    .A2(_03181_),
    .B1(_03182_),
    .C1(_03169_),
    .X(_03183_));
 sky130_fd_sc_hd__o211ai_2 _19379_ (.A1(_03169_),
    .A2(_03182_),
    .B1(_03181_),
    .C1(_03180_),
    .Y(_03184_));
 sky130_fd_sc_hd__a21oi_1 _19380_ (.A1(_03111_),
    .A2(_05282_),
    .B1(_03174_),
    .Y(_03185_));
 sky130_fd_sc_hd__nor2_1 _19381_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_03186_));
 sky130_fd_sc_hd__and2_1 _19382_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(_03187_));
 sky130_fd_sc_hd__nor2_1 _19383_ (.A(_03186_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__xnor2_1 _19384_ (.A(_03172_),
    .B(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__o21a_1 _19385_ (.A1(_03175_),
    .A2(_03185_),
    .B1(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__inv_2 _19386_ (.A(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__or3_1 _19387_ (.A(_03175_),
    .B(_03189_),
    .C(_03185_),
    .X(_03192_));
 sky130_fd_sc_hd__a32o_1 _19388_ (.A1(_02425_),
    .A2(_03191_),
    .A3(_03192_),
    .B1(_02406_),
    .B2(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_03193_));
 sky130_fd_sc_hd__a31o_1 _19389_ (.A1(_02478_),
    .A2(_03183_),
    .A3(_03184_),
    .B1(_03193_),
    .X(_00939_));
 sky130_fd_sc_hd__buf_2 _19390_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_03194_));
 sky130_fd_sc_hd__buf_2 _19391_ (.A(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_4 _19392_ (.A(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__xnor2_1 _19393_ (.A(_03196_),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_03197_));
 sky130_fd_sc_hd__a21oi_1 _19394_ (.A1(_03180_),
    .A2(_03184_),
    .B1(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__a311oi_1 _19395_ (.A1(_03180_),
    .A2(_03184_),
    .A3(_03197_),
    .B1(_03198_),
    .C1(_08113_),
    .Y(_03199_));
 sky130_fd_sc_hd__xor2_1 _19396_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_03200_));
 sky130_fd_sc_hd__o31ai_1 _19397_ (.A1(_03172_),
    .A2(_03186_),
    .A3(_03187_),
    .B1(_03191_),
    .Y(_03201_));
 sky130_fd_sc_hd__xnor2_1 _19398_ (.A(_03200_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__xnor2_1 _19399_ (.A(_03186_),
    .B(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__a21o_1 _19400_ (.A1(_08113_),
    .A2(_03203_),
    .B1(_02406_),
    .X(_03204_));
 sky130_fd_sc_hd__o22a_1 _19401_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(_02432_),
    .B1(_03199_),
    .B2(_03204_),
    .X(_00940_));
 sky130_fd_sc_hd__and2_1 _19402_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_03205_));
 sky130_fd_sc_hd__nor2_1 _19403_ (.A(_03194_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_03206_));
 sky130_fd_sc_hd__o21ai_1 _19404_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(_03194_),
    .Y(_03207_));
 sky130_fd_sc_hd__o21bai_1 _19405_ (.A1(_03194_),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1_N(_03184_),
    .Y(_03208_));
 sky130_fd_sc_hd__o211ai_1 _19406_ (.A1(_03205_),
    .A2(_03206_),
    .B1(_03207_),
    .C1(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__a211o_1 _19407_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03205_),
    .C1(_03206_),
    .X(_03210_));
 sky130_fd_sc_hd__or2_1 _19408_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_03111_),
    .X(_03211_));
 sky130_fd_sc_hd__nand2_1 _19409_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_03111_),
    .Y(_03212_));
 sky130_fd_sc_hd__and4bb_1 _19410_ (.A_N(\rbzero.debug_overlay.vplaneY[-2] ),
    .B_N(\rbzero.debug_overlay.vplaneY[-6] ),
    .C(_03211_),
    .D(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__a2bb2o_1 _19411_ (.A1_N(\rbzero.debug_overlay.vplaneY[-2] ),
    .A2_N(\rbzero.debug_overlay.vplaneY[-6] ),
    .B1(_03211_),
    .B2(_03212_),
    .X(_03214_));
 sky130_fd_sc_hd__and2b_1 _19412_ (.A_N(_03213_),
    .B(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__o21a_1 _19413_ (.A1(_03190_),
    .A2(_03200_),
    .B1(_03186_),
    .X(_03216_));
 sky130_fd_sc_hd__a21o_1 _19414_ (.A1(_03200_),
    .A2(_03201_),
    .B1(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__and2_1 _19415_ (.A(_03215_),
    .B(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__o21ai_1 _19416_ (.A1(_03215_),
    .A2(_03217_),
    .B1(_02425_),
    .Y(_03219_));
 sky130_fd_sc_hd__a2bb2o_1 _19417_ (.A1_N(_03218_),
    .A2_N(_03219_),
    .B1(\rbzero.wall_tracer.rayAddendY[3] ),
    .B2(_02405_),
    .X(_03220_));
 sky130_fd_sc_hd__a31o_1 _19418_ (.A1(_02478_),
    .A2(_03209_),
    .A3(_03210_),
    .B1(_03220_),
    .X(_00941_));
 sky130_fd_sc_hd__nand2_1 _19419_ (.A(_03196_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_03221_));
 sky130_fd_sc_hd__xor2_1 _19420_ (.A(_03194_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_03222_));
 sky130_fd_sc_hd__a21oi_1 _19421_ (.A1(_03221_),
    .A2(_03210_),
    .B1(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__a31o_1 _19422_ (.A1(_03221_),
    .A2(_03210_),
    .A3(_03222_),
    .B1(_08111_),
    .X(_03224_));
 sky130_fd_sc_hd__nor2_1 _19423_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_03111_),
    .Y(_03225_));
 sky130_fd_sc_hd__xor2_1 _19424_ (.A(_03167_),
    .B(_03127_),
    .X(_03226_));
 sky130_fd_sc_hd__or2_1 _19425_ (.A(_03213_),
    .B(_03218_),
    .X(_03227_));
 sky130_fd_sc_hd__xnor2_1 _19426_ (.A(_03226_),
    .B(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__xnor2_1 _19427_ (.A(_03225_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__o22a_1 _19428_ (.A1(_03223_),
    .A2(_03224_),
    .B1(_03229_),
    .B2(_04469_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _19429_ (.A0(\rbzero.wall_tracer.rayAddendY[4] ),
    .A1(_03230_),
    .S(_02431_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_1 _19430_ (.A(_03231_),
    .X(_00942_));
 sky130_fd_sc_hd__nand2_1 _19431_ (.A(_03194_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_03232_));
 sky130_fd_sc_hd__or2_1 _19432_ (.A(_03194_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_03233_));
 sky130_fd_sc_hd__nand2_1 _19433_ (.A(_03232_),
    .B(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__or2b_1 _19434_ (.A(_03210_),
    .B_N(_03222_),
    .X(_03235_));
 sky130_fd_sc_hd__o21ai_1 _19435_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_03196_),
    .Y(_03236_));
 sky130_fd_sc_hd__nand3_1 _19436_ (.A(_03234_),
    .B(_03235_),
    .C(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__a21o_1 _19437_ (.A1(_03235_),
    .A2(_03236_),
    .B1(_03234_),
    .X(_03238_));
 sky130_fd_sc_hd__nor2_1 _19438_ (.A(_03194_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .Y(_03239_));
 sky130_fd_sc_hd__and2_1 _19439_ (.A(_03194_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_03240_));
 sky130_fd_sc_hd__o22a_1 _19440_ (.A1(_03167_),
    .A2(_03127_),
    .B1(_03239_),
    .B2(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__nor4_1 _19441_ (.A(_03167_),
    .B(_03127_),
    .C(_03239_),
    .D(_03240_),
    .Y(_03242_));
 sky130_fd_sc_hd__nor2_1 _19442_ (.A(_03241_),
    .B(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__o21a_1 _19443_ (.A1(_03218_),
    .A2(_03226_),
    .B1(_03225_),
    .X(_03244_));
 sky130_fd_sc_hd__a21oi_1 _19444_ (.A1(_03226_),
    .A2(_03227_),
    .B1(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__xnor2_1 _19445_ (.A(_03243_),
    .B(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__a22o_1 _19446_ (.A1(\rbzero.wall_tracer.rayAddendY[5] ),
    .A2(_02405_),
    .B1(_03246_),
    .B2(_02439_),
    .X(_03247_));
 sky130_fd_sc_hd__a31o_1 _19447_ (.A1(_02478_),
    .A2(_03237_),
    .A3(_03238_),
    .B1(_03247_),
    .X(_00943_));
 sky130_fd_sc_hd__xnor2_1 _19448_ (.A(_03195_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_03248_));
 sky130_fd_sc_hd__a21oi_1 _19449_ (.A1(_03232_),
    .A2(_03238_),
    .B1(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__a31o_1 _19450_ (.A1(_03232_),
    .A2(_03238_),
    .A3(_03248_),
    .B1(_08111_),
    .X(_03250_));
 sky130_fd_sc_hd__or2_1 _19451_ (.A(_03194_),
    .B(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_03251_));
 sky130_fd_sc_hd__nand2_1 _19452_ (.A(_03195_),
    .B(\rbzero.debug_overlay.vplaneY[-2] ),
    .Y(_03252_));
 sky130_fd_sc_hd__a21o_1 _19453_ (.A1(_03251_),
    .A2(_03252_),
    .B1(_03239_),
    .X(_03253_));
 sky130_fd_sc_hd__nand2_1 _19454_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(_03239_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand2_1 _19455_ (.A(_03253_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__o21bai_1 _19456_ (.A1(_03241_),
    .A2(_03245_),
    .B1_N(_03242_),
    .Y(_03256_));
 sky130_fd_sc_hd__xnor2_1 _19457_ (.A(_03255_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__a2bb2o_1 _19458_ (.A1_N(_03249_),
    .A2_N(_03250_),
    .B1(_03257_),
    .B2(_08112_),
    .X(_03258_));
 sky130_fd_sc_hd__mux2_1 _19459_ (.A0(\rbzero.wall_tracer.rayAddendY[6] ),
    .A1(_03258_),
    .S(_02431_),
    .X(_03259_));
 sky130_fd_sc_hd__clkbuf_1 _19460_ (.A(_03259_),
    .X(_00944_));
 sky130_fd_sc_hd__nor3_1 _19461_ (.A(_03234_),
    .B(_03235_),
    .C(_03248_),
    .Y(_03260_));
 sky130_fd_sc_hd__o41a_1 _19462_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[5] ),
    .A3(\rbzero.wall_tracer.rayAddendY[4] ),
    .A4(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_03195_),
    .X(_03261_));
 sky130_fd_sc_hd__nand2_1 _19463_ (.A(_03195_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_03262_));
 sky130_fd_sc_hd__or2_1 _19464_ (.A(_03195_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_03263_));
 sky130_fd_sc_hd__o211ai_2 _19465_ (.A1(_03260_),
    .A2(_03261_),
    .B1(_03262_),
    .C1(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__a211o_1 _19466_ (.A1(_03262_),
    .A2(_03263_),
    .B1(_03260_),
    .C1(_03261_),
    .X(_03265_));
 sky130_fd_sc_hd__inv_2 _19467_ (.A(_03254_),
    .Y(_03266_));
 sky130_fd_sc_hd__and3_1 _19468_ (.A(_03253_),
    .B(_03254_),
    .C(_03256_),
    .X(_03267_));
 sky130_fd_sc_hd__nor2_1 _19469_ (.A(_03195_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .Y(_03268_));
 sky130_fd_sc_hd__and2_1 _19470_ (.A(_03195_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_03269_));
 sky130_fd_sc_hd__o21ai_1 _19471_ (.A1(_03268_),
    .A2(_03269_),
    .B1(_03251_),
    .Y(_03270_));
 sky130_fd_sc_hd__or3_1 _19472_ (.A(_03251_),
    .B(_03268_),
    .C(_03269_),
    .X(_03271_));
 sky130_fd_sc_hd__o211ai_2 _19473_ (.A1(_03266_),
    .A2(_03267_),
    .B1(_03270_),
    .C1(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__a211o_1 _19474_ (.A1(_03270_),
    .A2(_03271_),
    .B1(_03266_),
    .C1(_03267_),
    .X(_03273_));
 sky130_fd_sc_hd__a32o_1 _19475_ (.A1(_02425_),
    .A2(_03272_),
    .A3(_03273_),
    .B1(_02406_),
    .B2(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_03274_));
 sky130_fd_sc_hd__a31o_1 _19476_ (.A1(_02478_),
    .A2(_03264_),
    .A3(_03265_),
    .B1(_03274_),
    .X(_00945_));
 sky130_fd_sc_hd__xnor2_1 _19477_ (.A(_03195_),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_03275_));
 sky130_fd_sc_hd__a21oi_1 _19478_ (.A1(_03262_),
    .A2(_03264_),
    .B1(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__a31o_1 _19479_ (.A1(_03262_),
    .A2(_03264_),
    .A3(_03275_),
    .B1(_08112_),
    .X(_03277_));
 sky130_fd_sc_hd__nor2_1 _19480_ (.A(_03276_),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__inv_2 _19481_ (.A(_03167_),
    .Y(_03279_));
 sky130_fd_sc_hd__a21oi_1 _19482_ (.A1(_03167_),
    .A2(\rbzero.debug_overlay.vplaneY[-1] ),
    .B1(_03195_),
    .Y(_03280_));
 sky130_fd_sc_hd__a21oi_1 _19483_ (.A1(_03196_),
    .A2(_03167_),
    .B1(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__a21oi_1 _19484_ (.A1(_03279_),
    .A2(_03268_),
    .B1(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__a21o_1 _19485_ (.A1(_03271_),
    .A2(_03272_),
    .B1(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__nand3_1 _19486_ (.A(_03271_),
    .B(_03272_),
    .C(_03282_),
    .Y(_03284_));
 sky130_fd_sc_hd__a31o_1 _19487_ (.A1(_02425_),
    .A2(_03283_),
    .A3(_03284_),
    .B1(_02405_),
    .X(_03285_));
 sky130_fd_sc_hd__o22a_1 _19488_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(_02432_),
    .B1(_03278_),
    .B2(_03285_),
    .X(_00946_));
 sky130_fd_sc_hd__or2_1 _19489_ (.A(_03196_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_03286_));
 sky130_fd_sc_hd__nand2_1 _19490_ (.A(_03196_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2_1 _19491_ (.A(_03286_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__o21ai_1 _19492_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(\rbzero.wall_tracer.rayAddendY[7] ),
    .B1(_03196_),
    .Y(_03289_));
 sky130_fd_sc_hd__o21ai_1 _19493_ (.A1(_03264_),
    .A2(_03275_),
    .B1(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__xnor2_1 _19494_ (.A(_03288_),
    .B(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__inv_2 _19495_ (.A(_03196_),
    .Y(_03292_));
 sky130_fd_sc_hd__a21oi_1 _19496_ (.A1(_03292_),
    .A2(_03279_),
    .B1(_03283_),
    .Y(_03293_));
 sky130_fd_sc_hd__a211o_1 _19497_ (.A1(_03280_),
    .A2(_03283_),
    .B1(_03293_),
    .C1(_04469_),
    .X(_03294_));
 sky130_fd_sc_hd__o221a_1 _19498_ (.A1(\rbzero.wall_tracer.rayAddendY[9] ),
    .A2(_02432_),
    .B1(_09731_),
    .B2(_03291_),
    .C1(_03294_),
    .X(_00947_));
 sky130_fd_sc_hd__a21bo_1 _19499_ (.A1(_03286_),
    .A2(_03290_),
    .B1_N(_03287_),
    .X(_03295_));
 sky130_fd_sc_hd__xnor2_1 _19500_ (.A(_03196_),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_03296_));
 sky130_fd_sc_hd__xnor2_1 _19501_ (.A(_03295_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__o211a_1 _19502_ (.A1(_03167_),
    .A2(_03283_),
    .B1(_08112_),
    .C1(_03292_),
    .X(_03298_));
 sky130_fd_sc_hd__o22a_1 _19503_ (.A1(_02439_),
    .A2(_03297_),
    .B1(_03298_),
    .B2(_09728_),
    .X(_03299_));
 sky130_fd_sc_hd__a21o_1 _19504_ (.A1(\rbzero.wall_tracer.rayAddendY[10] ),
    .A2(_09725_),
    .B1(_03299_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _19505_ (.A0(\rbzero.debug_overlay.playerX[0] ),
    .A1(_06164_),
    .S(_09784_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _19506_ (.A0(_06108_),
    .A1(_03300_),
    .S(_09826_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_1 _19507_ (.A(_03301_),
    .X(_00949_));
 sky130_fd_sc_hd__nor2_1 _19508_ (.A(_06108_),
    .B(_09745_),
    .Y(_03302_));
 sky130_fd_sc_hd__or3_1 _19509_ (.A(_06102_),
    .B(_09746_),
    .C(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__o211a_1 _19510_ (.A1(_04998_),
    .A2(_08101_),
    .B1(_09826_),
    .C1(_03303_),
    .X(_03304_));
 sky130_fd_sc_hd__a21oi_1 _19511_ (.A1(_06122_),
    .A2(_09763_),
    .B1(_03304_),
    .Y(_00950_));
 sky130_fd_sc_hd__xnor2_1 _19512_ (.A(_09747_),
    .B(_09750_),
    .Y(_03305_));
 sky130_fd_sc_hd__or2_1 _19513_ (.A(_09824_),
    .B(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__o211a_1 _19514_ (.A1(_05000_),
    .A2(_08101_),
    .B1(_09826_),
    .C1(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__a21oi_1 _19515_ (.A1(_06146_),
    .A2(_09763_),
    .B1(_03307_),
    .Y(_00951_));
 sky130_fd_sc_hd__or2_1 _19516_ (.A(_09744_),
    .B(_09752_),
    .X(_03308_));
 sky130_fd_sc_hd__xnor2_1 _19517_ (.A(_09751_),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__mux2_1 _19518_ (.A0(\rbzero.debug_overlay.playerX[3] ),
    .A1(_03309_),
    .S(_09784_),
    .X(_03310_));
 sky130_fd_sc_hd__mux2_1 _19519_ (.A0(_06105_),
    .A1(_03310_),
    .S(_09826_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_1 _19520_ (.A(_03311_),
    .X(_00952_));
 sky130_fd_sc_hd__nor2_1 _19521_ (.A(_09743_),
    .B(_09753_),
    .Y(_03312_));
 sky130_fd_sc_hd__and2_1 _19522_ (.A(_09743_),
    .B(_09753_),
    .X(_03313_));
 sky130_fd_sc_hd__or2_1 _19523_ (.A(_06101_),
    .B(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__a2bb2o_1 _19524_ (.A1_N(_03312_),
    .A2_N(_03314_),
    .B1(\rbzero.debug_overlay.playerX[4] ),
    .B2(_09824_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _19525_ (.A0(\rbzero.map_rom.i_col[4] ),
    .A1(_03315_),
    .S(_09826_),
    .X(_03316_));
 sky130_fd_sc_hd__clkbuf_1 _19526_ (.A(_03316_),
    .X(_00953_));
 sky130_fd_sc_hd__a21oi_1 _19527_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(_09100_),
    .B1(_03313_),
    .Y(_03317_));
 sky130_fd_sc_hd__nor2_1 _19528_ (.A(_09742_),
    .B(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__a21o_1 _19529_ (.A1(_09742_),
    .A2(_03317_),
    .B1(_06102_),
    .X(_03319_));
 sky130_fd_sc_hd__o22a_1 _19530_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_08100_),
    .B1(_03318_),
    .B2(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _19531_ (.A0(\rbzero.wall_tracer.mapX[5] ),
    .A1(_03320_),
    .S(_09782_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_1 _19532_ (.A(_03321_),
    .X(_00954_));
 sky130_fd_sc_hd__nor2_2 _19533_ (.A(net41),
    .B(net40),
    .Y(_03322_));
 sky130_fd_sc_hd__and3_1 _19534_ (.A(\rbzero.pov.ready ),
    .B(_02681_),
    .C(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__a21o_2 _19535_ (.A1(net40),
    .A2(_02682_),
    .B1(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_4 _19536_ (.A(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__inv_2 _19537_ (.A(\rbzero.pov.ready_buffer[59] ),
    .Y(_03326_));
 sky130_fd_sc_hd__nor2_1 _19538_ (.A(_02685_),
    .B(_03322_),
    .Y(_03327_));
 sky130_fd_sc_hd__buf_4 _19539_ (.A(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_1 _19540_ (.A0(_03326_),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__nand2_1 _19541_ (.A(_03329_),
    .B(_03325_),
    .Y(_03330_));
 sky130_fd_sc_hd__o211a_1 _19542_ (.A1(\rbzero.debug_overlay.playerX[-9] ),
    .A2(_03325_),
    .B1(_03330_),
    .C1(_03096_),
    .X(_00955_));
 sky130_fd_sc_hd__a21oi_1 _19543_ (.A1(net40),
    .A2(_02682_),
    .B1(_03323_),
    .Y(_03331_));
 sky130_fd_sc_hd__buf_2 _19544_ (.A(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _19545_ (.A0(\rbzero.pov.ready_buffer[60] ),
    .A1(_08167_),
    .S(_03328_),
    .X(_03333_));
 sky130_fd_sc_hd__or2_1 _19546_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(_03324_),
    .X(_03334_));
 sky130_fd_sc_hd__o211a_1 _19547_ (.A1(_03332_),
    .A2(_03333_),
    .B1(_03334_),
    .C1(_03096_),
    .X(_00956_));
 sky130_fd_sc_hd__clkbuf_4 _19548_ (.A(_03327_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _19549_ (.A0(\rbzero.pov.ready_buffer[61] ),
    .A1(_08181_),
    .S(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__or2_1 _19550_ (.A(_03332_),
    .B(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__o211a_1 _19551_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_03325_),
    .B1(_03337_),
    .C1(_03096_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _19552_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(_08201_),
    .S(_03335_),
    .X(_03338_));
 sky130_fd_sc_hd__or2_1 _19553_ (.A(_03332_),
    .B(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__o211a_1 _19554_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_03325_),
    .B1(_03339_),
    .C1(_03096_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _19555_ (.A0(\rbzero.pov.ready_buffer[63] ),
    .A1(_08219_),
    .S(_03335_),
    .X(_03340_));
 sky130_fd_sc_hd__or2_1 _19556_ (.A(_03332_),
    .B(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__o211a_1 _19557_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_03325_),
    .B1(_03341_),
    .C1(_03096_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _19558_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(_08239_),
    .S(_03335_),
    .X(_03342_));
 sky130_fd_sc_hd__or2_1 _19559_ (.A(_03331_),
    .B(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__o211a_1 _19560_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_03325_),
    .B1(_03343_),
    .C1(_03096_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _19561_ (.A0(\rbzero.pov.ready_buffer[65] ),
    .A1(_08264_),
    .S(_03335_),
    .X(_03344_));
 sky130_fd_sc_hd__or2_1 _19562_ (.A(_03331_),
    .B(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__clkbuf_4 _19563_ (.A(_02997_),
    .X(_03346_));
 sky130_fd_sc_hd__o211a_1 _19564_ (.A1(\rbzero.debug_overlay.playerX[-3] ),
    .A2(_03325_),
    .B1(_03345_),
    .C1(_03346_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _19565_ (.A0(\rbzero.pov.ready_buffer[66] ),
    .A1(_08293_),
    .S(_03335_),
    .X(_03347_));
 sky130_fd_sc_hd__or2_1 _19566_ (.A(_03331_),
    .B(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__o211a_1 _19567_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_03325_),
    .B1(_03348_),
    .C1(_03346_),
    .X(_00962_));
 sky130_fd_sc_hd__clkbuf_4 _19568_ (.A(_03335_),
    .X(_03349_));
 sky130_fd_sc_hd__or2_1 _19569_ (.A(_02685_),
    .B(_03322_),
    .X(_03350_));
 sky130_fd_sc_hd__or2_1 _19570_ (.A(_08305_),
    .B(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__o211a_1 _19571_ (.A1(\rbzero.pov.ready_buffer[67] ),
    .A2(_03349_),
    .B1(_03324_),
    .C1(_03351_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_4 _19572_ (.A(_04450_),
    .X(_03353_));
 sky130_fd_sc_hd__a211o_1 _19573_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_03332_),
    .B1(_03352_),
    .C1(_03353_),
    .X(_00963_));
 sky130_fd_sc_hd__and2_1 _19574_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_08303_),
    .X(_03354_));
 sky130_fd_sc_hd__or2_1 _19575_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_08303_),
    .X(_03355_));
 sky130_fd_sc_hd__or3b_1 _19576_ (.A(_03354_),
    .B(_03350_),
    .C_N(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__o211a_1 _19577_ (.A1(\rbzero.pov.ready_buffer[68] ),
    .A2(_03349_),
    .B1(_03324_),
    .C1(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__a211o_1 _19578_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03332_),
    .B1(_03357_),
    .C1(_03353_),
    .X(_00964_));
 sky130_fd_sc_hd__clkbuf_4 _19579_ (.A(_03350_),
    .X(_03358_));
 sky130_fd_sc_hd__nor2_1 _19580_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03355_),
    .Y(_03359_));
 sky130_fd_sc_hd__and2_1 _19581_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03355_),
    .X(_03360_));
 sky130_fd_sc_hd__or2_1 _19582_ (.A(\rbzero.pov.ready_buffer[69] ),
    .B(_03335_),
    .X(_03361_));
 sky130_fd_sc_hd__o311a_1 _19583_ (.A1(_03358_),
    .A2(_03359_),
    .A3(_03360_),
    .B1(_03324_),
    .C1(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__a211o_1 _19584_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03332_),
    .B1(_03362_),
    .C1(_03353_),
    .X(_00965_));
 sky130_fd_sc_hd__or3_1 _19585_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .B(\rbzero.debug_overlay.playerX[1] ),
    .C(_03355_),
    .X(_03363_));
 sky130_fd_sc_hd__o21ai_1 _19586_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03355_),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .Y(_03364_));
 sky130_fd_sc_hd__a21oi_1 _19587_ (.A1(_03363_),
    .A2(_03364_),
    .B1(_03358_),
    .Y(_03365_));
 sky130_fd_sc_hd__a211o_1 _19588_ (.A1(\rbzero.pov.ready_buffer[70] ),
    .A2(_03358_),
    .B1(_03332_),
    .C1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__o211a_1 _19589_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_03325_),
    .B1(_03366_),
    .C1(_03346_),
    .X(_00966_));
 sky130_fd_sc_hd__inv_2 _19590_ (.A(net40),
    .Y(_03367_));
 sky130_fd_sc_hd__nand2_1 _19591_ (.A(\rbzero.pov.ready ),
    .B(_03322_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _19592_ (.A(_05711_),
    .B(_04675_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand3_1 _19593_ (.A(_05770_),
    .B(_05769_),
    .C(_09709_),
    .Y(_03370_));
 sky130_fd_sc_hd__or2_1 _19594_ (.A(_03369_),
    .B(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__a211o_1 _19595_ (.A1(_03367_),
    .A2(_03368_),
    .B1(_03371_),
    .C1(_02678_),
    .X(_03372_));
 sky130_fd_sc_hd__or2_1 _19596_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_03363_),
    .X(_03373_));
 sky130_fd_sc_hd__and2b_1 _19597_ (.A_N(_03322_),
    .B(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__a2bb2o_1 _19598_ (.A1_N(_03372_),
    .A2_N(_03374_),
    .B1(_03363_),
    .B2(\rbzero.debug_overlay.playerX[3] ),
    .X(_03375_));
 sky130_fd_sc_hd__o21a_1 _19599_ (.A1(\rbzero.pov.ready_buffer[71] ),
    .A2(_03349_),
    .B1(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__a211o_1 _19600_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03332_),
    .B1(_03376_),
    .C1(_03353_),
    .X(_00967_));
 sky130_fd_sc_hd__o21a_1 _19601_ (.A1(_03332_),
    .A2(_03374_),
    .B1(\rbzero.debug_overlay.playerX[4] ),
    .X(_03377_));
 sky130_fd_sc_hd__o21bai_1 _19602_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_03373_),
    .B1_N(_03322_),
    .Y(_03378_));
 sky130_fd_sc_hd__o211a_1 _19603_ (.A1(\rbzero.pov.ready_buffer[72] ),
    .A2(_03349_),
    .B1(_03325_),
    .C1(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__o21a_1 _19604_ (.A1(_03377_),
    .A2(_03379_),
    .B1(_02639_),
    .X(_00968_));
 sky130_fd_sc_hd__a21bo_1 _19605_ (.A1(_03324_),
    .A2(_03378_),
    .B1_N(\rbzero.debug_overlay.playerX[5] ),
    .X(_03380_));
 sky130_fd_sc_hd__inv_2 _19606_ (.A(\rbzero.pov.ready_buffer[73] ),
    .Y(_03381_));
 sky130_fd_sc_hd__o31a_1 _19607_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(\rbzero.debug_overlay.playerX[4] ),
    .A3(_03373_),
    .B1(_03335_),
    .X(_03382_));
 sky130_fd_sc_hd__a211o_1 _19608_ (.A1(_03381_),
    .A2(_03358_),
    .B1(_03382_),
    .C1(_03372_),
    .X(_03383_));
 sky130_fd_sc_hd__a21oi_1 _19609_ (.A1(_03380_),
    .A2(_03383_),
    .B1(_03353_),
    .Y(_00969_));
 sky130_fd_sc_hd__clkbuf_4 _19610_ (.A(_03323_),
    .X(_03384_));
 sky130_fd_sc_hd__a21oi_4 _19611_ (.A1(net41),
    .A2(_02682_),
    .B1(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__clkbuf_4 _19612_ (.A(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _19613_ (.A0(\rbzero.pov.ready_buffer[44] ),
    .A1(_08417_),
    .S(_03328_),
    .X(_03387_));
 sky130_fd_sc_hd__nand2_1 _19614_ (.A(_08417_),
    .B(_03386_),
    .Y(_03388_));
 sky130_fd_sc_hd__o211a_1 _19615_ (.A1(_03386_),
    .A2(_03387_),
    .B1(_03388_),
    .C1(_03346_),
    .X(_00970_));
 sky130_fd_sc_hd__a21o_1 _19616_ (.A1(net41),
    .A2(_02682_),
    .B1(_03323_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_4 _19617_ (.A(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__nand2_1 _19618_ (.A(\rbzero.pov.ready_buffer[45] ),
    .B(_03358_),
    .Y(_03391_));
 sky130_fd_sc_hd__o211ai_1 _19619_ (.A1(_08157_),
    .A2(_03358_),
    .B1(_03390_),
    .C1(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__o211a_1 _19620_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(_03390_),
    .B1(_03392_),
    .C1(_03346_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _19621_ (.A0(\rbzero.pov.ready_buffer[46] ),
    .A1(_08186_),
    .S(_03328_),
    .X(_03393_));
 sky130_fd_sc_hd__or2_1 _19622_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(_03390_),
    .X(_03394_));
 sky130_fd_sc_hd__o211a_1 _19623_ (.A1(_03386_),
    .A2(_03393_),
    .B1(_03394_),
    .C1(_03346_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _19624_ (.A0(\rbzero.pov.ready_buffer[47] ),
    .A1(_08195_),
    .S(_03328_),
    .X(_03395_));
 sky130_fd_sc_hd__or2_1 _19625_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_03390_),
    .X(_03396_));
 sky130_fd_sc_hd__o211a_1 _19626_ (.A1(_03386_),
    .A2(_03395_),
    .B1(_03396_),
    .C1(_03346_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _19627_ (.A0(\rbzero.pov.ready_buffer[48] ),
    .A1(_08215_),
    .S(_03328_),
    .X(_03397_));
 sky130_fd_sc_hd__or2_1 _19628_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_03389_),
    .X(_03398_));
 sky130_fd_sc_hd__o211a_1 _19629_ (.A1(_03386_),
    .A2(_03397_),
    .B1(_03398_),
    .C1(_03346_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _19630_ (.A0(\rbzero.pov.ready_buffer[49] ),
    .A1(_08233_),
    .S(_03328_),
    .X(_03399_));
 sky130_fd_sc_hd__or2_1 _19631_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(_03389_),
    .X(_03400_));
 sky130_fd_sc_hd__o211a_1 _19632_ (.A1(_03386_),
    .A2(_03399_),
    .B1(_03400_),
    .C1(_03346_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _19633_ (.A0(\rbzero.pov.ready_buffer[50] ),
    .A1(_08258_),
    .S(_03328_),
    .X(_03401_));
 sky130_fd_sc_hd__nand2_1 _19634_ (.A(_05056_),
    .B(_03385_),
    .Y(_03402_));
 sky130_fd_sc_hd__o211a_1 _19635_ (.A1(_03386_),
    .A2(_03401_),
    .B1(_03402_),
    .C1(_03346_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _19636_ (.A0(\rbzero.pov.ready_buffer[51] ),
    .A1(_08289_),
    .S(_03328_),
    .X(_03403_));
 sky130_fd_sc_hd__or2_1 _19637_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_03389_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_4 _19638_ (.A(_02997_),
    .X(_03405_));
 sky130_fd_sc_hd__o211a_1 _19639_ (.A1(_03386_),
    .A2(_03403_),
    .B1(_03404_),
    .C1(_03405_),
    .X(_00977_));
 sky130_fd_sc_hd__a21oi_1 _19640_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_03385_),
    .B1(_02731_),
    .Y(_03406_));
 sky130_fd_sc_hd__nor2_1 _19641_ (.A(\rbzero.pov.ready_buffer[52] ),
    .B(_03349_),
    .Y(_03407_));
 sky130_fd_sc_hd__a211o_1 _19642_ (.A1(_08300_),
    .A2(_03349_),
    .B1(_03385_),
    .C1(_03407_),
    .X(_03408_));
 sky130_fd_sc_hd__nand2_1 _19643_ (.A(_03406_),
    .B(_03408_),
    .Y(_00978_));
 sky130_fd_sc_hd__or2_1 _19644_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08298_),
    .X(_03409_));
 sky130_fd_sc_hd__nand2_1 _19645_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08298_),
    .Y(_03410_));
 sky130_fd_sc_hd__a21oi_1 _19646_ (.A1(_03409_),
    .A2(_03410_),
    .B1(_03358_),
    .Y(_03411_));
 sky130_fd_sc_hd__a211o_1 _19647_ (.A1(\rbzero.pov.ready_buffer[53] ),
    .A2(_03358_),
    .B1(_03385_),
    .C1(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__o211a_1 _19648_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_03390_),
    .B1(_03412_),
    .C1(_03405_),
    .X(_00979_));
 sky130_fd_sc_hd__and2_1 _19649_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(_03409_),
    .X(_03413_));
 sky130_fd_sc_hd__nor2_1 _19650_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(_03409_),
    .Y(_03414_));
 sky130_fd_sc_hd__or2_1 _19651_ (.A(_03350_),
    .B(_03414_),
    .X(_03415_));
 sky130_fd_sc_hd__o221a_1 _19652_ (.A1(\rbzero.pov.ready_buffer[54] ),
    .A2(_03349_),
    .B1(_03413_),
    .B2(_03415_),
    .C1(_03390_),
    .X(_03416_));
 sky130_fd_sc_hd__a211o_1 _19653_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03386_),
    .B1(_03416_),
    .C1(_03353_),
    .X(_00980_));
 sky130_fd_sc_hd__a21o_1 _19654_ (.A1(_03390_),
    .A2(_03415_),
    .B1(_06127_),
    .X(_03417_));
 sky130_fd_sc_hd__nand2_1 _19655_ (.A(_06127_),
    .B(_03414_),
    .Y(_03418_));
 sky130_fd_sc_hd__nor2_1 _19656_ (.A(\rbzero.pov.ready_buffer[55] ),
    .B(_03328_),
    .Y(_03419_));
 sky130_fd_sc_hd__a211o_1 _19657_ (.A1(_03349_),
    .A2(_03418_),
    .B1(_03419_),
    .C1(_03385_),
    .X(_03420_));
 sky130_fd_sc_hd__a21oi_1 _19658_ (.A1(_03417_),
    .A2(_03420_),
    .B1(_03353_),
    .Y(_00981_));
 sky130_fd_sc_hd__or2_1 _19659_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .B(_03418_),
    .X(_03421_));
 sky130_fd_sc_hd__and2b_1 _19660_ (.A_N(_03322_),
    .B(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__inv_2 _19661_ (.A(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21o_1 _19662_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03418_),
    .B1(_02732_),
    .X(_03424_));
 sky130_fd_sc_hd__o221a_1 _19663_ (.A1(\rbzero.pov.ready_buffer[56] ),
    .A2(_03349_),
    .B1(_03423_),
    .B2(_03424_),
    .C1(_03390_),
    .X(_03425_));
 sky130_fd_sc_hd__a211o_1 _19664_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03386_),
    .B1(_03425_),
    .C1(_03353_),
    .X(_00982_));
 sky130_fd_sc_hd__o21a_1 _19665_ (.A1(_03385_),
    .A2(_03422_),
    .B1(\rbzero.debug_overlay.playerY[4] ),
    .X(_03426_));
 sky130_fd_sc_hd__a41o_1 _19666_ (.A1(_04997_),
    .A2(_04993_),
    .A3(_06127_),
    .A4(_03414_),
    .B1(_03322_),
    .X(_03427_));
 sky130_fd_sc_hd__o211a_1 _19667_ (.A1(\rbzero.pov.ready_buffer[57] ),
    .A2(_03349_),
    .B1(_03390_),
    .C1(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__o21a_1 _19668_ (.A1(_03426_),
    .A2(_03428_),
    .B1(_02639_),
    .X(_00983_));
 sky130_fd_sc_hd__a21o_1 _19669_ (.A1(_03390_),
    .A2(_03427_),
    .B1(_06123_),
    .X(_03429_));
 sky130_fd_sc_hd__inv_2 _19670_ (.A(\rbzero.pov.ready_buffer[58] ),
    .Y(_03430_));
 sky130_fd_sc_hd__o31a_1 _19671_ (.A1(\rbzero.debug_overlay.playerY[5] ),
    .A2(\rbzero.debug_overlay.playerY[4] ),
    .A3(_03421_),
    .B1(_03335_),
    .X(_03431_));
 sky130_fd_sc_hd__a211o_1 _19672_ (.A1(_03430_),
    .A2(_03358_),
    .B1(_03385_),
    .C1(_03431_),
    .X(_03432_));
 sky130_fd_sc_hd__a21oi_1 _19673_ (.A1(_03429_),
    .A2(_03432_),
    .B1(_03353_),
    .Y(_00984_));
 sky130_fd_sc_hd__clkbuf_2 _19674_ (.A(_03384_),
    .X(_03433_));
 sky130_fd_sc_hd__or2b_1 _19675_ (.A(\rbzero.pov.ready_buffer[33] ),
    .B_N(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__o211a_1 _19676_ (.A1(\rbzero.debug_overlay.facingX[-9] ),
    .A2(_03433_),
    .B1(_03434_),
    .C1(_03405_),
    .X(_00985_));
 sky130_fd_sc_hd__or3b_1 _19677_ (.A(_03327_),
    .B(_02685_),
    .C_N(\rbzero.pov.ready ),
    .X(_03435_));
 sky130_fd_sc_hd__buf_2 _19678_ (.A(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__buf_2 _19679_ (.A(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__or2_1 _19680_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(_03433_),
    .X(_03438_));
 sky130_fd_sc_hd__o211a_1 _19681_ (.A1(\rbzero.pov.ready_buffer[34] ),
    .A2(_03437_),
    .B1(_03438_),
    .C1(_03405_),
    .X(_00986_));
 sky130_fd_sc_hd__or2_1 _19682_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(_03433_),
    .X(_03439_));
 sky130_fd_sc_hd__o211a_1 _19683_ (.A1(\rbzero.pov.ready_buffer[35] ),
    .A2(_03437_),
    .B1(_03439_),
    .C1(_03405_),
    .X(_00987_));
 sky130_fd_sc_hd__or2_1 _19684_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(_03433_),
    .X(_03440_));
 sky130_fd_sc_hd__o211a_1 _19685_ (.A1(\rbzero.pov.ready_buffer[36] ),
    .A2(_03437_),
    .B1(_03440_),
    .C1(_03405_),
    .X(_00988_));
 sky130_fd_sc_hd__buf_2 _19686_ (.A(_03436_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_2 _19687_ (.A(_03384_),
    .X(_03442_));
 sky130_fd_sc_hd__and2_1 _19688_ (.A(\rbzero.pov.ready_buffer[37] ),
    .B(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__buf_2 _19689_ (.A(_04450_),
    .X(_03444_));
 sky130_fd_sc_hd__a211o_1 _19690_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_03441_),
    .B1(_03443_),
    .C1(_03444_),
    .X(_00989_));
 sky130_fd_sc_hd__and2_1 _19691_ (.A(\rbzero.pov.ready_buffer[38] ),
    .B(_03442_),
    .X(_03445_));
 sky130_fd_sc_hd__a211o_1 _19692_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_03441_),
    .B1(_03445_),
    .C1(_03444_),
    .X(_00990_));
 sky130_fd_sc_hd__and2_1 _19693_ (.A(\rbzero.pov.ready_buffer[39] ),
    .B(_03442_),
    .X(_03446_));
 sky130_fd_sc_hd__a211o_1 _19694_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_03441_),
    .B1(_03446_),
    .C1(_03444_),
    .X(_00991_));
 sky130_fd_sc_hd__or2_1 _19695_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(_03433_),
    .X(_03447_));
 sky130_fd_sc_hd__o211a_1 _19696_ (.A1(net514),
    .A2(_03437_),
    .B1(_03447_),
    .C1(_03405_),
    .X(_00992_));
 sky130_fd_sc_hd__and2_1 _19697_ (.A(\rbzero.pov.ready_buffer[41] ),
    .B(_03442_),
    .X(_03448_));
 sky130_fd_sc_hd__a211o_1 _19698_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(_03441_),
    .B1(_03448_),
    .C1(_03444_),
    .X(_00993_));
 sky130_fd_sc_hd__or2_1 _19699_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(_03433_),
    .X(_03449_));
 sky130_fd_sc_hd__o211a_1 _19700_ (.A1(\rbzero.pov.ready_buffer[42] ),
    .A2(_03437_),
    .B1(_03449_),
    .C1(_03405_),
    .X(_00994_));
 sky130_fd_sc_hd__or2_1 _19701_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(_03433_),
    .X(_03450_));
 sky130_fd_sc_hd__o211a_1 _19702_ (.A1(\rbzero.pov.ready_buffer[43] ),
    .A2(_03437_),
    .B1(_03450_),
    .C1(_03405_),
    .X(_00995_));
 sky130_fd_sc_hd__clkbuf_2 _19703_ (.A(_03384_),
    .X(_03451_));
 sky130_fd_sc_hd__and2_1 _19704_ (.A(\rbzero.pov.ready_buffer[22] ),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__a211o_1 _19705_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(_03441_),
    .B1(_03452_),
    .C1(_03444_),
    .X(_00996_));
 sky130_fd_sc_hd__or2_1 _19706_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_03433_),
    .X(_03453_));
 sky130_fd_sc_hd__o211a_1 _19707_ (.A1(\rbzero.pov.ready_buffer[23] ),
    .A2(_03437_),
    .B1(_03453_),
    .C1(_03405_),
    .X(_00997_));
 sky130_fd_sc_hd__and2_1 _19708_ (.A(\rbzero.pov.ready_buffer[24] ),
    .B(_03451_),
    .X(_03454_));
 sky130_fd_sc_hd__a211o_1 _19709_ (.A1(\rbzero.debug_overlay.facingY[-7] ),
    .A2(_03441_),
    .B1(_03454_),
    .C1(_03444_),
    .X(_00998_));
 sky130_fd_sc_hd__clkbuf_4 _19710_ (.A(_03436_),
    .X(_03455_));
 sky130_fd_sc_hd__and2_1 _19711_ (.A(\rbzero.pov.ready_buffer[25] ),
    .B(_03451_),
    .X(_03456_));
 sky130_fd_sc_hd__a211o_1 _19712_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03444_),
    .X(_00999_));
 sky130_fd_sc_hd__and2_1 _19713_ (.A(\rbzero.pov.ready_buffer[26] ),
    .B(_03451_),
    .X(_03457_));
 sky130_fd_sc_hd__a211o_1 _19714_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_03455_),
    .B1(_03457_),
    .C1(_03444_),
    .X(_01000_));
 sky130_fd_sc_hd__or2_1 _19715_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(_03433_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_4 _19716_ (.A(_02638_),
    .X(_03459_));
 sky130_fd_sc_hd__o211a_1 _19717_ (.A1(\rbzero.pov.ready_buffer[27] ),
    .A2(_03437_),
    .B1(_03458_),
    .C1(_03459_),
    .X(_01001_));
 sky130_fd_sc_hd__clkbuf_2 _19718_ (.A(_03384_),
    .X(_03460_));
 sky130_fd_sc_hd__or2_1 _19719_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__o211a_1 _19720_ (.A1(\rbzero.pov.ready_buffer[28] ),
    .A2(_03437_),
    .B1(_03461_),
    .C1(_03459_),
    .X(_01002_));
 sky130_fd_sc_hd__and2_1 _19721_ (.A(\rbzero.pov.ready_buffer[29] ),
    .B(_03451_),
    .X(_03462_));
 sky130_fd_sc_hd__a211o_1 _19722_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(_03455_),
    .B1(_03462_),
    .C1(_03444_),
    .X(_01003_));
 sky130_fd_sc_hd__or2_1 _19723_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(_03460_),
    .X(_03463_));
 sky130_fd_sc_hd__o211a_1 _19724_ (.A1(\rbzero.pov.ready_buffer[30] ),
    .A2(_03437_),
    .B1(_03463_),
    .C1(_03459_),
    .X(_01004_));
 sky130_fd_sc_hd__and2_1 _19725_ (.A(\rbzero.pov.ready_buffer[31] ),
    .B(_03451_),
    .X(_03464_));
 sky130_fd_sc_hd__a211o_1 _19726_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_03455_),
    .B1(_03464_),
    .C1(_03444_),
    .X(_01005_));
 sky130_fd_sc_hd__and2_1 _19727_ (.A(\rbzero.pov.ready_buffer[32] ),
    .B(_03451_),
    .X(_03465_));
 sky130_fd_sc_hd__buf_4 _19728_ (.A(_04450_),
    .X(_03466_));
 sky130_fd_sc_hd__a211o_1 _19729_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_03455_),
    .B1(_03465_),
    .C1(_03466_),
    .X(_01006_));
 sky130_fd_sc_hd__and2_1 _19730_ (.A(\rbzero.pov.ready_buffer[11] ),
    .B(_03451_),
    .X(_03467_));
 sky130_fd_sc_hd__a211o_1 _19731_ (.A1(_05290_),
    .A2(_03455_),
    .B1(_03467_),
    .C1(_03466_),
    .X(_01007_));
 sky130_fd_sc_hd__buf_2 _19732_ (.A(_03436_),
    .X(_03468_));
 sky130_fd_sc_hd__or2_1 _19733_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(_03460_),
    .X(_03469_));
 sky130_fd_sc_hd__o211a_1 _19734_ (.A1(\rbzero.pov.ready_buffer[12] ),
    .A2(_03468_),
    .B1(_03469_),
    .C1(_03459_),
    .X(_01008_));
 sky130_fd_sc_hd__or2_1 _19735_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_03460_),
    .X(_03470_));
 sky130_fd_sc_hd__o211a_1 _19736_ (.A1(\rbzero.pov.ready_buffer[13] ),
    .A2(_03468_),
    .B1(_03470_),
    .C1(_03459_),
    .X(_01009_));
 sky130_fd_sc_hd__or2_1 _19737_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .B(_03460_),
    .X(_03471_));
 sky130_fd_sc_hd__o211a_1 _19738_ (.A1(\rbzero.pov.ready_buffer[14] ),
    .A2(_03468_),
    .B1(_03471_),
    .C1(_03459_),
    .X(_01010_));
 sky130_fd_sc_hd__and2_1 _19739_ (.A(\rbzero.pov.ready_buffer[15] ),
    .B(_03451_),
    .X(_03472_));
 sky130_fd_sc_hd__a211o_1 _19740_ (.A1(_05291_),
    .A2(_03455_),
    .B1(_03472_),
    .C1(_03466_),
    .X(_01011_));
 sky130_fd_sc_hd__and2_1 _19741_ (.A(\rbzero.pov.ready_buffer[16] ),
    .B(_03451_),
    .X(_03473_));
 sky130_fd_sc_hd__a211o_1 _19742_ (.A1(_05292_),
    .A2(_03455_),
    .B1(_03473_),
    .C1(_03466_),
    .X(_01012_));
 sky130_fd_sc_hd__or2_1 _19743_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(_03460_),
    .X(_03474_));
 sky130_fd_sc_hd__o211a_1 _19744_ (.A1(\rbzero.pov.ready_buffer[17] ),
    .A2(_03468_),
    .B1(_03474_),
    .C1(_03459_),
    .X(_01013_));
 sky130_fd_sc_hd__and2_1 _19745_ (.A(\rbzero.pov.ready_buffer[18] ),
    .B(_03384_),
    .X(_03475_));
 sky130_fd_sc_hd__a211o_1 _19746_ (.A1(_02443_),
    .A2(_03455_),
    .B1(_03475_),
    .C1(_03466_),
    .X(_01014_));
 sky130_fd_sc_hd__or2_1 _19747_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_03460_),
    .X(_03476_));
 sky130_fd_sc_hd__o211a_1 _19748_ (.A1(\rbzero.pov.ready_buffer[19] ),
    .A2(_03468_),
    .B1(_03476_),
    .C1(_03459_),
    .X(_01015_));
 sky130_fd_sc_hd__or2_1 _19749_ (.A(_02465_),
    .B(_03460_),
    .X(_03477_));
 sky130_fd_sc_hd__o211a_1 _19750_ (.A1(\rbzero.pov.ready_buffer[20] ),
    .A2(_03468_),
    .B1(_03477_),
    .C1(_03459_),
    .X(_01016_));
 sky130_fd_sc_hd__or2_1 _19751_ (.A(_02495_),
    .B(_03460_),
    .X(_03478_));
 sky130_fd_sc_hd__o211a_1 _19752_ (.A1(\rbzero.pov.ready_buffer[21] ),
    .A2(_03468_),
    .B1(_03478_),
    .C1(_03459_),
    .X(_01017_));
 sky130_fd_sc_hd__or2_1 _19753_ (.A(_05282_),
    .B(_03460_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_4 _19754_ (.A(_02638_),
    .X(_03480_));
 sky130_fd_sc_hd__o211a_1 _19755_ (.A1(\rbzero.pov.ready_buffer[0] ),
    .A2(_03468_),
    .B1(_03479_),
    .C1(_03480_),
    .X(_01018_));
 sky130_fd_sc_hd__or2_1 _19756_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_03442_),
    .X(_03481_));
 sky130_fd_sc_hd__o211a_1 _19757_ (.A1(\rbzero.pov.ready_buffer[1] ),
    .A2(_03468_),
    .B1(_03481_),
    .C1(_03480_),
    .X(_01019_));
 sky130_fd_sc_hd__or2_1 _19758_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03442_),
    .X(_03482_));
 sky130_fd_sc_hd__o211a_1 _19759_ (.A1(\rbzero.pov.ready_buffer[2] ),
    .A2(_03468_),
    .B1(_03482_),
    .C1(_03480_),
    .X(_01020_));
 sky130_fd_sc_hd__and2_1 _19760_ (.A(\rbzero.pov.ready_buffer[3] ),
    .B(_03384_),
    .X(_03483_));
 sky130_fd_sc_hd__a211o_1 _19761_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(_03455_),
    .B1(_03483_),
    .C1(_03466_),
    .X(_01021_));
 sky130_fd_sc_hd__and2_1 _19762_ (.A(\rbzero.pov.ready_buffer[4] ),
    .B(_03384_),
    .X(_03484_));
 sky130_fd_sc_hd__a211o_1 _19763_ (.A1(_03111_),
    .A2(_03436_),
    .B1(_03484_),
    .C1(_03466_),
    .X(_01022_));
 sky130_fd_sc_hd__and2_1 _19764_ (.A(\rbzero.pov.ready_buffer[5] ),
    .B(_03384_),
    .X(_03485_));
 sky130_fd_sc_hd__a211o_1 _19765_ (.A1(_03127_),
    .A2(_03436_),
    .B1(_03485_),
    .C1(_03466_),
    .X(_01023_));
 sky130_fd_sc_hd__or2_1 _19766_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(_03442_),
    .X(_03486_));
 sky130_fd_sc_hd__o211a_1 _19767_ (.A1(\rbzero.pov.ready_buffer[6] ),
    .A2(_03441_),
    .B1(_03486_),
    .C1(_03480_),
    .X(_01024_));
 sky130_fd_sc_hd__and2_1 _19768_ (.A(\rbzero.pov.ready_buffer[7] ),
    .B(_03384_),
    .X(_03487_));
 sky130_fd_sc_hd__a211o_1 _19769_ (.A1(\rbzero.debug_overlay.vplaneY[-2] ),
    .A2(_03436_),
    .B1(_03487_),
    .C1(_03466_),
    .X(_01025_));
 sky130_fd_sc_hd__or2_1 _19770_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_03442_),
    .X(_03488_));
 sky130_fd_sc_hd__o211a_1 _19771_ (.A1(\rbzero.pov.ready_buffer[8] ),
    .A2(_03441_),
    .B1(_03488_),
    .C1(_03480_),
    .X(_01026_));
 sky130_fd_sc_hd__or2_1 _19772_ (.A(_03167_),
    .B(_03442_),
    .X(_03489_));
 sky130_fd_sc_hd__o211a_1 _19773_ (.A1(\rbzero.pov.ready_buffer[9] ),
    .A2(_03441_),
    .B1(_03489_),
    .C1(_03480_),
    .X(_01027_));
 sky130_fd_sc_hd__or2_1 _19774_ (.A(_03196_),
    .B(_03442_),
    .X(_03490_));
 sky130_fd_sc_hd__o211a_1 _19775_ (.A1(\rbzero.pov.ready_buffer[10] ),
    .A2(_03441_),
    .B1(_03490_),
    .C1(_03480_),
    .X(_01028_));
 sky130_fd_sc_hd__and2b_1 _19776_ (.A_N(\rbzero.pov.sclk_buffer[2] ),
    .B(\rbzero.pov.sclk_buffer[1] ),
    .X(_03491_));
 sky130_fd_sc_hd__and2_1 _19777_ (.A(\rbzero.pov.spi_counter[0] ),
    .B(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__nor2_2 _19778_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(_04094_),
    .Y(_03493_));
 sky130_fd_sc_hd__o21ai_1 _19779_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03491_),
    .B1(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__nor2_1 _19780_ (.A(_03492_),
    .B(_03494_),
    .Y(_01029_));
 sky130_fd_sc_hd__and3_1 _19781_ (.A(\rbzero.pov.spi_counter[1] ),
    .B(\rbzero.pov.spi_counter[0] ),
    .C(_03491_),
    .X(_03495_));
 sky130_fd_sc_hd__clkinv_2 _19782_ (.A(\rbzero.pov.spi_counter[6] ),
    .Y(_03496_));
 sky130_fd_sc_hd__or4b_1 _19783_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[2] ),
    .C(\rbzero.pov.spi_counter[1] ),
    .D_N(\rbzero.pov.spi_counter[3] ),
    .X(_03497_));
 sky130_fd_sc_hd__or4b_1 _19784_ (.A(_03496_),
    .B(_03497_),
    .C(\rbzero.pov.spi_counter[5] ),
    .D_N(_03492_),
    .X(_03498_));
 sky130_fd_sc_hd__and2_1 _19785_ (.A(_03493_),
    .B(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__o21ai_1 _19786_ (.A1(\rbzero.pov.spi_counter[1] ),
    .A2(_03492_),
    .B1(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__nor2_1 _19787_ (.A(_03495_),
    .B(_03500_),
    .Y(_01030_));
 sky130_fd_sc_hd__and3_1 _19788_ (.A(\rbzero.pov.spi_counter[2] ),
    .B(\rbzero.pov.spi_counter[1] ),
    .C(_03492_),
    .X(_03501_));
 sky130_fd_sc_hd__o21ai_1 _19789_ (.A1(\rbzero.pov.spi_counter[2] ),
    .A2(_03495_),
    .B1(_03493_),
    .Y(_03502_));
 sky130_fd_sc_hd__nor2_1 _19790_ (.A(_03501_),
    .B(_03502_),
    .Y(_01031_));
 sky130_fd_sc_hd__and2_1 _19791_ (.A(\rbzero.pov.spi_counter[3] ),
    .B(_03501_),
    .X(_03503_));
 sky130_fd_sc_hd__o21ai_1 _19792_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_03501_),
    .B1(_03499_),
    .Y(_03504_));
 sky130_fd_sc_hd__nor2_1 _19793_ (.A(_03503_),
    .B(_03504_),
    .Y(_01032_));
 sky130_fd_sc_hd__and3_1 _19794_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[3] ),
    .C(_03501_),
    .X(_03505_));
 sky130_fd_sc_hd__o21ai_1 _19795_ (.A1(\rbzero.pov.spi_counter[4] ),
    .A2(_03503_),
    .B1(_03493_),
    .Y(_03506_));
 sky130_fd_sc_hd__nor2_1 _19796_ (.A(_03505_),
    .B(_03506_),
    .Y(_01033_));
 sky130_fd_sc_hd__and2_1 _19797_ (.A(\rbzero.pov.spi_counter[5] ),
    .B(_03505_),
    .X(_03507_));
 sky130_fd_sc_hd__o21ai_1 _19798_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_03505_),
    .B1(_03493_),
    .Y(_03508_));
 sky130_fd_sc_hd__nor2_1 _19799_ (.A(_03507_),
    .B(_03508_),
    .Y(_01034_));
 sky130_fd_sc_hd__a21boi_1 _19800_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03507_),
    .B1_N(_03499_),
    .Y(_03509_));
 sky130_fd_sc_hd__o21a_1 _19801_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03507_),
    .B1(_03509_),
    .X(_01035_));
 sky130_fd_sc_hd__and2b_1 _19802_ (.A_N(\rbzero.pov.ss_buffer[1] ),
    .B(_03491_),
    .X(_03510_));
 sky130_fd_sc_hd__buf_4 _19803_ (.A(_03510_),
    .X(_03511_));
 sky130_fd_sc_hd__buf_2 _19804_ (.A(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__or3b_1 _19805_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(\rbzero.pov.sclk_buffer[2] ),
    .C_N(\rbzero.pov.sclk_buffer[1] ),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_4 _19806_ (.A(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_2 _19807_ (.A(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__or2_1 _19808_ (.A(\rbzero.pov.mosi ),
    .B(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__o211a_1 _19809_ (.A1(\rbzero.pov.spi_buffer[0] ),
    .A2(_03512_),
    .B1(_03516_),
    .C1(_03480_),
    .X(_01036_));
 sky130_fd_sc_hd__or2_1 _19810_ (.A(\rbzero.pov.spi_buffer[0] ),
    .B(_03515_),
    .X(_03517_));
 sky130_fd_sc_hd__o211a_1 _19811_ (.A1(\rbzero.pov.spi_buffer[1] ),
    .A2(_03512_),
    .B1(_03517_),
    .C1(_03480_),
    .X(_01037_));
 sky130_fd_sc_hd__or2_1 _19812_ (.A(\rbzero.pov.spi_buffer[1] ),
    .B(_03515_),
    .X(_03518_));
 sky130_fd_sc_hd__o211a_1 _19813_ (.A1(\rbzero.pov.spi_buffer[2] ),
    .A2(_03512_),
    .B1(_03518_),
    .C1(_03480_),
    .X(_01038_));
 sky130_fd_sc_hd__or2_1 _19814_ (.A(\rbzero.pov.spi_buffer[2] ),
    .B(_03515_),
    .X(_03519_));
 sky130_fd_sc_hd__buf_2 _19815_ (.A(_02638_),
    .X(_03520_));
 sky130_fd_sc_hd__o211a_1 _19816_ (.A1(\rbzero.pov.spi_buffer[3] ),
    .A2(_03512_),
    .B1(_03519_),
    .C1(_03520_),
    .X(_01039_));
 sky130_fd_sc_hd__or2_1 _19817_ (.A(\rbzero.pov.spi_buffer[3] ),
    .B(_03515_),
    .X(_03521_));
 sky130_fd_sc_hd__o211a_1 _19818_ (.A1(\rbzero.pov.spi_buffer[4] ),
    .A2(_03512_),
    .B1(_03521_),
    .C1(_03520_),
    .X(_01040_));
 sky130_fd_sc_hd__or2_1 _19819_ (.A(\rbzero.pov.spi_buffer[4] ),
    .B(_03515_),
    .X(_03522_));
 sky130_fd_sc_hd__o211a_1 _19820_ (.A1(\rbzero.pov.spi_buffer[5] ),
    .A2(_03512_),
    .B1(_03522_),
    .C1(_03520_),
    .X(_01041_));
 sky130_fd_sc_hd__or2_1 _19821_ (.A(\rbzero.pov.spi_buffer[5] ),
    .B(_03515_),
    .X(_03523_));
 sky130_fd_sc_hd__o211a_1 _19822_ (.A1(\rbzero.pov.spi_buffer[6] ),
    .A2(_03512_),
    .B1(_03523_),
    .C1(_03520_),
    .X(_01042_));
 sky130_fd_sc_hd__or2_1 _19823_ (.A(\rbzero.pov.spi_buffer[6] ),
    .B(_03515_),
    .X(_03524_));
 sky130_fd_sc_hd__o211a_1 _19824_ (.A1(\rbzero.pov.spi_buffer[7] ),
    .A2(_03512_),
    .B1(_03524_),
    .C1(_03520_),
    .X(_01043_));
 sky130_fd_sc_hd__or2_1 _19825_ (.A(\rbzero.pov.spi_buffer[7] ),
    .B(_03515_),
    .X(_03525_));
 sky130_fd_sc_hd__o211a_1 _19826_ (.A1(\rbzero.pov.spi_buffer[8] ),
    .A2(_03512_),
    .B1(_03525_),
    .C1(_03520_),
    .X(_01044_));
 sky130_fd_sc_hd__or2_1 _19827_ (.A(\rbzero.pov.spi_buffer[8] ),
    .B(_03515_),
    .X(_03526_));
 sky130_fd_sc_hd__o211a_1 _19828_ (.A1(\rbzero.pov.spi_buffer[9] ),
    .A2(_03512_),
    .B1(_03526_),
    .C1(_03520_),
    .X(_01045_));
 sky130_fd_sc_hd__buf_2 _19829_ (.A(_03511_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_2 _19830_ (.A(_03514_),
    .X(_03528_));
 sky130_fd_sc_hd__or2_1 _19831_ (.A(\rbzero.pov.spi_buffer[9] ),
    .B(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__o211a_1 _19832_ (.A1(\rbzero.pov.spi_buffer[10] ),
    .A2(_03527_),
    .B1(_03529_),
    .C1(_03520_),
    .X(_01046_));
 sky130_fd_sc_hd__or2_1 _19833_ (.A(\rbzero.pov.spi_buffer[10] ),
    .B(_03528_),
    .X(_03530_));
 sky130_fd_sc_hd__o211a_1 _19834_ (.A1(\rbzero.pov.spi_buffer[11] ),
    .A2(_03527_),
    .B1(_03530_),
    .C1(_03520_),
    .X(_01047_));
 sky130_fd_sc_hd__or2_1 _19835_ (.A(\rbzero.pov.spi_buffer[11] ),
    .B(_03528_),
    .X(_03531_));
 sky130_fd_sc_hd__o211a_1 _19836_ (.A1(\rbzero.pov.spi_buffer[12] ),
    .A2(_03527_),
    .B1(_03531_),
    .C1(_03520_),
    .X(_01048_));
 sky130_fd_sc_hd__or2_1 _19837_ (.A(\rbzero.pov.spi_buffer[12] ),
    .B(_03528_),
    .X(_03532_));
 sky130_fd_sc_hd__buf_2 _19838_ (.A(_02638_),
    .X(_03533_));
 sky130_fd_sc_hd__o211a_1 _19839_ (.A1(\rbzero.pov.spi_buffer[13] ),
    .A2(_03527_),
    .B1(_03532_),
    .C1(_03533_),
    .X(_01049_));
 sky130_fd_sc_hd__or2_1 _19840_ (.A(\rbzero.pov.spi_buffer[13] ),
    .B(_03528_),
    .X(_03534_));
 sky130_fd_sc_hd__o211a_1 _19841_ (.A1(\rbzero.pov.spi_buffer[14] ),
    .A2(_03527_),
    .B1(_03534_),
    .C1(_03533_),
    .X(_01050_));
 sky130_fd_sc_hd__or2_1 _19842_ (.A(\rbzero.pov.spi_buffer[14] ),
    .B(_03528_),
    .X(_03535_));
 sky130_fd_sc_hd__o211a_1 _19843_ (.A1(\rbzero.pov.spi_buffer[15] ),
    .A2(_03527_),
    .B1(_03535_),
    .C1(_03533_),
    .X(_01051_));
 sky130_fd_sc_hd__or2_1 _19844_ (.A(\rbzero.pov.spi_buffer[15] ),
    .B(_03528_),
    .X(_03536_));
 sky130_fd_sc_hd__o211a_1 _19845_ (.A1(\rbzero.pov.spi_buffer[16] ),
    .A2(_03527_),
    .B1(_03536_),
    .C1(_03533_),
    .X(_01052_));
 sky130_fd_sc_hd__or2_1 _19846_ (.A(\rbzero.pov.spi_buffer[16] ),
    .B(_03528_),
    .X(_03537_));
 sky130_fd_sc_hd__o211a_1 _19847_ (.A1(\rbzero.pov.spi_buffer[17] ),
    .A2(_03527_),
    .B1(_03537_),
    .C1(_03533_),
    .X(_01053_));
 sky130_fd_sc_hd__or2_1 _19848_ (.A(\rbzero.pov.spi_buffer[17] ),
    .B(_03528_),
    .X(_03538_));
 sky130_fd_sc_hd__o211a_1 _19849_ (.A1(\rbzero.pov.spi_buffer[18] ),
    .A2(_03527_),
    .B1(_03538_),
    .C1(_03533_),
    .X(_01054_));
 sky130_fd_sc_hd__or2_1 _19850_ (.A(\rbzero.pov.spi_buffer[18] ),
    .B(_03528_),
    .X(_03539_));
 sky130_fd_sc_hd__o211a_1 _19851_ (.A1(\rbzero.pov.spi_buffer[19] ),
    .A2(_03527_),
    .B1(_03539_),
    .C1(_03533_),
    .X(_01055_));
 sky130_fd_sc_hd__buf_2 _19852_ (.A(_03511_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_2 _19853_ (.A(_03514_),
    .X(_03541_));
 sky130_fd_sc_hd__or2_1 _19854_ (.A(\rbzero.pov.spi_buffer[19] ),
    .B(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__o211a_1 _19855_ (.A1(\rbzero.pov.spi_buffer[20] ),
    .A2(_03540_),
    .B1(_03542_),
    .C1(_03533_),
    .X(_01056_));
 sky130_fd_sc_hd__or2_1 _19856_ (.A(\rbzero.pov.spi_buffer[20] ),
    .B(_03541_),
    .X(_03543_));
 sky130_fd_sc_hd__o211a_1 _19857_ (.A1(\rbzero.pov.spi_buffer[21] ),
    .A2(_03540_),
    .B1(_03543_),
    .C1(_03533_),
    .X(_01057_));
 sky130_fd_sc_hd__or2_1 _19858_ (.A(\rbzero.pov.spi_buffer[21] ),
    .B(_03541_),
    .X(_03544_));
 sky130_fd_sc_hd__o211a_1 _19859_ (.A1(\rbzero.pov.spi_buffer[22] ),
    .A2(_03540_),
    .B1(_03544_),
    .C1(_03533_),
    .X(_01058_));
 sky130_fd_sc_hd__or2_1 _19860_ (.A(\rbzero.pov.spi_buffer[22] ),
    .B(_03541_),
    .X(_03545_));
 sky130_fd_sc_hd__buf_2 _19861_ (.A(_02638_),
    .X(_03546_));
 sky130_fd_sc_hd__o211a_1 _19862_ (.A1(\rbzero.pov.spi_buffer[23] ),
    .A2(_03540_),
    .B1(_03545_),
    .C1(_03546_),
    .X(_01059_));
 sky130_fd_sc_hd__or2_1 _19863_ (.A(\rbzero.pov.spi_buffer[23] ),
    .B(_03541_),
    .X(_03547_));
 sky130_fd_sc_hd__o211a_1 _19864_ (.A1(\rbzero.pov.spi_buffer[24] ),
    .A2(_03540_),
    .B1(_03547_),
    .C1(_03546_),
    .X(_01060_));
 sky130_fd_sc_hd__or2_1 _19865_ (.A(\rbzero.pov.spi_buffer[24] ),
    .B(_03541_),
    .X(_03548_));
 sky130_fd_sc_hd__o211a_1 _19866_ (.A1(\rbzero.pov.spi_buffer[25] ),
    .A2(_03540_),
    .B1(_03548_),
    .C1(_03546_),
    .X(_01061_));
 sky130_fd_sc_hd__or2_1 _19867_ (.A(\rbzero.pov.spi_buffer[25] ),
    .B(_03541_),
    .X(_03549_));
 sky130_fd_sc_hd__o211a_1 _19868_ (.A1(\rbzero.pov.spi_buffer[26] ),
    .A2(_03540_),
    .B1(_03549_),
    .C1(_03546_),
    .X(_01062_));
 sky130_fd_sc_hd__or2_1 _19869_ (.A(\rbzero.pov.spi_buffer[26] ),
    .B(_03541_),
    .X(_03550_));
 sky130_fd_sc_hd__o211a_1 _19870_ (.A1(\rbzero.pov.spi_buffer[27] ),
    .A2(_03540_),
    .B1(_03550_),
    .C1(_03546_),
    .X(_01063_));
 sky130_fd_sc_hd__or2_1 _19871_ (.A(\rbzero.pov.spi_buffer[27] ),
    .B(_03541_),
    .X(_03551_));
 sky130_fd_sc_hd__o211a_1 _19872_ (.A1(\rbzero.pov.spi_buffer[28] ),
    .A2(_03540_),
    .B1(_03551_),
    .C1(_03546_),
    .X(_01064_));
 sky130_fd_sc_hd__or2_1 _19873_ (.A(\rbzero.pov.spi_buffer[28] ),
    .B(_03541_),
    .X(_03552_));
 sky130_fd_sc_hd__o211a_1 _19874_ (.A1(\rbzero.pov.spi_buffer[29] ),
    .A2(_03540_),
    .B1(_03552_),
    .C1(_03546_),
    .X(_01065_));
 sky130_fd_sc_hd__buf_2 _19875_ (.A(_03511_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_2 _19876_ (.A(_03514_),
    .X(_03554_));
 sky130_fd_sc_hd__or2_1 _19877_ (.A(\rbzero.pov.spi_buffer[29] ),
    .B(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__o211a_1 _19878_ (.A1(\rbzero.pov.spi_buffer[30] ),
    .A2(_03553_),
    .B1(_03555_),
    .C1(_03546_),
    .X(_01066_));
 sky130_fd_sc_hd__or2_1 _19879_ (.A(\rbzero.pov.spi_buffer[30] ),
    .B(_03554_),
    .X(_03556_));
 sky130_fd_sc_hd__o211a_1 _19880_ (.A1(\rbzero.pov.spi_buffer[31] ),
    .A2(_03553_),
    .B1(_03556_),
    .C1(_03546_),
    .X(_01067_));
 sky130_fd_sc_hd__or2_1 _19881_ (.A(\rbzero.pov.spi_buffer[31] ),
    .B(_03554_),
    .X(_03557_));
 sky130_fd_sc_hd__o211a_1 _19882_ (.A1(\rbzero.pov.spi_buffer[32] ),
    .A2(_03553_),
    .B1(_03557_),
    .C1(_03546_),
    .X(_01068_));
 sky130_fd_sc_hd__or2_1 _19883_ (.A(\rbzero.pov.spi_buffer[32] ),
    .B(_03554_),
    .X(_03558_));
 sky130_fd_sc_hd__buf_2 _19884_ (.A(_02638_),
    .X(_03559_));
 sky130_fd_sc_hd__o211a_1 _19885_ (.A1(\rbzero.pov.spi_buffer[33] ),
    .A2(_03553_),
    .B1(_03558_),
    .C1(_03559_),
    .X(_01069_));
 sky130_fd_sc_hd__or2_1 _19886_ (.A(\rbzero.pov.spi_buffer[33] ),
    .B(_03554_),
    .X(_03560_));
 sky130_fd_sc_hd__o211a_1 _19887_ (.A1(\rbzero.pov.spi_buffer[34] ),
    .A2(_03553_),
    .B1(_03560_),
    .C1(_03559_),
    .X(_01070_));
 sky130_fd_sc_hd__or2_1 _19888_ (.A(\rbzero.pov.spi_buffer[34] ),
    .B(_03554_),
    .X(_03561_));
 sky130_fd_sc_hd__o211a_1 _19889_ (.A1(\rbzero.pov.spi_buffer[35] ),
    .A2(_03553_),
    .B1(_03561_),
    .C1(_03559_),
    .X(_01071_));
 sky130_fd_sc_hd__or2_1 _19890_ (.A(\rbzero.pov.spi_buffer[35] ),
    .B(_03554_),
    .X(_03562_));
 sky130_fd_sc_hd__o211a_1 _19891_ (.A1(\rbzero.pov.spi_buffer[36] ),
    .A2(_03553_),
    .B1(_03562_),
    .C1(_03559_),
    .X(_01072_));
 sky130_fd_sc_hd__or2_1 _19892_ (.A(\rbzero.pov.spi_buffer[36] ),
    .B(_03554_),
    .X(_03563_));
 sky130_fd_sc_hd__o211a_1 _19893_ (.A1(\rbzero.pov.spi_buffer[37] ),
    .A2(_03553_),
    .B1(_03563_),
    .C1(_03559_),
    .X(_01073_));
 sky130_fd_sc_hd__or2_1 _19894_ (.A(\rbzero.pov.spi_buffer[37] ),
    .B(_03554_),
    .X(_03564_));
 sky130_fd_sc_hd__o211a_1 _19895_ (.A1(\rbzero.pov.spi_buffer[38] ),
    .A2(_03553_),
    .B1(_03564_),
    .C1(_03559_),
    .X(_01074_));
 sky130_fd_sc_hd__or2_1 _19896_ (.A(\rbzero.pov.spi_buffer[38] ),
    .B(_03554_),
    .X(_03565_));
 sky130_fd_sc_hd__o211a_1 _19897_ (.A1(\rbzero.pov.spi_buffer[39] ),
    .A2(_03553_),
    .B1(_03565_),
    .C1(_03559_),
    .X(_01075_));
 sky130_fd_sc_hd__buf_2 _19898_ (.A(_03511_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_2 _19899_ (.A(_03514_),
    .X(_03567_));
 sky130_fd_sc_hd__or2_1 _19900_ (.A(\rbzero.pov.spi_buffer[39] ),
    .B(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__o211a_1 _19901_ (.A1(\rbzero.pov.spi_buffer[40] ),
    .A2(_03566_),
    .B1(_03568_),
    .C1(_03559_),
    .X(_01076_));
 sky130_fd_sc_hd__or2_1 _19902_ (.A(\rbzero.pov.spi_buffer[40] ),
    .B(_03567_),
    .X(_03569_));
 sky130_fd_sc_hd__o211a_1 _19903_ (.A1(\rbzero.pov.spi_buffer[41] ),
    .A2(_03566_),
    .B1(_03569_),
    .C1(_03559_),
    .X(_01077_));
 sky130_fd_sc_hd__or2_1 _19904_ (.A(\rbzero.pov.spi_buffer[41] ),
    .B(_03567_),
    .X(_03570_));
 sky130_fd_sc_hd__o211a_1 _19905_ (.A1(\rbzero.pov.spi_buffer[42] ),
    .A2(_03566_),
    .B1(_03570_),
    .C1(_03559_),
    .X(_01078_));
 sky130_fd_sc_hd__or2_1 _19906_ (.A(\rbzero.pov.spi_buffer[42] ),
    .B(_03567_),
    .X(_03571_));
 sky130_fd_sc_hd__buf_2 _19907_ (.A(_02638_),
    .X(_03572_));
 sky130_fd_sc_hd__o211a_1 _19908_ (.A1(\rbzero.pov.spi_buffer[43] ),
    .A2(_03566_),
    .B1(_03571_),
    .C1(_03572_),
    .X(_01079_));
 sky130_fd_sc_hd__or2_1 _19909_ (.A(\rbzero.pov.spi_buffer[43] ),
    .B(_03567_),
    .X(_03573_));
 sky130_fd_sc_hd__o211a_1 _19910_ (.A1(\rbzero.pov.spi_buffer[44] ),
    .A2(_03566_),
    .B1(_03573_),
    .C1(_03572_),
    .X(_01080_));
 sky130_fd_sc_hd__or2_1 _19911_ (.A(\rbzero.pov.spi_buffer[44] ),
    .B(_03567_),
    .X(_03574_));
 sky130_fd_sc_hd__o211a_1 _19912_ (.A1(\rbzero.pov.spi_buffer[45] ),
    .A2(_03566_),
    .B1(_03574_),
    .C1(_03572_),
    .X(_01081_));
 sky130_fd_sc_hd__or2_1 _19913_ (.A(\rbzero.pov.spi_buffer[45] ),
    .B(_03567_),
    .X(_03575_));
 sky130_fd_sc_hd__o211a_1 _19914_ (.A1(\rbzero.pov.spi_buffer[46] ),
    .A2(_03566_),
    .B1(_03575_),
    .C1(_03572_),
    .X(_01082_));
 sky130_fd_sc_hd__or2_1 _19915_ (.A(\rbzero.pov.spi_buffer[46] ),
    .B(_03567_),
    .X(_03576_));
 sky130_fd_sc_hd__o211a_1 _19916_ (.A1(\rbzero.pov.spi_buffer[47] ),
    .A2(_03566_),
    .B1(_03576_),
    .C1(_03572_),
    .X(_01083_));
 sky130_fd_sc_hd__or2_1 _19917_ (.A(\rbzero.pov.spi_buffer[47] ),
    .B(_03567_),
    .X(_03577_));
 sky130_fd_sc_hd__o211a_1 _19918_ (.A1(\rbzero.pov.spi_buffer[48] ),
    .A2(_03566_),
    .B1(_03577_),
    .C1(_03572_),
    .X(_01084_));
 sky130_fd_sc_hd__or2_1 _19919_ (.A(\rbzero.pov.spi_buffer[48] ),
    .B(_03567_),
    .X(_03578_));
 sky130_fd_sc_hd__o211a_1 _19920_ (.A1(\rbzero.pov.spi_buffer[49] ),
    .A2(_03566_),
    .B1(_03578_),
    .C1(_03572_),
    .X(_01085_));
 sky130_fd_sc_hd__buf_2 _19921_ (.A(_03511_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_2 _19922_ (.A(_03514_),
    .X(_03580_));
 sky130_fd_sc_hd__or2_1 _19923_ (.A(\rbzero.pov.spi_buffer[49] ),
    .B(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__o211a_1 _19924_ (.A1(\rbzero.pov.spi_buffer[50] ),
    .A2(_03579_),
    .B1(_03581_),
    .C1(_03572_),
    .X(_01086_));
 sky130_fd_sc_hd__or2_1 _19925_ (.A(\rbzero.pov.spi_buffer[50] ),
    .B(_03580_),
    .X(_03582_));
 sky130_fd_sc_hd__o211a_1 _19926_ (.A1(\rbzero.pov.spi_buffer[51] ),
    .A2(_03579_),
    .B1(_03582_),
    .C1(_03572_),
    .X(_01087_));
 sky130_fd_sc_hd__or2_1 _19927_ (.A(\rbzero.pov.spi_buffer[51] ),
    .B(_03580_),
    .X(_03583_));
 sky130_fd_sc_hd__o211a_1 _19928_ (.A1(\rbzero.pov.spi_buffer[52] ),
    .A2(_03579_),
    .B1(_03583_),
    .C1(_03572_),
    .X(_01088_));
 sky130_fd_sc_hd__or2_1 _19929_ (.A(\rbzero.pov.spi_buffer[52] ),
    .B(_03580_),
    .X(_03584_));
 sky130_fd_sc_hd__buf_2 _19930_ (.A(_02638_),
    .X(_03585_));
 sky130_fd_sc_hd__o211a_1 _19931_ (.A1(\rbzero.pov.spi_buffer[53] ),
    .A2(_03579_),
    .B1(_03584_),
    .C1(_03585_),
    .X(_01089_));
 sky130_fd_sc_hd__or2_1 _19932_ (.A(\rbzero.pov.spi_buffer[53] ),
    .B(_03580_),
    .X(_03586_));
 sky130_fd_sc_hd__o211a_1 _19933_ (.A1(\rbzero.pov.spi_buffer[54] ),
    .A2(_03579_),
    .B1(_03586_),
    .C1(_03585_),
    .X(_01090_));
 sky130_fd_sc_hd__or2_1 _19934_ (.A(\rbzero.pov.spi_buffer[54] ),
    .B(_03580_),
    .X(_03587_));
 sky130_fd_sc_hd__o211a_1 _19935_ (.A1(\rbzero.pov.spi_buffer[55] ),
    .A2(_03579_),
    .B1(_03587_),
    .C1(_03585_),
    .X(_01091_));
 sky130_fd_sc_hd__or2_1 _19936_ (.A(\rbzero.pov.spi_buffer[55] ),
    .B(_03580_),
    .X(_03588_));
 sky130_fd_sc_hd__o211a_1 _19937_ (.A1(\rbzero.pov.spi_buffer[56] ),
    .A2(_03579_),
    .B1(_03588_),
    .C1(_03585_),
    .X(_01092_));
 sky130_fd_sc_hd__or2_1 _19938_ (.A(\rbzero.pov.spi_buffer[56] ),
    .B(_03580_),
    .X(_03589_));
 sky130_fd_sc_hd__o211a_1 _19939_ (.A1(\rbzero.pov.spi_buffer[57] ),
    .A2(_03579_),
    .B1(_03589_),
    .C1(_03585_),
    .X(_01093_));
 sky130_fd_sc_hd__or2_1 _19940_ (.A(\rbzero.pov.spi_buffer[57] ),
    .B(_03580_),
    .X(_03590_));
 sky130_fd_sc_hd__o211a_1 _19941_ (.A1(\rbzero.pov.spi_buffer[58] ),
    .A2(_03579_),
    .B1(_03590_),
    .C1(_03585_),
    .X(_01094_));
 sky130_fd_sc_hd__or2_1 _19942_ (.A(\rbzero.pov.spi_buffer[58] ),
    .B(_03580_),
    .X(_03591_));
 sky130_fd_sc_hd__o211a_1 _19943_ (.A1(\rbzero.pov.spi_buffer[59] ),
    .A2(_03579_),
    .B1(_03591_),
    .C1(_03585_),
    .X(_01095_));
 sky130_fd_sc_hd__buf_2 _19944_ (.A(_03510_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_2 _19945_ (.A(_03513_),
    .X(_03593_));
 sky130_fd_sc_hd__or2_1 _19946_ (.A(\rbzero.pov.spi_buffer[59] ),
    .B(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__o211a_1 _19947_ (.A1(\rbzero.pov.spi_buffer[60] ),
    .A2(_03592_),
    .B1(_03594_),
    .C1(_03585_),
    .X(_01096_));
 sky130_fd_sc_hd__or2_1 _19948_ (.A(\rbzero.pov.spi_buffer[60] ),
    .B(_03593_),
    .X(_03595_));
 sky130_fd_sc_hd__o211a_1 _19949_ (.A1(\rbzero.pov.spi_buffer[61] ),
    .A2(_03592_),
    .B1(_03595_),
    .C1(_03585_),
    .X(_01097_));
 sky130_fd_sc_hd__or2_1 _19950_ (.A(\rbzero.pov.spi_buffer[61] ),
    .B(_03593_),
    .X(_03596_));
 sky130_fd_sc_hd__o211a_1 _19951_ (.A1(\rbzero.pov.spi_buffer[62] ),
    .A2(_03592_),
    .B1(_03596_),
    .C1(_03585_),
    .X(_01098_));
 sky130_fd_sc_hd__or2_1 _19952_ (.A(\rbzero.pov.spi_buffer[62] ),
    .B(_03593_),
    .X(_03597_));
 sky130_fd_sc_hd__buf_2 _19953_ (.A(_02638_),
    .X(_03598_));
 sky130_fd_sc_hd__o211a_1 _19954_ (.A1(\rbzero.pov.spi_buffer[63] ),
    .A2(_03592_),
    .B1(_03597_),
    .C1(_03598_),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _19955_ (.A(\rbzero.pov.spi_buffer[63] ),
    .B(_03593_),
    .X(_03599_));
 sky130_fd_sc_hd__o211a_1 _19956_ (.A1(\rbzero.pov.spi_buffer[64] ),
    .A2(_03592_),
    .B1(_03599_),
    .C1(_03598_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_1 _19957_ (.A(\rbzero.pov.spi_buffer[64] ),
    .B(_03593_),
    .X(_03600_));
 sky130_fd_sc_hd__o211a_1 _19958_ (.A1(\rbzero.pov.spi_buffer[65] ),
    .A2(_03592_),
    .B1(_03600_),
    .C1(_03598_),
    .X(_01101_));
 sky130_fd_sc_hd__or2_1 _19959_ (.A(\rbzero.pov.spi_buffer[65] ),
    .B(_03593_),
    .X(_03601_));
 sky130_fd_sc_hd__o211a_1 _19960_ (.A1(\rbzero.pov.spi_buffer[66] ),
    .A2(_03592_),
    .B1(_03601_),
    .C1(_03598_),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _19961_ (.A(\rbzero.pov.spi_buffer[66] ),
    .B(_03593_),
    .X(_03602_));
 sky130_fd_sc_hd__o211a_1 _19962_ (.A1(\rbzero.pov.spi_buffer[67] ),
    .A2(_03592_),
    .B1(_03602_),
    .C1(_03598_),
    .X(_01103_));
 sky130_fd_sc_hd__or2_1 _19963_ (.A(\rbzero.pov.spi_buffer[67] ),
    .B(_03593_),
    .X(_03603_));
 sky130_fd_sc_hd__o211a_1 _19964_ (.A1(\rbzero.pov.spi_buffer[68] ),
    .A2(_03592_),
    .B1(_03603_),
    .C1(_03598_),
    .X(_01104_));
 sky130_fd_sc_hd__or2_1 _19965_ (.A(\rbzero.pov.spi_buffer[68] ),
    .B(_03593_),
    .X(_03604_));
 sky130_fd_sc_hd__o211a_1 _19966_ (.A1(\rbzero.pov.spi_buffer[69] ),
    .A2(_03592_),
    .B1(_03604_),
    .C1(_03598_),
    .X(_01105_));
 sky130_fd_sc_hd__or2_1 _19967_ (.A(\rbzero.pov.spi_buffer[69] ),
    .B(_03514_),
    .X(_03605_));
 sky130_fd_sc_hd__o211a_1 _19968_ (.A1(\rbzero.pov.spi_buffer[70] ),
    .A2(_03511_),
    .B1(_03605_),
    .C1(_03598_),
    .X(_01106_));
 sky130_fd_sc_hd__or2_1 _19969_ (.A(\rbzero.pov.spi_buffer[70] ),
    .B(_03514_),
    .X(_03606_));
 sky130_fd_sc_hd__o211a_1 _19970_ (.A1(\rbzero.pov.spi_buffer[71] ),
    .A2(_03511_),
    .B1(_03606_),
    .C1(_03598_),
    .X(_01107_));
 sky130_fd_sc_hd__or2_1 _19971_ (.A(\rbzero.pov.spi_buffer[71] ),
    .B(_03514_),
    .X(_03607_));
 sky130_fd_sc_hd__o211a_1 _19972_ (.A1(\rbzero.pov.spi_buffer[72] ),
    .A2(_03511_),
    .B1(_03607_),
    .C1(_03598_),
    .X(_01108_));
 sky130_fd_sc_hd__or2_1 _19973_ (.A(\rbzero.pov.spi_buffer[72] ),
    .B(_03514_),
    .X(_03608_));
 sky130_fd_sc_hd__o211a_1 _19974_ (.A1(\rbzero.pov.spi_buffer[73] ),
    .A2(_03511_),
    .B1(_03608_),
    .C1(_02901_),
    .X(_01109_));
 sky130_fd_sc_hd__buf_1 _19975_ (.A(clknet_1_0__leaf__05762_),
    .X(_03609_));
 sky130_fd_sc_hd__buf_1 _19976_ (.A(clknet_1_0__leaf__03609_),
    .X(_03610_));
 sky130_fd_sc_hd__inv_2 _19978__29 (.A(clknet_1_0__leaf__03610_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _19979__30 (.A(clknet_1_0__leaf__03610_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _19980__31 (.A(clknet_1_0__leaf__03610_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _19981__32 (.A(clknet_1_1__leaf__03610_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _19982__33 (.A(clknet_1_1__leaf__03610_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _19983__34 (.A(clknet_1_1__leaf__03610_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _19984__35 (.A(clknet_1_1__leaf__03610_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _19985__36 (.A(clknet_1_1__leaf__03610_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _19986__37 (.A(clknet_1_1__leaf__03610_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _19988__38 (.A(clknet_1_1__leaf__03611_),
    .Y(net164));
 sky130_fd_sc_hd__buf_1 _19987_ (.A(clknet_1_1__leaf__03609_),
    .X(_03611_));
 sky130_fd_sc_hd__inv_2 _19989__39 (.A(clknet_1_1__leaf__03611_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _19990__40 (.A(clknet_1_1__leaf__03611_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _19991__41 (.A(clknet_1_0__leaf__03611_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _19992__42 (.A(clknet_1_0__leaf__03611_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _19993__43 (.A(clknet_1_0__leaf__03611_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _19994__44 (.A(clknet_1_0__leaf__03611_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _19995__45 (.A(clknet_1_1__leaf__03611_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _19996__46 (.A(clknet_1_1__leaf__03611_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _19997__47 (.A(clknet_1_0__leaf__03611_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _19999__48 (.A(clknet_1_1__leaf__03612_),
    .Y(net174));
 sky130_fd_sc_hd__buf_1 _19998_ (.A(clknet_1_0__leaf__03609_),
    .X(_03612_));
 sky130_fd_sc_hd__inv_2 _20000__49 (.A(clknet_1_0__leaf__03612_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _20001__50 (.A(clknet_1_0__leaf__03612_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _20002__51 (.A(clknet_1_0__leaf__03612_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _20003__52 (.A(clknet_1_1__leaf__03612_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _20004__53 (.A(clknet_1_0__leaf__03612_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _20005__54 (.A(clknet_1_0__leaf__03612_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _20006__55 (.A(clknet_1_0__leaf__03612_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _20007__56 (.A(clknet_1_1__leaf__03612_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _20008__57 (.A(clknet_1_1__leaf__03612_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _20010__58 (.A(clknet_1_1__leaf__03613_),
    .Y(net184));
 sky130_fd_sc_hd__buf_1 _20009_ (.A(clknet_1_0__leaf__03609_),
    .X(_03613_));
 sky130_fd_sc_hd__inv_2 _20011__59 (.A(clknet_1_0__leaf__03613_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _20012__60 (.A(clknet_1_0__leaf__03613_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _20013__61 (.A(clknet_1_0__leaf__03613_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _20014__62 (.A(clknet_1_0__leaf__03613_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _20015__63 (.A(clknet_1_0__leaf__03613_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _20016__64 (.A(clknet_1_1__leaf__03613_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _20017__65 (.A(clknet_1_1__leaf__03613_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _20018__66 (.A(clknet_1_1__leaf__03613_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _20019__67 (.A(clknet_1_1__leaf__03613_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _20021__68 (.A(clknet_1_1__leaf__03614_),
    .Y(net194));
 sky130_fd_sc_hd__buf_1 _20020_ (.A(clknet_1_0__leaf__03609_),
    .X(_03614_));
 sky130_fd_sc_hd__inv_2 _20022__69 (.A(clknet_1_1__leaf__03614_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _20023__70 (.A(clknet_1_1__leaf__03614_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _20024__71 (.A(clknet_1_1__leaf__03614_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _20025__72 (.A(clknet_1_1__leaf__03614_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _20026__73 (.A(clknet_1_0__leaf__03614_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _20027__74 (.A(clknet_1_0__leaf__03614_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _20028__75 (.A(clknet_1_0__leaf__03614_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _20029__76 (.A(clknet_1_0__leaf__03614_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _20030__77 (.A(clknet_1_0__leaf__03614_),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _20032__78 (.A(clknet_1_0__leaf__03615_),
    .Y(net204));
 sky130_fd_sc_hd__buf_1 _20031_ (.A(clknet_1_0__leaf__03609_),
    .X(_03615_));
 sky130_fd_sc_hd__inv_2 _20033__79 (.A(clknet_1_1__leaf__03615_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _20034__80 (.A(clknet_1_1__leaf__03615_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _20035__81 (.A(clknet_1_1__leaf__03615_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _20036__82 (.A(clknet_1_1__leaf__03615_),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _20037__83 (.A(clknet_1_1__leaf__03615_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _20038__84 (.A(clknet_1_0__leaf__03615_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _20039__85 (.A(clknet_1_0__leaf__03615_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _20040__86 (.A(clknet_1_0__leaf__03615_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _20041__87 (.A(clknet_1_0__leaf__03615_),
    .Y(net213));
 sky130_fd_sc_hd__inv_2 _20044__88 (.A(clknet_1_0__leaf__03617_),
    .Y(net214));
 sky130_fd_sc_hd__buf_1 _20042_ (.A(clknet_1_1__leaf__05762_),
    .X(_03616_));
 sky130_fd_sc_hd__buf_1 _20043_ (.A(clknet_1_0__leaf__03616_),
    .X(_03617_));
 sky130_fd_sc_hd__inv_2 _20045__89 (.A(clknet_1_0__leaf__03617_),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _20046__90 (.A(clknet_1_0__leaf__03617_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _20047__91 (.A(clknet_1_0__leaf__03617_),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _20340__92 (.A(clknet_1_1__leaf__03617_),
    .Y(net218));
 sky130_fd_sc_hd__buf_4 _20048_ (.A(\rbzero.pov.spi_done ),
    .X(_03618_));
 sky130_fd_sc_hd__o211a_1 _20049_ (.A1(_03618_),
    .A2(\rbzero.pov.ready ),
    .B1(_02901_),
    .C1(_03358_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _20050_ (.A0(\rbzero.pov.ready_buffer[0] ),
    .A1(\rbzero.pov.spi_buffer[0] ),
    .S(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__and2_1 _20051_ (.A(_08093_),
    .B(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_1 _20052_ (.A(_03620_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _20053_ (.A0(\rbzero.pov.ready_buffer[1] ),
    .A1(\rbzero.pov.spi_buffer[1] ),
    .S(_03618_),
    .X(_03621_));
 sky130_fd_sc_hd__and2_1 _20054_ (.A(_08093_),
    .B(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__clkbuf_1 _20055_ (.A(_03622_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _20056_ (.A0(\rbzero.pov.ready_buffer[2] ),
    .A1(\rbzero.pov.spi_buffer[2] ),
    .S(_03618_),
    .X(_03623_));
 sky130_fd_sc_hd__and2_1 _20057_ (.A(_08093_),
    .B(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__clkbuf_1 _20058_ (.A(_03624_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _20059_ (.A0(\rbzero.pov.ready_buffer[3] ),
    .A1(\rbzero.pov.spi_buffer[3] ),
    .S(_03618_),
    .X(_03625_));
 sky130_fd_sc_hd__and2_1 _20060_ (.A(_08093_),
    .B(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _20061_ (.A(_03626_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _20062_ (.A0(\rbzero.pov.ready_buffer[4] ),
    .A1(\rbzero.pov.spi_buffer[4] ),
    .S(_03618_),
    .X(_03627_));
 sky130_fd_sc_hd__and2_1 _20063_ (.A(_08093_),
    .B(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__clkbuf_1 _20064_ (.A(_03628_),
    .X(_01179_));
 sky130_fd_sc_hd__clkbuf_2 _20065_ (.A(_08092_),
    .X(_03629_));
 sky130_fd_sc_hd__mux2_1 _20066_ (.A0(\rbzero.pov.ready_buffer[5] ),
    .A1(\rbzero.pov.spi_buffer[5] ),
    .S(_03618_),
    .X(_03630_));
 sky130_fd_sc_hd__and2_1 _20067_ (.A(_03629_),
    .B(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _20068_ (.A(_03631_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _20069_ (.A0(\rbzero.pov.ready_buffer[6] ),
    .A1(\rbzero.pov.spi_buffer[6] ),
    .S(_03618_),
    .X(_03632_));
 sky130_fd_sc_hd__and2_1 _20070_ (.A(_03629_),
    .B(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_1 _20071_ (.A(_03633_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _20072_ (.A0(\rbzero.pov.ready_buffer[7] ),
    .A1(\rbzero.pov.spi_buffer[7] ),
    .S(_03618_),
    .X(_03634_));
 sky130_fd_sc_hd__and2_1 _20073_ (.A(_03629_),
    .B(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_1 _20074_ (.A(_03635_),
    .X(_01182_));
 sky130_fd_sc_hd__buf_4 _20075_ (.A(\rbzero.pov.spi_done ),
    .X(_03636_));
 sky130_fd_sc_hd__clkbuf_4 _20076_ (.A(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__mux2_1 _20077_ (.A0(\rbzero.pov.ready_buffer[8] ),
    .A1(\rbzero.pov.spi_buffer[8] ),
    .S(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__and2_1 _20078_ (.A(_03629_),
    .B(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__clkbuf_1 _20079_ (.A(_03639_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _20080_ (.A0(\rbzero.pov.ready_buffer[9] ),
    .A1(\rbzero.pov.spi_buffer[9] ),
    .S(_03637_),
    .X(_03640_));
 sky130_fd_sc_hd__and2_1 _20081_ (.A(_03629_),
    .B(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _20082_ (.A(_03641_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _20083_ (.A0(\rbzero.pov.ready_buffer[10] ),
    .A1(\rbzero.pov.spi_buffer[10] ),
    .S(_03637_),
    .X(_03642_));
 sky130_fd_sc_hd__and2_1 _20084_ (.A(_03629_),
    .B(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__clkbuf_1 _20085_ (.A(_03643_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _20086_ (.A0(\rbzero.pov.ready_buffer[11] ),
    .A1(\rbzero.pov.spi_buffer[11] ),
    .S(_03637_),
    .X(_03644_));
 sky130_fd_sc_hd__and2_1 _20087_ (.A(_03629_),
    .B(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _20088_ (.A(_03645_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _20089_ (.A0(\rbzero.pov.ready_buffer[12] ),
    .A1(\rbzero.pov.spi_buffer[12] ),
    .S(_03637_),
    .X(_03646_));
 sky130_fd_sc_hd__and2_1 _20090_ (.A(_03629_),
    .B(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_1 _20091_ (.A(_03647_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _20092_ (.A0(\rbzero.pov.ready_buffer[13] ),
    .A1(\rbzero.pov.spi_buffer[13] ),
    .S(_03637_),
    .X(_03648_));
 sky130_fd_sc_hd__and2_1 _20093_ (.A(_03629_),
    .B(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _20094_ (.A(_03649_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _20095_ (.A0(\rbzero.pov.ready_buffer[14] ),
    .A1(\rbzero.pov.spi_buffer[14] ),
    .S(_03637_),
    .X(_03650_));
 sky130_fd_sc_hd__and2_1 _20096_ (.A(_03629_),
    .B(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _20097_ (.A(_03651_),
    .X(_01189_));
 sky130_fd_sc_hd__clkbuf_2 _20098_ (.A(_08092_),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _20099_ (.A0(\rbzero.pov.ready_buffer[15] ),
    .A1(\rbzero.pov.spi_buffer[15] ),
    .S(_03637_),
    .X(_03653_));
 sky130_fd_sc_hd__and2_1 _20100_ (.A(_03652_),
    .B(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__clkbuf_1 _20101_ (.A(_03654_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _20102_ (.A0(\rbzero.pov.ready_buffer[16] ),
    .A1(\rbzero.pov.spi_buffer[16] ),
    .S(_03637_),
    .X(_03655_));
 sky130_fd_sc_hd__and2_1 _20103_ (.A(_03652_),
    .B(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_1 _20104_ (.A(_03656_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _20105_ (.A0(\rbzero.pov.ready_buffer[17] ),
    .A1(\rbzero.pov.spi_buffer[17] ),
    .S(_03637_),
    .X(_03657_));
 sky130_fd_sc_hd__and2_1 _20106_ (.A(_03652_),
    .B(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_1 _20107_ (.A(_03658_),
    .X(_01192_));
 sky130_fd_sc_hd__clkbuf_4 _20108_ (.A(_03636_),
    .X(_03659_));
 sky130_fd_sc_hd__mux2_1 _20109_ (.A0(\rbzero.pov.ready_buffer[18] ),
    .A1(\rbzero.pov.spi_buffer[18] ),
    .S(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__and2_1 _20110_ (.A(_03652_),
    .B(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_1 _20111_ (.A(_03661_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _20112_ (.A0(\rbzero.pov.ready_buffer[19] ),
    .A1(\rbzero.pov.spi_buffer[19] ),
    .S(_03659_),
    .X(_03662_));
 sky130_fd_sc_hd__and2_1 _20113_ (.A(_03652_),
    .B(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__clkbuf_1 _20114_ (.A(_03663_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _20115_ (.A0(\rbzero.pov.ready_buffer[20] ),
    .A1(\rbzero.pov.spi_buffer[20] ),
    .S(_03659_),
    .X(_03664_));
 sky130_fd_sc_hd__and2_1 _20116_ (.A(_03652_),
    .B(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__clkbuf_1 _20117_ (.A(_03665_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _20118_ (.A0(\rbzero.pov.ready_buffer[21] ),
    .A1(\rbzero.pov.spi_buffer[21] ),
    .S(_03659_),
    .X(_03666_));
 sky130_fd_sc_hd__and2_1 _20119_ (.A(_03652_),
    .B(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__clkbuf_1 _20120_ (.A(_03667_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _20121_ (.A0(\rbzero.pov.ready_buffer[22] ),
    .A1(\rbzero.pov.spi_buffer[22] ),
    .S(_03659_),
    .X(_03668_));
 sky130_fd_sc_hd__and2_1 _20122_ (.A(_03652_),
    .B(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_1 _20123_ (.A(_03669_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _20124_ (.A0(\rbzero.pov.ready_buffer[23] ),
    .A1(\rbzero.pov.spi_buffer[23] ),
    .S(_03659_),
    .X(_03670_));
 sky130_fd_sc_hd__and2_1 _20125_ (.A(_03652_),
    .B(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__clkbuf_1 _20126_ (.A(_03671_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _20127_ (.A0(\rbzero.pov.ready_buffer[24] ),
    .A1(\rbzero.pov.spi_buffer[24] ),
    .S(_03659_),
    .X(_03672_));
 sky130_fd_sc_hd__and2_1 _20128_ (.A(_03652_),
    .B(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__clkbuf_1 _20129_ (.A(_03673_),
    .X(_01199_));
 sky130_fd_sc_hd__clkbuf_2 _20130_ (.A(_08092_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _20131_ (.A0(\rbzero.pov.ready_buffer[25] ),
    .A1(\rbzero.pov.spi_buffer[25] ),
    .S(_03659_),
    .X(_03675_));
 sky130_fd_sc_hd__and2_1 _20132_ (.A(_03674_),
    .B(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__clkbuf_1 _20133_ (.A(_03676_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _20134_ (.A0(\rbzero.pov.ready_buffer[26] ),
    .A1(\rbzero.pov.spi_buffer[26] ),
    .S(_03659_),
    .X(_03677_));
 sky130_fd_sc_hd__and2_1 _20135_ (.A(_03674_),
    .B(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_1 _20136_ (.A(_03678_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _20137_ (.A0(\rbzero.pov.ready_buffer[27] ),
    .A1(\rbzero.pov.spi_buffer[27] ),
    .S(_03659_),
    .X(_03679_));
 sky130_fd_sc_hd__and2_1 _20138_ (.A(_03674_),
    .B(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_1 _20139_ (.A(_03680_),
    .X(_01202_));
 sky130_fd_sc_hd__clkbuf_4 _20140_ (.A(_03636_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _20141_ (.A0(\rbzero.pov.ready_buffer[28] ),
    .A1(\rbzero.pov.spi_buffer[28] ),
    .S(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__and2_1 _20142_ (.A(_03674_),
    .B(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _20143_ (.A(_03683_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _20144_ (.A0(\rbzero.pov.ready_buffer[29] ),
    .A1(\rbzero.pov.spi_buffer[29] ),
    .S(_03681_),
    .X(_03684_));
 sky130_fd_sc_hd__and2_1 _20145_ (.A(_03674_),
    .B(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__clkbuf_1 _20146_ (.A(_03685_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _20147_ (.A0(\rbzero.pov.ready_buffer[30] ),
    .A1(\rbzero.pov.spi_buffer[30] ),
    .S(_03681_),
    .X(_03686_));
 sky130_fd_sc_hd__and2_1 _20148_ (.A(_03674_),
    .B(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_1 _20149_ (.A(_03687_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _20150_ (.A0(\rbzero.pov.ready_buffer[31] ),
    .A1(\rbzero.pov.spi_buffer[31] ),
    .S(_03681_),
    .X(_03688_));
 sky130_fd_sc_hd__and2_1 _20151_ (.A(_03674_),
    .B(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _20152_ (.A(_03689_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _20153_ (.A0(\rbzero.pov.ready_buffer[32] ),
    .A1(\rbzero.pov.spi_buffer[32] ),
    .S(_03681_),
    .X(_03690_));
 sky130_fd_sc_hd__and2_1 _20154_ (.A(_03674_),
    .B(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__clkbuf_1 _20155_ (.A(_03691_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _20156_ (.A0(\rbzero.pov.ready_buffer[33] ),
    .A1(\rbzero.pov.spi_buffer[33] ),
    .S(_03681_),
    .X(_03692_));
 sky130_fd_sc_hd__and2_1 _20157_ (.A(_03674_),
    .B(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__clkbuf_1 _20158_ (.A(_03693_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _20159_ (.A0(\rbzero.pov.ready_buffer[34] ),
    .A1(\rbzero.pov.spi_buffer[34] ),
    .S(_03681_),
    .X(_03694_));
 sky130_fd_sc_hd__and2_1 _20160_ (.A(_03674_),
    .B(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_1 _20161_ (.A(_03695_),
    .X(_01209_));
 sky130_fd_sc_hd__buf_2 _20162_ (.A(_08092_),
    .X(_03696_));
 sky130_fd_sc_hd__mux2_1 _20163_ (.A0(\rbzero.pov.ready_buffer[35] ),
    .A1(\rbzero.pov.spi_buffer[35] ),
    .S(_03681_),
    .X(_03697_));
 sky130_fd_sc_hd__and2_1 _20164_ (.A(_03696_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_1 _20165_ (.A(_03698_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _20166_ (.A0(\rbzero.pov.ready_buffer[36] ),
    .A1(\rbzero.pov.spi_buffer[36] ),
    .S(_03681_),
    .X(_03699_));
 sky130_fd_sc_hd__and2_1 _20167_ (.A(_03696_),
    .B(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_1 _20168_ (.A(_03700_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _20169_ (.A0(\rbzero.pov.ready_buffer[37] ),
    .A1(\rbzero.pov.spi_buffer[37] ),
    .S(_03681_),
    .X(_03701_));
 sky130_fd_sc_hd__and2_1 _20170_ (.A(_03696_),
    .B(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__clkbuf_1 _20171_ (.A(_03702_),
    .X(_01212_));
 sky130_fd_sc_hd__buf_4 _20172_ (.A(_03636_),
    .X(_03703_));
 sky130_fd_sc_hd__mux2_1 _20173_ (.A0(\rbzero.pov.ready_buffer[38] ),
    .A1(\rbzero.pov.spi_buffer[38] ),
    .S(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__and2_1 _20174_ (.A(_03696_),
    .B(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_1 _20175_ (.A(_03705_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _20176_ (.A0(\rbzero.pov.ready_buffer[39] ),
    .A1(\rbzero.pov.spi_buffer[39] ),
    .S(_03703_),
    .X(_03706_));
 sky130_fd_sc_hd__and2_1 _20177_ (.A(_03696_),
    .B(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_1 _20178_ (.A(_03707_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _20179_ (.A0(\rbzero.pov.ready_buffer[40] ),
    .A1(\rbzero.pov.spi_buffer[40] ),
    .S(_03703_),
    .X(_03708_));
 sky130_fd_sc_hd__and2_1 _20180_ (.A(_03696_),
    .B(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_1 _20181_ (.A(_03709_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _20182_ (.A0(\rbzero.pov.ready_buffer[41] ),
    .A1(\rbzero.pov.spi_buffer[41] ),
    .S(_03703_),
    .X(_03710_));
 sky130_fd_sc_hd__and2_1 _20183_ (.A(_03696_),
    .B(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_1 _20184_ (.A(_03711_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _20185_ (.A0(\rbzero.pov.ready_buffer[42] ),
    .A1(\rbzero.pov.spi_buffer[42] ),
    .S(_03703_),
    .X(_03712_));
 sky130_fd_sc_hd__and2_1 _20186_ (.A(_03696_),
    .B(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _20187_ (.A(_03713_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _20188_ (.A0(\rbzero.pov.ready_buffer[43] ),
    .A1(\rbzero.pov.spi_buffer[43] ),
    .S(_03703_),
    .X(_03714_));
 sky130_fd_sc_hd__and2_1 _20189_ (.A(_03696_),
    .B(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_1 _20190_ (.A(_03715_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _20191_ (.A0(\rbzero.pov.ready_buffer[44] ),
    .A1(\rbzero.pov.spi_buffer[44] ),
    .S(_03703_),
    .X(_03716_));
 sky130_fd_sc_hd__and2_1 _20192_ (.A(_03696_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_1 _20193_ (.A(_03717_),
    .X(_01219_));
 sky130_fd_sc_hd__buf_2 _20194_ (.A(_08092_),
    .X(_03718_));
 sky130_fd_sc_hd__mux2_1 _20195_ (.A0(\rbzero.pov.ready_buffer[45] ),
    .A1(\rbzero.pov.spi_buffer[45] ),
    .S(_03703_),
    .X(_03719_));
 sky130_fd_sc_hd__and2_1 _20196_ (.A(_03718_),
    .B(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _20197_ (.A(_03720_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _20198_ (.A0(\rbzero.pov.ready_buffer[46] ),
    .A1(\rbzero.pov.spi_buffer[46] ),
    .S(_03703_),
    .X(_03721_));
 sky130_fd_sc_hd__and2_1 _20199_ (.A(_03718_),
    .B(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_1 _20200_ (.A(_03722_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _20201_ (.A0(\rbzero.pov.ready_buffer[47] ),
    .A1(\rbzero.pov.spi_buffer[47] ),
    .S(_03703_),
    .X(_03723_));
 sky130_fd_sc_hd__and2_1 _20202_ (.A(_03718_),
    .B(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _20203_ (.A(_03724_),
    .X(_01222_));
 sky130_fd_sc_hd__buf_4 _20204_ (.A(\rbzero.pov.spi_done ),
    .X(_03725_));
 sky130_fd_sc_hd__mux2_1 _20205_ (.A0(\rbzero.pov.ready_buffer[48] ),
    .A1(\rbzero.pov.spi_buffer[48] ),
    .S(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__and2_1 _20206_ (.A(_03718_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _20207_ (.A(_03727_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _20208_ (.A0(\rbzero.pov.ready_buffer[49] ),
    .A1(\rbzero.pov.spi_buffer[49] ),
    .S(_03725_),
    .X(_03728_));
 sky130_fd_sc_hd__and2_1 _20209_ (.A(_03718_),
    .B(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__clkbuf_1 _20210_ (.A(_03729_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _20211_ (.A0(\rbzero.pov.ready_buffer[50] ),
    .A1(\rbzero.pov.spi_buffer[50] ),
    .S(_03725_),
    .X(_03730_));
 sky130_fd_sc_hd__and2_1 _20212_ (.A(_03718_),
    .B(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_1 _20213_ (.A(_03731_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _20214_ (.A0(\rbzero.pov.ready_buffer[51] ),
    .A1(\rbzero.pov.spi_buffer[51] ),
    .S(_03725_),
    .X(_03732_));
 sky130_fd_sc_hd__and2_1 _20215_ (.A(_03718_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__clkbuf_1 _20216_ (.A(_03733_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _20217_ (.A0(\rbzero.pov.ready_buffer[52] ),
    .A1(\rbzero.pov.spi_buffer[52] ),
    .S(_03725_),
    .X(_03734_));
 sky130_fd_sc_hd__and2_1 _20218_ (.A(_03718_),
    .B(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__clkbuf_1 _20219_ (.A(_03735_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _20220_ (.A0(\rbzero.pov.ready_buffer[53] ),
    .A1(\rbzero.pov.spi_buffer[53] ),
    .S(_03725_),
    .X(_03736_));
 sky130_fd_sc_hd__and2_1 _20221_ (.A(_03718_),
    .B(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__clkbuf_1 _20222_ (.A(_03737_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _20223_ (.A0(\rbzero.pov.ready_buffer[54] ),
    .A1(\rbzero.pov.spi_buffer[54] ),
    .S(_03725_),
    .X(_03738_));
 sky130_fd_sc_hd__and2_1 _20224_ (.A(_03718_),
    .B(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__clkbuf_1 _20225_ (.A(_03739_),
    .X(_01229_));
 sky130_fd_sc_hd__clkbuf_2 _20226_ (.A(_08091_),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _20227_ (.A0(\rbzero.pov.ready_buffer[55] ),
    .A1(\rbzero.pov.spi_buffer[55] ),
    .S(_03725_),
    .X(_03741_));
 sky130_fd_sc_hd__and2_1 _20228_ (.A(_03740_),
    .B(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__clkbuf_1 _20229_ (.A(_03742_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _20230_ (.A0(\rbzero.pov.ready_buffer[56] ),
    .A1(\rbzero.pov.spi_buffer[56] ),
    .S(_03725_),
    .X(_03743_));
 sky130_fd_sc_hd__and2_1 _20231_ (.A(_03740_),
    .B(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_1 _20232_ (.A(_03744_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _20233_ (.A0(\rbzero.pov.ready_buffer[57] ),
    .A1(\rbzero.pov.spi_buffer[57] ),
    .S(_03725_),
    .X(_03745_));
 sky130_fd_sc_hd__and2_1 _20234_ (.A(_03740_),
    .B(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _20235_ (.A(_03746_),
    .X(_01232_));
 sky130_fd_sc_hd__clkbuf_4 _20236_ (.A(\rbzero.pov.spi_done ),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_1 _20237_ (.A0(\rbzero.pov.ready_buffer[58] ),
    .A1(\rbzero.pov.spi_buffer[58] ),
    .S(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__and2_1 _20238_ (.A(_03740_),
    .B(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_1 _20239_ (.A(_03749_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _20240_ (.A0(\rbzero.pov.ready_buffer[59] ),
    .A1(\rbzero.pov.spi_buffer[59] ),
    .S(_03747_),
    .X(_03750_));
 sky130_fd_sc_hd__and2_1 _20241_ (.A(_03740_),
    .B(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_1 _20242_ (.A(_03751_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _20243_ (.A0(\rbzero.pov.ready_buffer[60] ),
    .A1(\rbzero.pov.spi_buffer[60] ),
    .S(_03747_),
    .X(_03752_));
 sky130_fd_sc_hd__and2_1 _20244_ (.A(_03740_),
    .B(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__clkbuf_1 _20245_ (.A(_03753_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _20246_ (.A0(\rbzero.pov.ready_buffer[61] ),
    .A1(\rbzero.pov.spi_buffer[61] ),
    .S(_03747_),
    .X(_03754_));
 sky130_fd_sc_hd__and2_1 _20247_ (.A(_03740_),
    .B(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _20248_ (.A(_03755_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _20249_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(\rbzero.pov.spi_buffer[62] ),
    .S(_03747_),
    .X(_03756_));
 sky130_fd_sc_hd__and2_1 _20250_ (.A(_03740_),
    .B(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _20251_ (.A(_03757_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _20252_ (.A0(\rbzero.pov.ready_buffer[63] ),
    .A1(\rbzero.pov.spi_buffer[63] ),
    .S(_03747_),
    .X(_03758_));
 sky130_fd_sc_hd__and2_1 _20253_ (.A(_03740_),
    .B(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_1 _20254_ (.A(_03759_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _20255_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(\rbzero.pov.spi_buffer[64] ),
    .S(_03747_),
    .X(_03760_));
 sky130_fd_sc_hd__and2_1 _20256_ (.A(_03740_),
    .B(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _20257_ (.A(_03761_),
    .X(_01239_));
 sky130_fd_sc_hd__clkbuf_4 _20258_ (.A(_08091_),
    .X(_03762_));
 sky130_fd_sc_hd__mux2_1 _20259_ (.A0(\rbzero.pov.ready_buffer[65] ),
    .A1(\rbzero.pov.spi_buffer[65] ),
    .S(_03747_),
    .X(_03763_));
 sky130_fd_sc_hd__and2_1 _20260_ (.A(_03762_),
    .B(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _20261_ (.A(_03764_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _20262_ (.A0(\rbzero.pov.ready_buffer[66] ),
    .A1(\rbzero.pov.spi_buffer[66] ),
    .S(_03747_),
    .X(_03765_));
 sky130_fd_sc_hd__and2_1 _20263_ (.A(_03762_),
    .B(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _20264_ (.A(_03766_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _20265_ (.A0(\rbzero.pov.ready_buffer[67] ),
    .A1(\rbzero.pov.spi_buffer[67] ),
    .S(_03747_),
    .X(_03767_));
 sky130_fd_sc_hd__and2_1 _20266_ (.A(_03762_),
    .B(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_1 _20267_ (.A(_03768_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _20268_ (.A0(\rbzero.pov.ready_buffer[68] ),
    .A1(\rbzero.pov.spi_buffer[68] ),
    .S(_03636_),
    .X(_03769_));
 sky130_fd_sc_hd__and2_1 _20269_ (.A(_03762_),
    .B(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _20270_ (.A(_03770_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _20271_ (.A0(\rbzero.pov.ready_buffer[69] ),
    .A1(\rbzero.pov.spi_buffer[69] ),
    .S(_03636_),
    .X(_03771_));
 sky130_fd_sc_hd__and2_1 _20272_ (.A(_03762_),
    .B(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _20273_ (.A(_03772_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _20274_ (.A0(\rbzero.pov.ready_buffer[70] ),
    .A1(\rbzero.pov.spi_buffer[70] ),
    .S(_03636_),
    .X(_03773_));
 sky130_fd_sc_hd__and2_1 _20275_ (.A(_03762_),
    .B(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_1 _20276_ (.A(_03774_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _20277_ (.A0(\rbzero.pov.ready_buffer[71] ),
    .A1(\rbzero.pov.spi_buffer[71] ),
    .S(_03636_),
    .X(_03775_));
 sky130_fd_sc_hd__and2_1 _20278_ (.A(_03762_),
    .B(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__clkbuf_1 _20279_ (.A(_03776_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _20280_ (.A0(\rbzero.pov.ready_buffer[72] ),
    .A1(\rbzero.pov.spi_buffer[72] ),
    .S(_03636_),
    .X(_03777_));
 sky130_fd_sc_hd__and2_1 _20281_ (.A(_03762_),
    .B(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__clkbuf_1 _20282_ (.A(_03778_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _20283_ (.A0(\rbzero.pov.ready_buffer[73] ),
    .A1(\rbzero.pov.spi_buffer[73] ),
    .S(_03636_),
    .X(_03779_));
 sky130_fd_sc_hd__and2_1 _20284_ (.A(_03762_),
    .B(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_1 _20285_ (.A(_03780_),
    .X(_01248_));
 sky130_fd_sc_hd__nor3b_1 _20286_ (.A(_03498_),
    .B(_03618_),
    .C_N(_03493_),
    .Y(_01249_));
 sky130_fd_sc_hd__and2_1 _20287_ (.A(_05698_),
    .B(_09712_),
    .X(_03781_));
 sky130_fd_sc_hd__clkbuf_1 _20288_ (.A(_03781_),
    .X(_01250_));
 sky130_fd_sc_hd__and2_1 _20289_ (.A(\rbzero.pov.mosi_buffer[0] ),
    .B(_09712_),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_1 _20290_ (.A(_03782_),
    .X(_01251_));
 sky130_fd_sc_hd__and4b_1 _20291_ (.A_N(_05716_),
    .B(_05715_),
    .C(_05071_),
    .D(_05078_),
    .X(_03783_));
 sky130_fd_sc_hd__a41o_1 _20292_ (.A1(_05711_),
    .A2(_05770_),
    .A3(_04676_),
    .A4(_03783_),
    .B1(\rbzero.vga_sync.vsync ),
    .X(_03784_));
 sky130_fd_sc_hd__or4b_1 _20293_ (.A(_05770_),
    .B(_05769_),
    .C(_03369_),
    .D_N(_03783_),
    .X(_03785_));
 sky130_fd_sc_hd__and3_1 _20294_ (.A(_02653_),
    .B(_03784_),
    .C(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__clkbuf_1 _20295_ (.A(_03786_),
    .X(_01252_));
 sky130_fd_sc_hd__inv_2 _20296_ (.A(_04689_),
    .Y(_03787_));
 sky130_fd_sc_hd__and4_1 _20297_ (.A(_04454_),
    .B(_04484_),
    .C(_04019_),
    .D(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__and4_1 _20298_ (.A(_04014_),
    .B(_04481_),
    .C(_05003_),
    .D(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__a31o_1 _20299_ (.A1(_04014_),
    .A2(_05172_),
    .A3(_03788_),
    .B1(_04450_),
    .X(_03790_));
 sky130_fd_sc_hd__o21ba_1 _20300_ (.A1(\rbzero.hsync ),
    .A2(_03789_),
    .B1_N(_03790_),
    .X(_01253_));
 sky130_fd_sc_hd__or3_1 _20301_ (.A(_05770_),
    .B(_05769_),
    .C(_03369_),
    .X(_03791_));
 sky130_fd_sc_hd__or3b_1 _20302_ (.A(_05715_),
    .B(_04671_),
    .C_N(_05716_),
    .X(_03792_));
 sky130_fd_sc_hd__or4_1 _20303_ (.A(_04683_),
    .B(_04681_),
    .C(_03791_),
    .D(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__a21oi_1 _20304_ (.A1(_09709_),
    .A2(_03793_),
    .B1(_05769_),
    .Y(_03794_));
 sky130_fd_sc_hd__a211oi_1 _20305_ (.A1(_05769_),
    .A2(_09709_),
    .B1(_03794_),
    .C1(_02731_),
    .Y(_01254_));
 sky130_fd_sc_hd__a21o_1 _20306_ (.A1(_05769_),
    .A2(_09709_),
    .B1(_05770_),
    .X(_03795_));
 sky130_fd_sc_hd__and3_1 _20307_ (.A(_02653_),
    .B(_03370_),
    .C(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__clkbuf_1 _20308_ (.A(_03796_),
    .X(_01255_));
 sky130_fd_sc_hd__nand2_1 _20309_ (.A(_05062_),
    .B(_03370_),
    .Y(_03797_));
 sky130_fd_sc_hd__a21o_1 _20310_ (.A1(_08091_),
    .A2(_03793_),
    .B1(_09716_),
    .X(_03798_));
 sky130_fd_sc_hd__o211a_1 _20311_ (.A1(_05062_),
    .A2(_03370_),
    .B1(_03797_),
    .C1(_03798_),
    .X(_01256_));
 sky130_fd_sc_hd__buf_4 _20312_ (.A(_09716_),
    .X(_03799_));
 sky130_fd_sc_hd__a31o_1 _20313_ (.A1(_04675_),
    .A2(_05770_),
    .A3(_05769_),
    .B1(_05711_),
    .X(_03800_));
 sky130_fd_sc_hd__and4b_1 _20314_ (.A_N(_02679_),
    .B(_03793_),
    .C(_03800_),
    .D(_09709_),
    .X(_03801_));
 sky130_fd_sc_hd__a22o_1 _20315_ (.A1(_05711_),
    .A2(_03799_),
    .B1(_03801_),
    .B2(_02901_),
    .X(_01257_));
 sky130_fd_sc_hd__nand2_1 _20316_ (.A(_05186_),
    .B(_02680_),
    .Y(_03802_));
 sky130_fd_sc_hd__or2_1 _20317_ (.A(_05186_),
    .B(_02680_),
    .X(_03803_));
 sky130_fd_sc_hd__a21oi_1 _20318_ (.A1(_03802_),
    .A2(_03803_),
    .B1(_03353_),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _20319_ (.A(_05074_),
    .B(_02680_),
    .Y(_03804_));
 sky130_fd_sc_hd__inv_2 _20320_ (.A(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__o2111a_1 _20321_ (.A1(_05016_),
    .A2(_03802_),
    .B1(_03805_),
    .C1(_02901_),
    .D1(_04681_),
    .X(_01259_));
 sky130_fd_sc_hd__o21ai_1 _20322_ (.A1(_04683_),
    .A2(_03804_),
    .B1(_02901_),
    .Y(_03806_));
 sky130_fd_sc_hd__nor2_1 _20323_ (.A(_05014_),
    .B(_03805_),
    .Y(_03807_));
 sky130_fd_sc_hd__nor2_1 _20324_ (.A(_03806_),
    .B(_03807_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_1 _20325_ (.A(_02676_),
    .B(_03804_),
    .Y(_03808_));
 sky130_fd_sc_hd__o211a_1 _20326_ (.A1(_04671_),
    .A2(_03807_),
    .B1(_03808_),
    .C1(_02901_),
    .X(_01261_));
 sky130_fd_sc_hd__nor2_1 _20327_ (.A(_05074_),
    .B(_03371_),
    .Y(_03809_));
 sky130_fd_sc_hd__and3_1 _20328_ (.A(_05715_),
    .B(_02676_),
    .C(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__a21o_1 _20329_ (.A1(_02676_),
    .A2(_03804_),
    .B1(_05715_),
    .X(_03811_));
 sky130_fd_sc_hd__and3b_1 _20330_ (.A_N(_03810_),
    .B(_08092_),
    .C(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_1 _20331_ (.A(_03812_),
    .X(_01262_));
 sky130_fd_sc_hd__a21boi_1 _20332_ (.A1(_05716_),
    .A2(_03810_),
    .B1_N(_03798_),
    .Y(_03813_));
 sky130_fd_sc_hd__o21a_1 _20333_ (.A1(_05716_),
    .A2(_03810_),
    .B1(_03813_),
    .X(_01263_));
 sky130_fd_sc_hd__and2_1 _20334_ (.A(net46),
    .B(_09712_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_1 _20335_ (.A(_03814_),
    .X(_01264_));
 sky130_fd_sc_hd__and2_1 _20336_ (.A(\rbzero.spi_registers.sclk_buffer[0] ),
    .B(_09712_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _20337_ (.A(_03815_),
    .X(_01265_));
 sky130_fd_sc_hd__and2_1 _20338_ (.A(\rbzero.spi_registers.sclk_buffer[1] ),
    .B(_09712_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _20339_ (.A(_03816_),
    .X(_01266_));
 sky130_fd_sc_hd__inv_2 _20341__93 (.A(clknet_1_1__leaf__03617_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _20342__94 (.A(clknet_1_1__leaf__03617_),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _20343__95 (.A(clknet_1_1__leaf__03617_),
    .Y(net221));
 sky130_fd_sc_hd__inv_2 _20344__96 (.A(clknet_1_1__leaf__03617_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _20345__97 (.A(clknet_1_1__leaf__03617_),
    .Y(net223));
 sky130_fd_sc_hd__inv_2 _20347__98 (.A(clknet_1_0__leaf__03817_),
    .Y(net224));
 sky130_fd_sc_hd__buf_1 _20346_ (.A(clknet_1_0__leaf__03616_),
    .X(_03817_));
 sky130_fd_sc_hd__inv_2 _20348__99 (.A(clknet_1_0__leaf__03817_),
    .Y(net225));
 sky130_fd_sc_hd__inv_2 _20349__100 (.A(clknet_1_0__leaf__03817_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _20350__101 (.A(clknet_1_0__leaf__03817_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _20351__102 (.A(clknet_1_1__leaf__03817_),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _20352__103 (.A(clknet_1_1__leaf__03817_),
    .Y(net229));
 sky130_fd_sc_hd__inv_2 _20353__104 (.A(clknet_1_1__leaf__03817_),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _20354__105 (.A(clknet_1_1__leaf__03817_),
    .Y(net231));
 sky130_fd_sc_hd__inv_2 _20355__106 (.A(clknet_1_1__leaf__03817_),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _20356__107 (.A(clknet_1_1__leaf__03817_),
    .Y(net233));
 sky130_fd_sc_hd__inv_2 _20358__108 (.A(clknet_1_0__leaf__03818_),
    .Y(net234));
 sky130_fd_sc_hd__buf_1 _20357_ (.A(clknet_1_0__leaf__03616_),
    .X(_03818_));
 sky130_fd_sc_hd__inv_2 _20359__109 (.A(clknet_1_0__leaf__03818_),
    .Y(net235));
 sky130_fd_sc_hd__inv_2 _20360__110 (.A(clknet_1_1__leaf__03818_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _20361__111 (.A(clknet_1_1__leaf__03818_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _20362__112 (.A(clknet_1_1__leaf__03818_),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _20363__113 (.A(clknet_1_1__leaf__03818_),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _20364__114 (.A(clknet_1_1__leaf__03818_),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _20365__115 (.A(clknet_1_0__leaf__03818_),
    .Y(net241));
 sky130_fd_sc_hd__inv_2 _20366__116 (.A(clknet_1_0__leaf__03818_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _20367__117 (.A(clknet_1_0__leaf__03818_),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _20369__118 (.A(clknet_1_0__leaf__03819_),
    .Y(net244));
 sky130_fd_sc_hd__buf_1 _20368_ (.A(clknet_1_0__leaf__03616_),
    .X(_03819_));
 sky130_fd_sc_hd__inv_2 _20370__119 (.A(clknet_1_0__leaf__03819_),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _20371__120 (.A(clknet_1_0__leaf__03819_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _20372__121 (.A(clknet_1_0__leaf__03819_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _20373__122 (.A(clknet_1_0__leaf__03819_),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _20374__123 (.A(clknet_1_1__leaf__03819_),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _20375__124 (.A(clknet_1_1__leaf__03819_),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _20376__125 (.A(clknet_1_1__leaf__03819_),
    .Y(net251));
 sky130_fd_sc_hd__inv_2 _20377__126 (.A(clknet_1_1__leaf__03819_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _20378__127 (.A(clknet_1_1__leaf__03819_),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _20380__128 (.A(clknet_1_0__leaf__03820_),
    .Y(net254));
 sky130_fd_sc_hd__buf_1 _20379_ (.A(clknet_1_0__leaf__03616_),
    .X(_03820_));
 sky130_fd_sc_hd__inv_2 _20381__129 (.A(clknet_1_1__leaf__03820_),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _20382__130 (.A(clknet_1_1__leaf__03820_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _20383__131 (.A(clknet_1_1__leaf__03820_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _20384__132 (.A(clknet_1_1__leaf__03820_),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _20385__133 (.A(clknet_1_1__leaf__03820_),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _20386__134 (.A(clknet_1_0__leaf__03820_),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _20387__135 (.A(clknet_1_0__leaf__03820_),
    .Y(net261));
 sky130_fd_sc_hd__inv_2 _20388__136 (.A(clknet_1_0__leaf__03820_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _20389__137 (.A(clknet_1_0__leaf__03820_),
    .Y(net263));
 sky130_fd_sc_hd__inv_2 _20391__138 (.A(clknet_1_0__leaf__03821_),
    .Y(net264));
 sky130_fd_sc_hd__buf_1 _20390_ (.A(clknet_1_0__leaf__03616_),
    .X(_03821_));
 sky130_fd_sc_hd__inv_2 _20392__139 (.A(clknet_1_0__leaf__03821_),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _20393__140 (.A(clknet_1_0__leaf__03821_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _20394__141 (.A(clknet_1_0__leaf__03821_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _20395__142 (.A(clknet_1_1__leaf__03821_),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _20396__143 (.A(clknet_1_1__leaf__03821_),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _20397__144 (.A(clknet_1_1__leaf__03821_),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _20398__145 (.A(clknet_1_1__leaf__03821_),
    .Y(net271));
 sky130_fd_sc_hd__inv_2 _20399__146 (.A(clknet_1_1__leaf__03821_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _20400__147 (.A(clknet_1_1__leaf__03821_),
    .Y(net273));
 sky130_fd_sc_hd__inv_2 _20402__148 (.A(clknet_1_0__leaf__03822_),
    .Y(net274));
 sky130_fd_sc_hd__buf_1 _20401_ (.A(clknet_1_1__leaf__03616_),
    .X(_03822_));
 sky130_fd_sc_hd__inv_2 _20403__149 (.A(clknet_1_0__leaf__03822_),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _20404__150 (.A(clknet_1_0__leaf__03822_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _20405__151 (.A(clknet_1_0__leaf__03822_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _20406__152 (.A(clknet_1_0__leaf__03822_),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _20407__153 (.A(clknet_1_0__leaf__03822_),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _20408__154 (.A(clknet_1_1__leaf__03822_),
    .Y(net280));
 sky130_fd_sc_hd__inv_2 _20409__155 (.A(clknet_1_1__leaf__03822_),
    .Y(net281));
 sky130_fd_sc_hd__inv_2 _20410__156 (.A(clknet_1_1__leaf__03822_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _20411__157 (.A(clknet_1_1__leaf__03822_),
    .Y(net283));
 sky130_fd_sc_hd__inv_2 _20413__158 (.A(clknet_1_1__leaf__03823_),
    .Y(net284));
 sky130_fd_sc_hd__buf_1 _20412_ (.A(clknet_1_1__leaf__03616_),
    .X(_03823_));
 sky130_fd_sc_hd__inv_2 _20414__159 (.A(clknet_1_1__leaf__03823_),
    .Y(net285));
 sky130_fd_sc_hd__inv_2 _20415__160 (.A(clknet_1_1__leaf__03823_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _20416__161 (.A(clknet_1_0__leaf__03823_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _20417__162 (.A(clknet_1_0__leaf__03823_),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _20418__163 (.A(clknet_1_0__leaf__03823_),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _20419__164 (.A(clknet_1_0__leaf__03823_),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _20420__165 (.A(clknet_1_1__leaf__03823_),
    .Y(net291));
 sky130_fd_sc_hd__inv_2 _20421__166 (.A(clknet_1_1__leaf__03823_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _20422__167 (.A(clknet_1_1__leaf__03823_),
    .Y(net293));
 sky130_fd_sc_hd__inv_2 _20424__168 (.A(clknet_1_0__leaf__03824_),
    .Y(net294));
 sky130_fd_sc_hd__buf_1 _20423_ (.A(clknet_1_1__leaf__03616_),
    .X(_03824_));
 sky130_fd_sc_hd__inv_2 _20425__169 (.A(clknet_1_0__leaf__03824_),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _20426__170 (.A(clknet_1_0__leaf__03824_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _20427__171 (.A(clknet_1_0__leaf__03824_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _20428__172 (.A(clknet_1_0__leaf__03824_),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _20429__173 (.A(clknet_1_0__leaf__03824_),
    .Y(net299));
 sky130_fd_sc_hd__inv_2 _20430__174 (.A(clknet_1_1__leaf__03824_),
    .Y(net300));
 sky130_fd_sc_hd__inv_2 _20431__175 (.A(clknet_1_1__leaf__03824_),
    .Y(net301));
 sky130_fd_sc_hd__inv_2 _20432__176 (.A(clknet_1_1__leaf__03824_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _20433__177 (.A(clknet_1_1__leaf__03824_),
    .Y(net303));
 sky130_fd_sc_hd__inv_2 _20435__178 (.A(clknet_1_1__leaf__03825_),
    .Y(net304));
 sky130_fd_sc_hd__buf_1 _20434_ (.A(clknet_1_1__leaf__03616_),
    .X(_03825_));
 sky130_fd_sc_hd__inv_2 _20436__179 (.A(clknet_1_1__leaf__03825_),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _20437__180 (.A(clknet_1_1__leaf__03825_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _20438__181 (.A(clknet_1_0__leaf__03825_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _20439__182 (.A(clknet_1_0__leaf__03825_),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _20440__183 (.A(clknet_1_0__leaf__03825_),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _20441__184 (.A(clknet_1_0__leaf__03825_),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 _20442__185 (.A(clknet_1_0__leaf__03825_),
    .Y(net311));
 sky130_fd_sc_hd__inv_2 _20443__186 (.A(clknet_1_1__leaf__03825_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _20444__187 (.A(clknet_1_1__leaf__03825_),
    .Y(net313));
 sky130_fd_sc_hd__inv_2 _20447__188 (.A(clknet_1_1__leaf__03827_),
    .Y(net314));
 sky130_fd_sc_hd__buf_1 _20445_ (.A(clknet_1_1__leaf__05762_),
    .X(_03826_));
 sky130_fd_sc_hd__buf_1 _20446_ (.A(clknet_1_1__leaf__03826_),
    .X(_03827_));
 sky130_fd_sc_hd__inv_2 _20448__189 (.A(clknet_1_1__leaf__03827_),
    .Y(net315));
 sky130_fd_sc_hd__inv_2 _20449__190 (.A(clknet_1_0__leaf__03827_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _20450__191 (.A(clknet_1_0__leaf__03827_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _20451__192 (.A(clknet_1_0__leaf__03827_),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _20452__193 (.A(clknet_1_0__leaf__03827_),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 _20453__194 (.A(clknet_1_0__leaf__03827_),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _20454__195 (.A(clknet_1_0__leaf__03827_),
    .Y(net321));
 sky130_fd_sc_hd__inv_2 _20455__196 (.A(clknet_1_1__leaf__03827_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _20456__197 (.A(clknet_1_1__leaf__03827_),
    .Y(net323));
 sky130_fd_sc_hd__inv_2 _20458__198 (.A(clknet_1_0__leaf__03828_),
    .Y(net324));
 sky130_fd_sc_hd__buf_1 _20457_ (.A(clknet_1_0__leaf__03826_),
    .X(_03828_));
 sky130_fd_sc_hd__inv_2 _20459__199 (.A(clknet_1_0__leaf__03828_),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _20460__200 (.A(clknet_1_1__leaf__03828_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _20461__201 (.A(clknet_1_1__leaf__03828_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _20462__202 (.A(clknet_1_1__leaf__03828_),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _20463__203 (.A(clknet_1_1__leaf__03828_),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _20464__204 (.A(clknet_1_1__leaf__03828_),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _20465__205 (.A(clknet_1_0__leaf__03828_),
    .Y(net331));
 sky130_fd_sc_hd__inv_2 _20466__206 (.A(clknet_1_0__leaf__03828_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _20467__207 (.A(clknet_1_0__leaf__03828_),
    .Y(net333));
 sky130_fd_sc_hd__inv_2 _20469__208 (.A(clknet_1_1__leaf__03829_),
    .Y(net334));
 sky130_fd_sc_hd__buf_1 _20468_ (.A(clknet_1_0__leaf__03826_),
    .X(_03829_));
 sky130_fd_sc_hd__inv_2 _20470__209 (.A(clknet_1_1__leaf__03829_),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _20471__210 (.A(clknet_1_1__leaf__03829_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _20472__211 (.A(clknet_1_1__leaf__03829_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _20473__212 (.A(clknet_1_1__leaf__03829_),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _20474__213 (.A(clknet_1_1__leaf__03829_),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _20475__214 (.A(clknet_1_0__leaf__03829_),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _20476__215 (.A(clknet_1_0__leaf__03829_),
    .Y(net341));
 sky130_fd_sc_hd__inv_2 _20477__216 (.A(clknet_1_0__leaf__03829_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _20478__217 (.A(clknet_1_0__leaf__03829_),
    .Y(net343));
 sky130_fd_sc_hd__inv_2 _20480__218 (.A(clknet_1_0__leaf__03830_),
    .Y(net344));
 sky130_fd_sc_hd__buf_1 _20479_ (.A(clknet_1_1__leaf__03826_),
    .X(_03830_));
 sky130_fd_sc_hd__inv_2 _20481__219 (.A(clknet_1_0__leaf__03830_),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _20482__220 (.A(clknet_1_1__leaf__03830_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _20483__221 (.A(clknet_1_1__leaf__03830_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _20484__222 (.A(clknet_1_1__leaf__03830_),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _20485__223 (.A(clknet_1_0__leaf__03830_),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _20486__224 (.A(clknet_1_0__leaf__03830_),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _20487__225 (.A(clknet_1_0__leaf__03830_),
    .Y(net351));
 sky130_fd_sc_hd__inv_2 _20488__226 (.A(clknet_1_0__leaf__03830_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _20489__227 (.A(clknet_1_1__leaf__03830_),
    .Y(net353));
 sky130_fd_sc_hd__inv_2 _20491__228 (.A(clknet_1_0__leaf__03831_),
    .Y(net354));
 sky130_fd_sc_hd__buf_1 _20490_ (.A(clknet_1_1__leaf__03826_),
    .X(_03831_));
 sky130_fd_sc_hd__inv_2 _20492__229 (.A(clknet_1_0__leaf__03831_),
    .Y(net355));
 sky130_fd_sc_hd__inv_2 _20493__230 (.A(clknet_1_1__leaf__03831_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _20494__231 (.A(clknet_1_1__leaf__03831_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _20495__232 (.A(clknet_1_1__leaf__03831_),
    .Y(net358));
 sky130_fd_sc_hd__inv_2 _20496__233 (.A(clknet_1_1__leaf__03831_),
    .Y(net359));
 sky130_fd_sc_hd__inv_2 _20497__234 (.A(clknet_1_1__leaf__03831_),
    .Y(net360));
 sky130_fd_sc_hd__inv_2 _20498__235 (.A(clknet_1_1__leaf__03831_),
    .Y(net361));
 sky130_fd_sc_hd__inv_2 _20499__236 (.A(clknet_1_0__leaf__03831_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _20500__237 (.A(clknet_1_0__leaf__03831_),
    .Y(net363));
 sky130_fd_sc_hd__inv_2 _20502__238 (.A(clknet_1_1__leaf__03832_),
    .Y(net364));
 sky130_fd_sc_hd__buf_1 _20501_ (.A(clknet_1_1__leaf__03826_),
    .X(_03832_));
 sky130_fd_sc_hd__inv_2 _20503__239 (.A(clknet_1_0__leaf__03832_),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _20504__240 (.A(clknet_1_0__leaf__03832_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _20505__241 (.A(clknet_1_1__leaf__03832_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _20506__242 (.A(clknet_1_1__leaf__03832_),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _20507__243 (.A(clknet_1_1__leaf__03832_),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _20508__244 (.A(clknet_1_1__leaf__03832_),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _20509__245 (.A(clknet_1_1__leaf__03832_),
    .Y(net371));
 sky130_fd_sc_hd__inv_2 _20510__246 (.A(clknet_1_0__leaf__03832_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _20511__247 (.A(clknet_1_0__leaf__03832_),
    .Y(net373));
 sky130_fd_sc_hd__inv_2 _20513__248 (.A(clknet_1_0__leaf__03833_),
    .Y(net374));
 sky130_fd_sc_hd__buf_1 _20512_ (.A(clknet_1_1__leaf__03826_),
    .X(_03833_));
 sky130_fd_sc_hd__inv_2 _20514__249 (.A(clknet_1_1__leaf__03833_),
    .Y(net375));
 sky130_fd_sc_hd__inv_2 _20515__250 (.A(clknet_1_1__leaf__03833_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _20516__251 (.A(clknet_1_1__leaf__03833_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _20517__252 (.A(clknet_1_0__leaf__03833_),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _20518__253 (.A(clknet_1_0__leaf__03833_),
    .Y(net379));
 sky130_fd_sc_hd__inv_2 _20519__254 (.A(clknet_1_0__leaf__03833_),
    .Y(net380));
 sky130_fd_sc_hd__inv_2 _20520__255 (.A(clknet_1_1__leaf__03833_),
    .Y(net381));
 sky130_fd_sc_hd__inv_2 _20521__256 (.A(clknet_1_1__leaf__03833_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _20522__257 (.A(clknet_1_0__leaf__03833_),
    .Y(net383));
 sky130_fd_sc_hd__inv_2 _20524__258 (.A(clknet_1_1__leaf__03834_),
    .Y(net384));
 sky130_fd_sc_hd__buf_1 _20523_ (.A(clknet_1_1__leaf__03826_),
    .X(_03834_));
 sky130_fd_sc_hd__inv_2 _20525__259 (.A(clknet_1_1__leaf__03834_),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _20526__260 (.A(clknet_1_0__leaf__03834_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _20527__261 (.A(clknet_1_0__leaf__03834_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _20528__262 (.A(clknet_1_0__leaf__03834_),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _20529__263 (.A(clknet_1_0__leaf__03834_),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _20530__264 (.A(clknet_1_0__leaf__03834_),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _20531__265 (.A(clknet_1_0__leaf__03834_),
    .Y(net391));
 sky130_fd_sc_hd__inv_2 _20532__266 (.A(clknet_1_1__leaf__03834_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _20533__267 (.A(clknet_1_1__leaf__03834_),
    .Y(net393));
 sky130_fd_sc_hd__inv_2 _20535__268 (.A(clknet_1_1__leaf__03835_),
    .Y(net394));
 sky130_fd_sc_hd__buf_1 _20534_ (.A(clknet_1_0__leaf__03826_),
    .X(_03835_));
 sky130_fd_sc_hd__inv_2 _20536__269 (.A(clknet_1_1__leaf__03835_),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _20537__270 (.A(clknet_1_0__leaf__03835_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _20538__271 (.A(clknet_1_0__leaf__03835_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _20539__272 (.A(clknet_1_0__leaf__03835_),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _20540__273 (.A(clknet_1_1__leaf__03835_),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _20541__274 (.A(clknet_1_1__leaf__03835_),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _20542__275 (.A(clknet_1_0__leaf__03835_),
    .Y(net401));
 sky130_fd_sc_hd__inv_2 _20543__276 (.A(clknet_1_0__leaf__03835_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _20544__277 (.A(clknet_1_0__leaf__03835_),
    .Y(net403));
 sky130_fd_sc_hd__inv_2 _20546__278 (.A(clknet_1_1__leaf__03836_),
    .Y(net404));
 sky130_fd_sc_hd__buf_1 _20545_ (.A(clknet_1_0__leaf__03826_),
    .X(_03836_));
 sky130_fd_sc_hd__inv_2 _20547__279 (.A(clknet_1_1__leaf__03836_),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _20548__280 (.A(clknet_1_1__leaf__03836_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _20549__281 (.A(clknet_1_1__leaf__03836_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _20550__282 (.A(clknet_1_0__leaf__03836_),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _20551__283 (.A(clknet_1_1__leaf__03836_),
    .Y(net409));
 sky130_fd_sc_hd__inv_2 _20552__284 (.A(clknet_1_0__leaf__03836_),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _20553__285 (.A(clknet_1_0__leaf__03836_),
    .Y(net411));
 sky130_fd_sc_hd__inv_2 _20554__286 (.A(clknet_1_0__leaf__03836_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _20555__287 (.A(clknet_1_0__leaf__03836_),
    .Y(net413));
 sky130_fd_sc_hd__inv_2 _20558__288 (.A(clknet_1_1__leaf__03838_),
    .Y(net414));
 sky130_fd_sc_hd__buf_1 _20556_ (.A(clknet_1_0__leaf__05762_),
    .X(_03837_));
 sky130_fd_sc_hd__buf_1 _20557_ (.A(clknet_1_0__leaf__03837_),
    .X(_03838_));
 sky130_fd_sc_hd__inv_2 _20559__289 (.A(clknet_1_0__leaf__03838_),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _20560__290 (.A(clknet_1_0__leaf__03838_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _20561__291 (.A(clknet_1_0__leaf__03838_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _20562__292 (.A(clknet_1_1__leaf__03838_),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _20563__293 (.A(clknet_1_1__leaf__03838_),
    .Y(net419));
 sky130_fd_sc_hd__inv_2 _20564__294 (.A(clknet_1_1__leaf__03838_),
    .Y(net420));
 sky130_fd_sc_hd__inv_2 _20565__295 (.A(clknet_1_0__leaf__03838_),
    .Y(net421));
 sky130_fd_sc_hd__inv_2 _20566__296 (.A(clknet_1_0__leaf__03838_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _20567__297 (.A(clknet_1_0__leaf__03838_),
    .Y(net423));
 sky130_fd_sc_hd__inv_2 _20569__298 (.A(clknet_1_0__leaf__03839_),
    .Y(net424));
 sky130_fd_sc_hd__buf_1 _20568_ (.A(clknet_1_0__leaf__03837_),
    .X(_03839_));
 sky130_fd_sc_hd__inv_2 _20570__299 (.A(clknet_1_0__leaf__03839_),
    .Y(net425));
 sky130_fd_sc_hd__inv_2 _20571__300 (.A(clknet_1_1__leaf__03839_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _20572__301 (.A(clknet_1_1__leaf__03839_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _20573__302 (.A(clknet_1_1__leaf__03839_),
    .Y(net428));
 sky130_fd_sc_hd__inv_2 _20574__303 (.A(clknet_1_1__leaf__03839_),
    .Y(net429));
 sky130_fd_sc_hd__inv_2 _20575__304 (.A(clknet_1_0__leaf__03839_),
    .Y(net430));
 sky130_fd_sc_hd__inv_2 _20576__305 (.A(clknet_1_0__leaf__03839_),
    .Y(net431));
 sky130_fd_sc_hd__inv_2 _20577__306 (.A(clknet_1_0__leaf__03839_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _20578__307 (.A(clknet_1_0__leaf__03839_),
    .Y(net433));
 sky130_fd_sc_hd__inv_2 _20580__308 (.A(clknet_1_0__leaf__03840_),
    .Y(net434));
 sky130_fd_sc_hd__buf_1 _20579_ (.A(clknet_1_0__leaf__03837_),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _20581__309 (.A(clknet_1_0__leaf__03840_),
    .Y(net435));
 sky130_fd_sc_hd__inv_2 _20582__310 (.A(clknet_1_0__leaf__03840_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _20583__311 (.A(clknet_1_0__leaf__03840_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _20584__312 (.A(clknet_1_0__leaf__03840_),
    .Y(net438));
 sky130_fd_sc_hd__inv_2 _20585__313 (.A(clknet_1_1__leaf__03840_),
    .Y(net439));
 sky130_fd_sc_hd__inv_2 _20586__314 (.A(clknet_1_1__leaf__03840_),
    .Y(net440));
 sky130_fd_sc_hd__inv_2 _20587__315 (.A(clknet_1_1__leaf__03840_),
    .Y(net441));
 sky130_fd_sc_hd__inv_2 _20588__316 (.A(clknet_1_1__leaf__03840_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _20589__317 (.A(clknet_1_1__leaf__03840_),
    .Y(net443));
 sky130_fd_sc_hd__inv_2 _20591__318 (.A(clknet_1_0__leaf__03841_),
    .Y(net444));
 sky130_fd_sc_hd__buf_1 _20590_ (.A(clknet_1_0__leaf__03837_),
    .X(_03841_));
 sky130_fd_sc_hd__inv_2 _20592__319 (.A(clknet_1_0__leaf__03841_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _20593__320 (.A(clknet_1_0__leaf__03841_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _20594__321 (.A(clknet_1_1__leaf__03841_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _20595__322 (.A(clknet_1_0__leaf__03841_),
    .Y(net448));
 sky130_fd_sc_hd__inv_2 _20596__323 (.A(clknet_1_1__leaf__03841_),
    .Y(net449));
 sky130_fd_sc_hd__inv_2 _20597__324 (.A(clknet_1_1__leaf__03841_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _20598__325 (.A(clknet_1_1__leaf__03841_),
    .Y(net451));
 sky130_fd_sc_hd__inv_2 _20599__326 (.A(clknet_1_1__leaf__03841_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _20600__327 (.A(clknet_1_1__leaf__03841_),
    .Y(net453));
 sky130_fd_sc_hd__inv_2 _20602__328 (.A(clknet_1_1__leaf__03842_),
    .Y(net454));
 sky130_fd_sc_hd__buf_1 _20601_ (.A(clknet_1_0__leaf__03837_),
    .X(_03842_));
 sky130_fd_sc_hd__inv_2 _20603__329 (.A(clknet_1_1__leaf__03842_),
    .Y(net455));
 sky130_fd_sc_hd__inv_2 _20604__330 (.A(clknet_1_1__leaf__03842_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _20605__331 (.A(clknet_1_1__leaf__03842_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _20606__332 (.A(clknet_1_0__leaf__03842_),
    .Y(net458));
 sky130_fd_sc_hd__inv_2 _20607__333 (.A(clknet_1_0__leaf__03842_),
    .Y(net459));
 sky130_fd_sc_hd__inv_2 _20608__334 (.A(clknet_1_0__leaf__03842_),
    .Y(net460));
 sky130_fd_sc_hd__inv_2 _20609__335 (.A(clknet_1_0__leaf__03842_),
    .Y(net461));
 sky130_fd_sc_hd__inv_2 _20610__336 (.A(clknet_1_0__leaf__03842_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _20611__337 (.A(clknet_1_0__leaf__03842_),
    .Y(net463));
 sky130_fd_sc_hd__inv_2 _20613__338 (.A(clknet_1_1__leaf__03843_),
    .Y(net464));
 sky130_fd_sc_hd__buf_1 _20612_ (.A(clknet_1_0__leaf__03837_),
    .X(_03843_));
 sky130_fd_sc_hd__inv_2 _20614__339 (.A(clknet_1_1__leaf__03843_),
    .Y(net465));
 sky130_fd_sc_hd__inv_2 _20615__340 (.A(clknet_1_1__leaf__03843_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _20616__341 (.A(clknet_1_1__leaf__03843_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _20617__342 (.A(clknet_1_0__leaf__03843_),
    .Y(net468));
 sky130_fd_sc_hd__inv_2 _20618__343 (.A(clknet_1_0__leaf__03843_),
    .Y(net469));
 sky130_fd_sc_hd__inv_2 _20619__344 (.A(clknet_1_0__leaf__03843_),
    .Y(net470));
 sky130_fd_sc_hd__inv_2 _20620__345 (.A(clknet_1_0__leaf__03843_),
    .Y(net471));
 sky130_fd_sc_hd__inv_2 _20621__346 (.A(clknet_1_0__leaf__03843_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _20622__347 (.A(clknet_1_0__leaf__03843_),
    .Y(net473));
 sky130_fd_sc_hd__inv_2 _20624__348 (.A(clknet_1_0__leaf__03844_),
    .Y(net474));
 sky130_fd_sc_hd__buf_1 _20623_ (.A(clknet_1_1__leaf__03837_),
    .X(_03844_));
 sky130_fd_sc_hd__inv_2 _20625__349 (.A(clknet_1_0__leaf__03844_),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _20626__350 (.A(clknet_1_0__leaf__03844_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _20627__351 (.A(clknet_1_0__leaf__03844_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _20628__352 (.A(clknet_1_0__leaf__03844_),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _20629__353 (.A(clknet_1_0__leaf__03844_),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _20630__354 (.A(clknet_1_1__leaf__03844_),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _20631__355 (.A(clknet_1_1__leaf__03844_),
    .Y(net481));
 sky130_fd_sc_hd__inv_2 _20632__356 (.A(clknet_1_1__leaf__03844_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _20633__357 (.A(clknet_1_1__leaf__03844_),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _20635__358 (.A(clknet_1_0__leaf__03845_),
    .Y(net484));
 sky130_fd_sc_hd__buf_1 _20634_ (.A(clknet_1_1__leaf__03837_),
    .X(_03845_));
 sky130_fd_sc_hd__inv_2 _20636__359 (.A(clknet_1_1__leaf__03845_),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _20637__360 (.A(clknet_1_1__leaf__03845_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _20638__361 (.A(clknet_1_1__leaf__03845_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _20639__362 (.A(clknet_1_1__leaf__03845_),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _20640__363 (.A(clknet_1_1__leaf__03845_),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _20641__364 (.A(clknet_1_0__leaf__03845_),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _20642__365 (.A(clknet_1_0__leaf__03845_),
    .Y(net491));
 sky130_fd_sc_hd__inv_2 _20643__366 (.A(clknet_1_0__leaf__03845_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _20644__367 (.A(clknet_1_0__leaf__03845_),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _20646__368 (.A(clknet_1_0__leaf__03846_),
    .Y(net494));
 sky130_fd_sc_hd__buf_1 _20645_ (.A(clknet_1_1__leaf__03837_),
    .X(_03846_));
 sky130_fd_sc_hd__inv_2 _20647__369 (.A(clknet_1_0__leaf__03846_),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _20648__370 (.A(clknet_1_1__leaf__03846_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _20649__371 (.A(clknet_1_1__leaf__03846_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _20650__372 (.A(clknet_1_1__leaf__03846_),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _20651__373 (.A(clknet_1_1__leaf__03846_),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _20652__374 (.A(clknet_1_1__leaf__03846_),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _20653__375 (.A(clknet_1_0__leaf__03846_),
    .Y(net501));
 sky130_fd_sc_hd__inv_2 _20654__376 (.A(clknet_1_0__leaf__03846_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _20655__377 (.A(clknet_1_0__leaf__03846_),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _20657__378 (.A(clknet_1_1__leaf__03847_),
    .Y(net504));
 sky130_fd_sc_hd__buf_1 _20656_ (.A(clknet_1_1__leaf__03837_),
    .X(_03847_));
 sky130_fd_sc_hd__inv_2 _20658__379 (.A(clknet_1_1__leaf__03847_),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _20659__380 (.A(clknet_1_1__leaf__03847_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _20660__381 (.A(clknet_1_1__leaf__03847_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _20661__382 (.A(clknet_1_1__leaf__03847_),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _20662__383 (.A(clknet_1_0__leaf__03847_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _20663__384 (.A(clknet_1_0__leaf__03847_),
    .Y(net510));
 sky130_fd_sc_hd__inv_2 _20664__385 (.A(clknet_1_0__leaf__03847_),
    .Y(net511));
 sky130_fd_sc_hd__inv_2 _20665__386 (.A(clknet_1_0__leaf__03847_),
    .Y(net512));
 sky130_fd_sc_hd__inv_2 _20666__387 (.A(clknet_1_0__leaf__03847_),
    .Y(net513));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__buf_1 _20667_ (.A(clknet_1_1__leaf__05762_),
    .X(_03848_));
 sky130_fd_sc_hd__inv_2 _20669__9 (.A(clknet_1_1__leaf__03848_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _20670__10 (.A(clknet_1_0__leaf__03848_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _20671__11 (.A(clknet_1_0__leaf__03848_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _20672__12 (.A(clknet_1_0__leaf__03848_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _20673__13 (.A(clknet_1_0__leaf__03848_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _20674__14 (.A(clknet_1_0__leaf__03848_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _20675__15 (.A(clknet_1_1__leaf__03848_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _20676__16 (.A(clknet_1_1__leaf__03848_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _20677__17 (.A(clknet_1_1__leaf__03848_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _20679__18 (.A(clknet_1_1__leaf__03849_),
    .Y(net144));
 sky130_fd_sc_hd__buf_1 _20678_ (.A(clknet_1_1__leaf__05762_),
    .X(_03849_));
 sky130_fd_sc_hd__inv_2 _20680__19 (.A(clknet_1_1__leaf__03849_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _20681__20 (.A(clknet_1_1__leaf__03849_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _20682__21 (.A(clknet_1_1__leaf__03849_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _20683__22 (.A(clknet_1_0__leaf__03849_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _20684__23 (.A(clknet_1_0__leaf__03849_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _20685__24 (.A(clknet_1_0__leaf__03849_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _20686__25 (.A(clknet_1_0__leaf__03849_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _20687__26 (.A(clknet_1_0__leaf__03849_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _20688__27 (.A(clknet_1_0__leaf__03849_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _19977__28 (.A(clknet_1_0__leaf__03610_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _20690__5 (.A(clknet_1_1__leaf__03609_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _20691__6 (.A(clknet_1_1__leaf__03609_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _20692__7 (.A(clknet_1_1__leaf__03609_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _20668__8 (.A(clknet_1_1__leaf__03848_),
    .Y(net134));
 sky130_fd_sc_hd__nor2_1 _20693_ (.A(\gpout5.clk_div[0] ),
    .B(net65),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _20694_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .Y(_03850_));
 sky130_fd_sc_hd__or2_1 _20695_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .X(_03851_));
 sky130_fd_sc_hd__and3_1 _20696_ (.A(_02653_),
    .B(_03850_),
    .C(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__clkbuf_1 _20697_ (.A(_03852_),
    .X(_01588_));
 sky130_fd_sc_hd__clkbuf_4 _20698_ (.A(_09716_),
    .X(_03853_));
 sky130_fd_sc_hd__nand2_1 _20699_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .Y(_03854_));
 sky130_fd_sc_hd__or2_1 _20700_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_4 _20701_ (.A(_04094_),
    .X(_03856_));
 sky130_fd_sc_hd__a32o_1 _20702_ (.A1(_03853_),
    .A2(_03854_),
    .A3(_03855_),
    .B1(_03856_),
    .B2(\rbzero.texV[-11] ),
    .X(_01589_));
 sky130_fd_sc_hd__or2_1 _20703_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .X(_03857_));
 sky130_fd_sc_hd__nand2_1 _20704_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03858_));
 sky130_fd_sc_hd__nand3b_1 _20705_ (.A_N(_03854_),
    .B(_03857_),
    .C(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__a21bo_1 _20706_ (.A1(_03857_),
    .A2(_03858_),
    .B1_N(_03854_),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_4 _20707_ (.A(_04094_),
    .X(_03861_));
 sky130_fd_sc_hd__a32o_1 _20708_ (.A1(_03853_),
    .A2(_03859_),
    .A3(_03860_),
    .B1(_03861_),
    .B2(\rbzero.texV[-10] ),
    .X(_01590_));
 sky130_fd_sc_hd__and2_1 _20709_ (.A(_03858_),
    .B(_03859_),
    .X(_03862_));
 sky130_fd_sc_hd__nor2_1 _20710_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03863_));
 sky130_fd_sc_hd__nand2_1 _20711_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03864_));
 sky130_fd_sc_hd__or2b_1 _20712_ (.A(_03863_),
    .B_N(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__xor2_1 _20713_ (.A(_03862_),
    .B(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__a22o_1 _20714_ (.A1(\rbzero.texV[-9] ),
    .A2(_03466_),
    .B1(_03799_),
    .B2(_03866_),
    .X(_01591_));
 sky130_fd_sc_hd__nor2_1 _20715_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _20716_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_03868_));
 sky130_fd_sc_hd__or2b_1 _20717_ (.A(_03867_),
    .B_N(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__o21a_1 _20718_ (.A1(_03862_),
    .A2(_03863_),
    .B1(_03864_),
    .X(_03870_));
 sky130_fd_sc_hd__or2_1 _20719_ (.A(_03869_),
    .B(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__a21oi_1 _20720_ (.A1(_03869_),
    .A2(_03870_),
    .B1(_09711_),
    .Y(_03872_));
 sky130_fd_sc_hd__a22o_1 _20721_ (.A1(\rbzero.texV[-8] ),
    .A2(_03856_),
    .B1(_03871_),
    .B2(_03872_),
    .X(_01592_));
 sky130_fd_sc_hd__nor2_1 _20722_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .Y(_03873_));
 sky130_fd_sc_hd__and2_1 _20723_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .X(_03874_));
 sky130_fd_sc_hd__o21a_1 _20724_ (.A1(_03867_),
    .A2(_03870_),
    .B1(_03868_),
    .X(_03875_));
 sky130_fd_sc_hd__o21ai_1 _20725_ (.A1(_03873_),
    .A2(_03874_),
    .B1(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__or3_1 _20726_ (.A(_03873_),
    .B(_03874_),
    .C(_03875_),
    .X(_03877_));
 sky130_fd_sc_hd__a32o_1 _20727_ (.A1(_03853_),
    .A2(_03876_),
    .A3(_03877_),
    .B1(_03861_),
    .B2(\rbzero.texV[-7] ),
    .X(_01593_));
 sky130_fd_sc_hd__xnor2_1 _20728_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_03878_));
 sky130_fd_sc_hd__o21bai_1 _20729_ (.A1(_03873_),
    .A2(_03875_),
    .B1_N(_03874_),
    .Y(_03879_));
 sky130_fd_sc_hd__xnor2_1 _20730_ (.A(_03878_),
    .B(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__a22o_1 _20731_ (.A1(\rbzero.texV[-6] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03880_),
    .X(_01594_));
 sky130_fd_sc_hd__nor2_1 _20732_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_03881_));
 sky130_fd_sc_hd__and2_1 _20733_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .X(_03882_));
 sky130_fd_sc_hd__a21o_1 _20734_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_03879_),
    .X(_03883_));
 sky130_fd_sc_hd__o21ai_1 _20735_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__or3_1 _20736_ (.A(_03881_),
    .B(_03882_),
    .C(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__o21ai_1 _20737_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03884_),
    .Y(_03886_));
 sky130_fd_sc_hd__a32o_1 _20738_ (.A1(_03853_),
    .A2(_03885_),
    .A3(_03886_),
    .B1(_03861_),
    .B2(\rbzero.texV[-5] ),
    .X(_01595_));
 sky130_fd_sc_hd__xnor2_1 _20739_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_03887_));
 sky130_fd_sc_hd__o21bai_1 _20740_ (.A1(_03881_),
    .A2(_03884_),
    .B1_N(_03882_),
    .Y(_03888_));
 sky130_fd_sc_hd__xnor2_1 _20741_ (.A(_03887_),
    .B(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__a22o_1 _20742_ (.A1(\rbzero.texV[-4] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03889_),
    .X(_01596_));
 sky130_fd_sc_hd__nor2_1 _20743_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _20744_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03891_));
 sky130_fd_sc_hd__and2b_1 _20745_ (.A_N(_03890_),
    .B(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__a21o_1 _20746_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_03888_),
    .X(_03893_));
 sky130_fd_sc_hd__o21ai_1 _20747_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(\rbzero.texV[-4] ),
    .B1(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__xnor2_1 _20748_ (.A(_03892_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__a22o_1 _20749_ (.A1(\rbzero.texV[-3] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03895_),
    .X(_01597_));
 sky130_fd_sc_hd__or2_1 _20750_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .X(_03896_));
 sky130_fd_sc_hd__nand2_1 _20751_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .Y(_03897_));
 sky130_fd_sc_hd__o21ai_1 _20752_ (.A1(_03890_),
    .A2(_03894_),
    .B1(_03891_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand3_1 _20753_ (.A(_03896_),
    .B(_03897_),
    .C(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__a21o_1 _20754_ (.A1(_03896_),
    .A2(_03897_),
    .B1(_03898_),
    .X(_03900_));
 sky130_fd_sc_hd__a32o_1 _20755_ (.A1(_03853_),
    .A2(_03899_),
    .A3(_03900_),
    .B1(_03861_),
    .B2(\rbzero.texV[-2] ),
    .X(_01598_));
 sky130_fd_sc_hd__nor2_1 _20756_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .Y(_03901_));
 sky130_fd_sc_hd__and2_1 _20757_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .X(_03902_));
 sky130_fd_sc_hd__or2_1 _20758_ (.A(_03901_),
    .B(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__a21boi_1 _20759_ (.A1(_03896_),
    .A2(_03898_),
    .B1_N(_03897_),
    .Y(_03904_));
 sky130_fd_sc_hd__xor2_1 _20760_ (.A(_03903_),
    .B(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__a22o_1 _20761_ (.A1(\rbzero.texV[-1] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03905_),
    .X(_01599_));
 sky130_fd_sc_hd__nor2_1 _20762_ (.A(_03903_),
    .B(_03904_),
    .Y(_03906_));
 sky130_fd_sc_hd__or2_1 _20763_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .X(_03907_));
 sky130_fd_sc_hd__nand2_1 _20764_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .Y(_03908_));
 sky130_fd_sc_hd__o211a_1 _20765_ (.A1(_03902_),
    .A2(_03906_),
    .B1(_03907_),
    .C1(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__inv_2 _20766_ (.A(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__a211o_1 _20767_ (.A1(_03907_),
    .A2(_03908_),
    .B1(_03902_),
    .C1(_03906_),
    .X(_03911_));
 sky130_fd_sc_hd__a32o_1 _20768_ (.A1(_03853_),
    .A2(_03910_),
    .A3(_03911_),
    .B1(_03861_),
    .B2(\rbzero.texV[0] ),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _20769_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .X(_03912_));
 sky130_fd_sc_hd__nand2_1 _20770_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .Y(_03913_));
 sky130_fd_sc_hd__nand2_1 _20771_ (.A(_03908_),
    .B(_03910_),
    .Y(_03914_));
 sky130_fd_sc_hd__and3_1 _20772_ (.A(_03912_),
    .B(_03913_),
    .C(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__inv_2 _20773_ (.A(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__a21o_1 _20774_ (.A1(_03912_),
    .A2(_03913_),
    .B1(_03914_),
    .X(_03917_));
 sky130_fd_sc_hd__a32o_1 _20775_ (.A1(_03853_),
    .A2(_03916_),
    .A3(_03917_),
    .B1(_03861_),
    .B2(\rbzero.texV[1] ),
    .X(_01601_));
 sky130_fd_sc_hd__or2_1 _20776_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .X(_03918_));
 sky130_fd_sc_hd__nand2_1 _20777_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _20778_ (.A(_03913_),
    .B(_03916_),
    .Y(_03920_));
 sky130_fd_sc_hd__and3_1 _20779_ (.A(_03918_),
    .B(_03919_),
    .C(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__inv_2 _20780_ (.A(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__a21o_1 _20781_ (.A1(_03918_),
    .A2(_03919_),
    .B1(_03920_),
    .X(_03923_));
 sky130_fd_sc_hd__a32o_1 _20782_ (.A1(_03853_),
    .A2(_03922_),
    .A3(_03923_),
    .B1(_03861_),
    .B2(\rbzero.texV[2] ),
    .X(_01602_));
 sky130_fd_sc_hd__or2_1 _20783_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .X(_03924_));
 sky130_fd_sc_hd__nand2_1 _20784_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _20785_ (.A(_03919_),
    .B(_03922_),
    .Y(_03926_));
 sky130_fd_sc_hd__a21o_1 _20786_ (.A1(_03924_),
    .A2(_03925_),
    .B1(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__and3_1 _20787_ (.A(_03924_),
    .B(_03925_),
    .C(_03926_),
    .X(_03928_));
 sky130_fd_sc_hd__inv_2 _20788_ (.A(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__a32o_1 _20789_ (.A1(_03853_),
    .A2(_03927_),
    .A3(_03929_),
    .B1(_03861_),
    .B2(\rbzero.texV[3] ),
    .X(_01603_));
 sky130_fd_sc_hd__or2_1 _20790_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_1 _20791_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _20792_ (.A(_03925_),
    .B(_03929_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand3_1 _20793_ (.A(_03930_),
    .B(_03931_),
    .C(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__a21o_1 _20794_ (.A1(_03930_),
    .A2(_03931_),
    .B1(_03932_),
    .X(_03934_));
 sky130_fd_sc_hd__a32o_1 _20795_ (.A1(_03853_),
    .A2(_03933_),
    .A3(_03934_),
    .B1(_03861_),
    .B2(\rbzero.texV[4] ),
    .X(_01604_));
 sky130_fd_sc_hd__a21boi_1 _20796_ (.A1(_03930_),
    .A2(_03932_),
    .B1_N(_03931_),
    .Y(_03935_));
 sky130_fd_sc_hd__nor2_1 _20797_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03936_));
 sky130_fd_sc_hd__nand2_1 _20798_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03937_));
 sky130_fd_sc_hd__and2b_1 _20799_ (.A_N(_03936_),
    .B(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__xnor2_1 _20800_ (.A(_03935_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__a22o_1 _20801_ (.A1(\rbzero.texV[5] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03939_),
    .X(_01605_));
 sky130_fd_sc_hd__or2_1 _20802_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .X(_03940_));
 sky130_fd_sc_hd__nand2_1 _20803_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_03941_));
 sky130_fd_sc_hd__nand2_1 _20804_ (.A(_03940_),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__o21ai_1 _20805_ (.A1(_03935_),
    .A2(_03936_),
    .B1(_03937_),
    .Y(_03943_));
 sky130_fd_sc_hd__xnor2_1 _20806_ (.A(_03942_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__a22o_1 _20807_ (.A1(\rbzero.texV[6] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03944_),
    .X(_01606_));
 sky130_fd_sc_hd__nor2_1 _20808_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03945_));
 sky130_fd_sc_hd__nand2_1 _20809_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03946_));
 sky130_fd_sc_hd__and2b_1 _20810_ (.A_N(_03945_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__a21boi_1 _20811_ (.A1(_03940_),
    .A2(_03943_),
    .B1_N(_03941_),
    .Y(_03948_));
 sky130_fd_sc_hd__xnor2_1 _20812_ (.A(_03947_),
    .B(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__a22o_1 _20813_ (.A1(\rbzero.texV[7] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03949_),
    .X(_01607_));
 sky130_fd_sc_hd__or2_1 _20814_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .X(_03950_));
 sky130_fd_sc_hd__nand2_1 _20815_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_03951_));
 sky130_fd_sc_hd__o21ai_1 _20816_ (.A1(_03945_),
    .A2(_03948_),
    .B1(_03946_),
    .Y(_03952_));
 sky130_fd_sc_hd__a21o_1 _20817_ (.A1(_03950_),
    .A2(_03951_),
    .B1(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__nand3_1 _20818_ (.A(_03950_),
    .B(_03951_),
    .C(_03952_),
    .Y(_03954_));
 sky130_fd_sc_hd__a32o_1 _20819_ (.A1(_09716_),
    .A2(_03953_),
    .A3(_03954_),
    .B1(_03861_),
    .B2(\rbzero.texV[8] ),
    .X(_01608_));
 sky130_fd_sc_hd__or2_1 _20820_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .X(_03955_));
 sky130_fd_sc_hd__nand2_1 _20821_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_03956_));
 sky130_fd_sc_hd__a21o_1 _20822_ (.A1(\rbzero.traced_texa[8] ),
    .A2(\rbzero.texV[8] ),
    .B1(_03952_),
    .X(_03957_));
 sky130_fd_sc_hd__a22o_1 _20823_ (.A1(_03955_),
    .A2(_03956_),
    .B1(_03957_),
    .B2(_03950_),
    .X(_03958_));
 sky130_fd_sc_hd__nand4_1 _20824_ (.A(_03950_),
    .B(_03955_),
    .C(_03956_),
    .D(_03957_),
    .Y(_03959_));
 sky130_fd_sc_hd__a32o_1 _20825_ (.A1(_09716_),
    .A2(_03958_),
    .A3(_03959_),
    .B1(_02731_),
    .B2(\rbzero.texV[9] ),
    .X(_01609_));
 sky130_fd_sc_hd__xnor2_1 _20826_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_03960_));
 sky130_fd_sc_hd__and3_1 _20827_ (.A(_03956_),
    .B(_03959_),
    .C(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__a21oi_1 _20828_ (.A1(_03956_),
    .A2(_03959_),
    .B1(_03960_),
    .Y(_03962_));
 sky130_fd_sc_hd__nor2_1 _20829_ (.A(_03961_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__a22o_1 _20830_ (.A1(\rbzero.texV[10] ),
    .A2(_03856_),
    .B1(_03799_),
    .B2(_03963_),
    .X(_01610_));
 sky130_fd_sc_hd__o21ai_1 _20831_ (.A1(_04472_),
    .A2(_08116_),
    .B1(_04471_),
    .Y(_03964_));
 sky130_fd_sc_hd__nand2_1 _20832_ (.A(_04471_),
    .B(_09709_),
    .Y(_03965_));
 sky130_fd_sc_hd__a21o_1 _20833_ (.A1(_04687_),
    .A2(_03965_),
    .B1(_06203_),
    .X(_03966_));
 sky130_fd_sc_hd__mux2_1 _20834_ (.A0(_03964_),
    .A1(_04471_),
    .S(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__and2_1 _20835_ (.A(_04478_),
    .B(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__clkbuf_1 _20836_ (.A(_03968_),
    .X(_01611_));
 sky130_fd_sc_hd__nand2_1 _20837_ (.A(_04472_),
    .B(_04471_),
    .Y(_03969_));
 sky130_fd_sc_hd__o211a_1 _20838_ (.A1(_03969_),
    .A2(_03966_),
    .B1(_04478_),
    .C1(_04465_),
    .X(_01612_));
 sky130_fd_sc_hd__nor2_1 _20839_ (.A(_03969_),
    .B(_03966_),
    .Y(_03970_));
 sky130_fd_sc_hd__a21oi_1 _20840_ (.A1(\rbzero.trace_state[2] ),
    .A2(_03970_),
    .B1(_08113_),
    .Y(_03971_));
 sky130_fd_sc_hd__o21a_1 _20841_ (.A1(\rbzero.trace_state[2] ),
    .A2(_03970_),
    .B1(_03971_),
    .X(_01613_));
 sky130_fd_sc_hd__o21ai_1 _20842_ (.A1(_04472_),
    .A2(_08116_),
    .B1(_04473_),
    .Y(_03972_));
 sky130_fd_sc_hd__o31a_1 _20843_ (.A1(_08406_),
    .A2(_03966_),
    .A3(_03972_),
    .B1(_01622_),
    .X(_01614_));
 sky130_fd_sc_hd__and2_2 _20844_ (.A(_03762_),
    .B(clknet_1_1__leaf__05731_),
    .X(_03973_));
 sky130_fd_sc_hd__buf_1 _20845_ (.A(_03973_),
    .X(_01615_));
 sky130_fd_sc_hd__and2_2 _20846_ (.A(_02371_),
    .B(clknet_1_1__leaf__05786_),
    .X(_03974_));
 sky130_fd_sc_hd__buf_1 _20847_ (.A(_03974_),
    .X(_01616_));
 sky130_fd_sc_hd__and2_2 _20848_ (.A(_02371_),
    .B(clknet_1_0__leaf__05839_),
    .X(_03975_));
 sky130_fd_sc_hd__buf_1 _20849_ (.A(_03975_),
    .X(_01617_));
 sky130_fd_sc_hd__and2_2 _20850_ (.A(_02371_),
    .B(clknet_1_1__leaf__05893_),
    .X(_03976_));
 sky130_fd_sc_hd__buf_1 _20851_ (.A(_03976_),
    .X(_01618_));
 sky130_fd_sc_hd__and2_2 _20852_ (.A(_02371_),
    .B(clknet_1_0__leaf__05944_),
    .X(_03977_));
 sky130_fd_sc_hd__buf_1 _20853_ (.A(_03977_),
    .X(_01619_));
 sky130_fd_sc_hd__and2_2 _20854_ (.A(_02371_),
    .B(clknet_1_0__leaf__05991_),
    .X(_03978_));
 sky130_fd_sc_hd__buf_1 _20855_ (.A(_03978_),
    .X(_01620_));
 sky130_fd_sc_hd__nor2_1 _20856_ (.A(\rbzero.hsync ),
    .B(net65),
    .Y(_01621_));
 sky130_fd_sc_hd__o2bb2ai_1 _20857_ (.A1_N(\rbzero.traced_texVinit[0] ),
    .A2_N(_09725_),
    .B1(_09731_),
    .B2(_09093_),
    .Y(_01623_));
 sky130_fd_sc_hd__a22o_1 _20858_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(_09738_),
    .B1(_09737_),
    .B2(_09086_),
    .X(_01624_));
 sky130_fd_sc_hd__a22o_1 _20859_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(_09738_),
    .B1(_09737_),
    .B2(_09082_),
    .X(_01625_));
 sky130_fd_sc_hd__a22o_1 _20860_ (.A1(\rbzero.traced_texVinit[3] ),
    .A2(_09738_),
    .B1(_09737_),
    .B2(_09834_),
    .X(_01626_));
 sky130_fd_sc_hd__buf_6 _20861_ (.A(_09728_),
    .X(_03979_));
 sky130_fd_sc_hd__inv_2 _20862_ (.A(_09324_),
    .Y(_03980_));
 sky130_fd_sc_hd__a22o_1 _20863_ (.A1(\rbzero.traced_texVinit[4] ),
    .A2(_09738_),
    .B1(_03979_),
    .B2(_03980_),
    .X(_01627_));
 sky130_fd_sc_hd__a2bb2o_1 _20864_ (.A1_N(_09446_),
    .A2_N(_09731_),
    .B1(_09725_),
    .B2(\rbzero.traced_texVinit[5] ),
    .X(_01628_));
 sky130_fd_sc_hd__buf_6 _20865_ (.A(_09724_),
    .X(_03981_));
 sky130_fd_sc_hd__a22o_1 _20866_ (.A1(\rbzero.traced_texVinit[6] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_09570_),
    .X(_01629_));
 sky130_fd_sc_hd__a2bb2o_1 _20867_ (.A1_N(_09702_),
    .A2_N(_09731_),
    .B1(_09725_),
    .B2(\rbzero.traced_texVinit[7] ),
    .X(_01630_));
 sky130_fd_sc_hd__a22o_1 _20868_ (.A1(\rbzero.traced_texVinit[8] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_09989_),
    .X(_01631_));
 sky130_fd_sc_hd__a22o_1 _20869_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_10105_),
    .X(_01632_));
 sky130_fd_sc_hd__a22o_1 _20870_ (.A1(\rbzero.traced_texVinit[10] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_10217_),
    .X(_01633_));
 sky130_fd_sc_hd__nor2_1 _20871_ (.A(\gpout0.clk_div[0] ),
    .B(net65),
    .Y(_01634_));
 sky130_fd_sc_hd__nand2_1 _20872_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .Y(_03982_));
 sky130_fd_sc_hd__or2_1 _20873_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .X(_03983_));
 sky130_fd_sc_hd__and3_1 _20874_ (.A(_02653_),
    .B(_03982_),
    .C(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__clkbuf_1 _20875_ (.A(_03984_),
    .X(_01635_));
 sky130_fd_sc_hd__xor2_1 _20876_ (.A(_05290_),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_03985_));
 sky130_fd_sc_hd__a22o_1 _20877_ (.A1(\rbzero.wall_tracer.rayAddendX[-9] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_03985_),
    .X(_01636_));
 sky130_fd_sc_hd__a22o_1 _20878_ (.A1(_05290_),
    .A2(\rbzero.wall_tracer.rayAddendX[-9] ),
    .B1(_02412_),
    .B2(_02413_),
    .X(_03986_));
 sky130_fd_sc_hd__nor2_1 _20879_ (.A(_09731_),
    .B(_02414_),
    .Y(_03987_));
 sky130_fd_sc_hd__a22o_1 _20880_ (.A1(\rbzero.wall_tracer.rayAddendX[-8] ),
    .A2(_03981_),
    .B1(_03986_),
    .B2(_03987_),
    .X(_01637_));
 sky130_fd_sc_hd__and2b_1 _20881_ (.A_N(_02411_),
    .B(_02416_),
    .X(_03988_));
 sky130_fd_sc_hd__xnor2_1 _20882_ (.A(_02415_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__a22o_1 _20883_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_03989_),
    .X(_01638_));
 sky130_fd_sc_hd__nand2_1 _20884_ (.A(_02410_),
    .B(_02418_),
    .Y(_03990_));
 sky130_fd_sc_hd__xnor2_1 _20885_ (.A(_02417_),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__a22o_1 _20886_ (.A1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_03991_),
    .X(_01639_));
 sky130_fd_sc_hd__xor2_1 _20887_ (.A(_05282_),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_03992_));
 sky130_fd_sc_hd__a22o_1 _20888_ (.A1(\rbzero.wall_tracer.rayAddendY[-9] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_03992_),
    .X(_01640_));
 sky130_fd_sc_hd__a22o_1 _20889_ (.A1(_05282_),
    .A2(\rbzero.wall_tracer.rayAddendY[-9] ),
    .B1(_03117_),
    .B2(_03118_),
    .X(_03993_));
 sky130_fd_sc_hd__a32o_1 _20890_ (.A1(_09728_),
    .A2(_03119_),
    .A3(_03993_),
    .B1(_02406_),
    .B2(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_01641_));
 sky130_fd_sc_hd__and2b_1 _20891_ (.A_N(_03116_),
    .B(_03121_),
    .X(_03994_));
 sky130_fd_sc_hd__xnor2_1 _20892_ (.A(_03120_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__a22o_1 _20893_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_03981_),
    .B1(_03979_),
    .B2(_03995_),
    .X(_01642_));
 sky130_fd_sc_hd__nand2_1 _20894_ (.A(_03115_),
    .B(_03123_),
    .Y(_03996_));
 sky130_fd_sc_hd__xnor2_1 _20895_ (.A(_03122_),
    .B(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__a22o_1 _20896_ (.A1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .A2(_02406_),
    .B1(_02478_),
    .B2(_03997_),
    .X(_01643_));
 sky130_fd_sc_hd__nor2_1 _20897_ (.A(\gpout1.clk_div[0] ),
    .B(net65),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _20898_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .Y(_03998_));
 sky130_fd_sc_hd__or2_1 _20899_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .X(_03999_));
 sky130_fd_sc_hd__and3_1 _20900_ (.A(_02653_),
    .B(_03998_),
    .C(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__clkbuf_1 _20901_ (.A(_04000_),
    .X(_01645_));
 sky130_fd_sc_hd__nor2_1 _20902_ (.A(\gpout2.clk_div[0] ),
    .B(net65),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _20903_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .Y(_04001_));
 sky130_fd_sc_hd__or2_1 _20904_ (.A(\gpout2.clk_div[0] ),
    .B(\gpout2.clk_div[1] ),
    .X(_04002_));
 sky130_fd_sc_hd__and3_1 _20905_ (.A(_02653_),
    .B(_04001_),
    .C(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__clkbuf_1 _20906_ (.A(_04003_),
    .X(_01647_));
 sky130_fd_sc_hd__nor2_1 _20907_ (.A(\gpout3.clk_div[0] ),
    .B(net65),
    .Y(_01648_));
 sky130_fd_sc_hd__nand2_1 _20908_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .Y(_04004_));
 sky130_fd_sc_hd__or2_1 _20909_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .X(_04005_));
 sky130_fd_sc_hd__and3_1 _20910_ (.A(_02653_),
    .B(_04004_),
    .C(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__clkbuf_1 _20911_ (.A(_04006_),
    .X(_01649_));
 sky130_fd_sc_hd__nor2_1 _20912_ (.A(\gpout4.clk_div[0] ),
    .B(net65),
    .Y(_01650_));
 sky130_fd_sc_hd__nand2_1 _20913_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .Y(_04007_));
 sky130_fd_sc_hd__or2_1 _20914_ (.A(\gpout4.clk_div[1] ),
    .B(\gpout4.clk_div[0] ),
    .X(_04008_));
 sky130_fd_sc_hd__and3_1 _20915_ (.A(_02653_),
    .B(_04007_),
    .C(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__clkbuf_1 _20916_ (.A(_04009_),
    .X(_01651_));
 sky130_fd_sc_hd__dfxtp_2 _20917_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00000_),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20918_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00001_),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20919_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00386_),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20920_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00387_),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20921_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00388_),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20922_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00389_),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20923_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00390_),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20924_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00391_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20925_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00392_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20926_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00393_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20927_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00394_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20928_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00395_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20929_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00396_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00397_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20931_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00398_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20932_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00399_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20933_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00400_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00401_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20935_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00402_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20936_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00403_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20937_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00404_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20938_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00405_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20939_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20940_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20941_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20942_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20943_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20944_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20945_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_4 _20946_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00413_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_4 _20947_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00414_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _20948_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00415_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20949_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00416_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _20950_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00417_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _20951_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00418_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _20952_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00419_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20953_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00420_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20954_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00421_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20955_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00422_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20956_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00423_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20957_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00424_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20958_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00425_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20959_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00426_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20960_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00427_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_4 _20961_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00428_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20962_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00429_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20963_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00430_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_4 _20964_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00431_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20965_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00432_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_4 _20966_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00433_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_4 _20967_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00434_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_2 _20969_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20970_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20973_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20976_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20977_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20979_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20984_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20985_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00457_),
    .Q(\reg_rgb[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00458_),
    .Q(\reg_rgb[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20992_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00459_),
    .Q(\reg_rgb[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20993_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00460_),
    .Q(\reg_rgb[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20994_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00461_),
    .Q(\reg_rgb[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20995_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00462_),
    .Q(\reg_rgb[23] ));
 sky130_fd_sc_hd__dfxtp_4 _20996_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00463_),
    .Q(\rbzero.wall_hot[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20997_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00464_),
    .Q(\rbzero.wall_hot[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20998_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00465_),
    .Q(\rbzero.side_hot ));
 sky130_fd_sc_hd__dfxtp_1 _20999_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00466_),
    .Q(\rbzero.texu_hot[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21000_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00467_),
    .Q(\rbzero.texu_hot[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21001_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00468_),
    .Q(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21002_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00469_),
    .Q(\rbzero.texu_hot[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21003_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00470_),
    .Q(\rbzero.texu_hot[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21004_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00471_),
    .Q(\rbzero.texu_hot[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21005_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00472_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21006_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00473_),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_4 _21007_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00474_),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21008_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00475_),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21009_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00476_),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21010_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00477_),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21011_ (.CLK(clknet_4_6_0_i_clk),
    .D(_00478_),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21012_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00479_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21013_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00480_),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_4 _21014_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00481_),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21015_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00482_),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _21016_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00483_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21017_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00484_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21018_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00485_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00486_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21020_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00487_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21021_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00488_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21022_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00489_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21023_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00490_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21024_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00491_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21025_ (.CLK(clknet_leaf_111_i_clk),
    .D(_00492_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21026_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00493_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21027_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00494_),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21028_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00495_),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21029_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00496_),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00497_),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21031_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00498_),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21032_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00499_),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21033_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00500_),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21034_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00501_),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00502_),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00503_),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21037_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00504_),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21038_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00505_),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21039_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00506_),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21040_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00507_),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21041_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00508_),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21042_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00509_),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21043_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00510_),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21044_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00511_),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21045_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00512_),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21046_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00513_),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21047_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00514_),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21048_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00515_),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21049_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00516_),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21050_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00517_),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21051_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00518_),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21052_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00519_),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21053_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00520_),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21054_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00521_),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21055_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00522_),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21056_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00523_),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21057_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00524_),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21058_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00525_),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21059_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00526_),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21060_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00527_),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21061_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00528_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21062_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00529_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00530_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00531_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00532_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00533_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00534_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21068_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00535_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00536_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00537_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21071_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00538_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00539_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21073_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00540_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21074_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21080_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21081_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21088_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21091_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21092_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21093_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21097_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21098_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21099_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21100_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21101_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21102_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21103_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21104_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21105_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00572_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21106_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00573_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21107_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00574_),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21108_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00575_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21109_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00576_),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21110_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00577_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21111_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00578_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21112_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00579_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21113_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00580_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21114_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00581_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21115_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00582_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21116_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00583_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21117_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00584_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21118_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00585_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21119_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00586_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21120_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00587_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00588_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21122_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00589_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00590_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00591_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21125_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00592_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00593_),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_2 _21127_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00594_),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_4 _21128_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00595_),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_2 _21129_ (.CLK(clknet_4_3_0_i_clk),
    .D(_00596_),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_4 _21130_ (.CLK(clknet_leaf_113_i_clk),
    .D(_00597_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21131_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00598_),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00599_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21133_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00600_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21134_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00601_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21135_ (.CLK(clknet_leaf_141_i_clk),
    .D(_00602_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21136_ (.CLK(clknet_leaf_141_i_clk),
    .D(_00603_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00604_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21138_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00605_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21139_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00606_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21140_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00607_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21141_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00608_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21142_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00609_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21143_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00610_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21144_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00611_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21145_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00612_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_4 _21146_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00613_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_4 _21147_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00614_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_4 _21148_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00615_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21149_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00616_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21150_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00617_),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _21151_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00618_),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21152_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00619_),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _21153_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00620_),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _21154_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00621_),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_2 _21155_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00622_),
    .Q(\rbzero.spi_registers.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _21156_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00623_),
    .Q(\rbzero.spi_registers.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21157_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00624_),
    .Q(\rbzero.spi_registers.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21158_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00625_),
    .Q(\rbzero.spi_registers.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21159_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00626_),
    .Q(\rbzero.spi_registers.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00627_),
    .Q(\rbzero.spi_registers.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00628_),
    .Q(\rbzero.spi_registers.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21162_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00629_),
    .Q(\rbzero.spi_registers.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21163_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00630_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21164_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00631_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00632_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21166_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00633_),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00634_),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00635_),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00636_),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00637_),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21171_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00638_),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00639_),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21173_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00640_),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00641_),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21175_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00642_),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21176_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00643_),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21177_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00644_),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00645_),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00646_),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00647_),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00648_),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21182_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00649_),
    .Q(\rbzero.map_overlay.i_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00650_),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21184_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00651_),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00652_),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00653_),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00654_),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00655_),
    .Q(\rbzero.map_overlay.i_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21189_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00656_),
    .Q(\rbzero.mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00657_),
    .Q(\rbzero.mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00658_),
    .Q(\rbzero.mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00659_),
    .Q(\rbzero.mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00660_),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00661_),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21195_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00662_),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21196_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00663_),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00664_),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21198_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00665_),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00666_),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00667_),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00668_),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00669_),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00670_),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00671_),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21205_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00672_),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21206_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00673_),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00674_),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00675_),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21209_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00676_),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21210_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00677_),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00678_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21212_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00679_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00680_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21214_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00681_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21215_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00682_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21216_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00683_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00684_),
    .Q(\rbzero.spi_registers.texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00685_),
    .Q(\rbzero.spi_registers.texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00686_),
    .Q(\rbzero.spi_registers.texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21220_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00687_),
    .Q(\rbzero.spi_registers.texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00688_),
    .Q(\rbzero.spi_registers.texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00689_),
    .Q(\rbzero.spi_registers.texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00690_),
    .Q(\rbzero.spi_registers.texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00691_),
    .Q(\rbzero.spi_registers.texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21225_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00692_),
    .Q(\rbzero.spi_registers.texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21226_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00693_),
    .Q(\rbzero.spi_registers.texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21227_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00694_),
    .Q(\rbzero.spi_registers.texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00695_),
    .Q(\rbzero.spi_registers.texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00696_),
    .Q(\rbzero.spi_registers.texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00697_),
    .Q(\rbzero.spi_registers.texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00698_),
    .Q(\rbzero.spi_registers.texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00699_),
    .Q(\rbzero.spi_registers.texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00700_),
    .Q(\rbzero.spi_registers.texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00701_),
    .Q(\rbzero.spi_registers.texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00702_),
    .Q(\rbzero.spi_registers.texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00703_),
    .Q(\rbzero.spi_registers.texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00704_),
    .Q(\rbzero.spi_registers.texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00705_),
    .Q(\rbzero.spi_registers.texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00706_),
    .Q(\rbzero.spi_registers.texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00707_),
    .Q(\rbzero.spi_registers.texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00708_),
    .Q(\rbzero.spi_registers.texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00709_),
    .Q(\rbzero.spi_registers.texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00710_),
    .Q(\rbzero.spi_registers.texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00711_),
    .Q(\rbzero.spi_registers.texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21245_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00712_),
    .Q(\rbzero.spi_registers.texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00713_),
    .Q(\rbzero.spi_registers.texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21247_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00714_),
    .Q(\rbzero.spi_registers.texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21248_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00715_),
    .Q(\rbzero.spi_registers.texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00716_),
    .Q(\rbzero.spi_registers.texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00717_),
    .Q(\rbzero.spi_registers.texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00718_),
    .Q(\rbzero.spi_registers.texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00719_),
    .Q(\rbzero.spi_registers.texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00720_),
    .Q(\rbzero.spi_registers.texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00721_),
    .Q(\rbzero.spi_registers.texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00722_),
    .Q(\rbzero.spi_registers.texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00723_),
    .Q(\rbzero.spi_registers.texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00724_),
    .Q(\rbzero.spi_registers.texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21258_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00725_),
    .Q(\rbzero.spi_registers.texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21259_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00726_),
    .Q(\rbzero.spi_registers.texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21260_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00727_),
    .Q(\rbzero.spi_registers.texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21261_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00728_),
    .Q(\rbzero.spi_registers.texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21262_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00729_),
    .Q(\rbzero.spi_registers.texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00730_),
    .Q(\rbzero.spi_registers.texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21264_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00731_),
    .Q(\rbzero.spi_registers.texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00732_),
    .Q(\rbzero.spi_registers.texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00733_),
    .Q(\rbzero.spi_registers.texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21267_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00734_),
    .Q(\rbzero.spi_registers.texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00735_),
    .Q(\rbzero.spi_registers.texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21269_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00736_),
    .Q(\rbzero.spi_registers.texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00737_),
    .Q(\rbzero.spi_registers.texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00738_),
    .Q(\rbzero.spi_registers.texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00739_),
    .Q(\rbzero.spi_registers.texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00740_),
    .Q(\rbzero.spi_registers.texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00741_),
    .Q(\rbzero.spi_registers.texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21275_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00742_),
    .Q(\rbzero.spi_registers.texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21276_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00743_),
    .Q(\rbzero.spi_registers.texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21277_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00744_),
    .Q(\rbzero.spi_registers.texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21278_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00745_),
    .Q(\rbzero.spi_registers.texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00746_),
    .Q(\rbzero.spi_registers.texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21280_ (.CLK(clknet_leaf_143_i_clk),
    .D(_00747_),
    .Q(\rbzero.spi_registers.texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(clknet_leaf_143_i_clk),
    .D(_00748_),
    .Q(\rbzero.spi_registers.texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00749_),
    .Q(\rbzero.spi_registers.texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00750_),
    .Q(\rbzero.spi_registers.texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00751_),
    .Q(\rbzero.spi_registers.texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00752_),
    .Q(\rbzero.spi_registers.texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00753_),
    .Q(\rbzero.spi_registers.texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00754_),
    .Q(\rbzero.spi_registers.texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00755_),
    .Q(\rbzero.spi_registers.texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00756_),
    .Q(\rbzero.spi_registers.texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00757_),
    .Q(\rbzero.spi_registers.texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00758_),
    .Q(\rbzero.spi_registers.texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00759_),
    .Q(\rbzero.spi_registers.texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21293_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00760_),
    .Q(\rbzero.spi_registers.texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21294_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00761_),
    .Q(\rbzero.spi_registers.texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00762_),
    .Q(\rbzero.spi_registers.texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00763_),
    .Q(\rbzero.spi_registers.texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21297_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00764_),
    .Q(\rbzero.spi_registers.texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00765_),
    .Q(\rbzero.spi_registers.texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00766_),
    .Q(\rbzero.spi_registers.texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00767_),
    .Q(\rbzero.spi_registers.texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21301_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00768_),
    .Q(\rbzero.spi_registers.texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00769_),
    .Q(\rbzero.spi_registers.texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00770_),
    .Q(\rbzero.spi_registers.texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00771_),
    .Q(\rbzero.spi_registers.texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00772_),
    .Q(\rbzero.spi_registers.texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(clknet_leaf_141_i_clk),
    .D(_00773_),
    .Q(\rbzero.spi_registers.texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00774_),
    .Q(\rbzero.spi_registers.texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(clknet_leaf_141_i_clk),
    .D(_00775_),
    .Q(\rbzero.spi_registers.texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21309_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00776_),
    .Q(\rbzero.spi_registers.texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21310_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00777_),
    .Q(\rbzero.spi_registers.texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00778_),
    .Q(\rbzero.spi_registers.texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00779_),
    .Q(\rbzero.spi_registers.texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00780_),
    .Q(\rbzero.spi_registers.buf_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00781_),
    .Q(\rbzero.spi_registers.buf_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00782_),
    .Q(\rbzero.spi_registers.buf_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00783_),
    .Q(\rbzero.spi_registers.buf_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00784_),
    .Q(\rbzero.spi_registers.buf_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00785_),
    .Q(\rbzero.spi_registers.buf_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00786_),
    .Q(\rbzero.spi_registers.buf_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00787_),
    .Q(\rbzero.spi_registers.buf_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00788_),
    .Q(\rbzero.spi_registers.buf_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00789_),
    .Q(\rbzero.spi_registers.buf_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(clknet_leaf_42_i_clk),
    .D(_00790_),
    .Q(\rbzero.spi_registers.buf_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00791_),
    .Q(\rbzero.spi_registers.buf_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00792_),
    .Q(\rbzero.spi_registers.buf_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00793_),
    .Q(\rbzero.spi_registers.buf_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00794_),
    .Q(\rbzero.spi_registers.buf_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(clknet_leaf_39_i_clk),
    .D(_00795_),
    .Q(\rbzero.spi_registers.buf_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00796_),
    .Q(\rbzero.spi_registers.buf_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00797_),
    .Q(\rbzero.spi_registers.buf_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00798_),
    .Q(\rbzero.spi_registers.buf_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00799_),
    .Q(\rbzero.spi_registers.buf_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00800_),
    .Q(\rbzero.spi_registers.buf_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00801_),
    .Q(\rbzero.spi_registers.buf_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00802_),
    .Q(\rbzero.spi_registers.buf_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00803_),
    .Q(\rbzero.spi_registers.buf_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00804_),
    .Q(\rbzero.spi_registers.buf_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00805_),
    .Q(\rbzero.spi_registers.buf_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00806_),
    .Q(\rbzero.spi_registers.buf_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00807_),
    .Q(\rbzero.spi_registers.buf_othery[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(clknet_leaf_40_i_clk),
    .D(_00808_),
    .Q(\rbzero.spi_registers.buf_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00809_),
    .Q(\rbzero.spi_registers.buf_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00810_),
    .Q(\rbzero.spi_registers.buf_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00811_),
    .Q(\rbzero.spi_registers.buf_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00812_),
    .Q(\rbzero.spi_registers.buf_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00813_),
    .Q(\rbzero.spi_registers.buf_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00814_),
    .Q(\rbzero.spi_registers.buf_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00815_),
    .Q(\rbzero.spi_registers.buf_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00816_),
    .Q(\rbzero.spi_registers.buf_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00817_),
    .Q(\rbzero.spi_registers.buf_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00818_),
    .Q(\rbzero.spi_registers.buf_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00819_),
    .Q(\rbzero.spi_registers.buf_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00820_),
    .Q(\rbzero.spi_registers.buf_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00821_),
    .Q(\rbzero.spi_registers.buf_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00822_),
    .Q(\rbzero.spi_registers.buf_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00823_),
    .Q(\rbzero.spi_registers.buf_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00824_),
    .Q(\rbzero.spi_registers.buf_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00825_),
    .Q(\rbzero.spi_registers.buf_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00826_),
    .Q(\rbzero.spi_registers.buf_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00827_),
    .Q(\rbzero.spi_registers.buf_mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00828_),
    .Q(\rbzero.spi_registers.buf_mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00829_),
    .Q(\rbzero.spi_registers.buf_mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00830_),
    .Q(\rbzero.spi_registers.buf_mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00831_),
    .Q(\rbzero.spi_registers.buf_texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00832_),
    .Q(\rbzero.spi_registers.buf_texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00833_),
    .Q(\rbzero.spi_registers.buf_texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00834_),
    .Q(\rbzero.spi_registers.buf_texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00835_),
    .Q(\rbzero.spi_registers.buf_texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00836_),
    .Q(\rbzero.spi_registers.buf_texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00837_),
    .Q(\rbzero.spi_registers.buf_texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00838_),
    .Q(\rbzero.spi_registers.buf_texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00839_),
    .Q(\rbzero.spi_registers.buf_texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00840_),
    .Q(\rbzero.spi_registers.buf_texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00841_),
    .Q(\rbzero.spi_registers.buf_texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00842_),
    .Q(\rbzero.spi_registers.buf_texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00843_),
    .Q(\rbzero.spi_registers.buf_texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00844_),
    .Q(\rbzero.spi_registers.buf_texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00845_),
    .Q(\rbzero.spi_registers.buf_texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00846_),
    .Q(\rbzero.spi_registers.buf_texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00847_),
    .Q(\rbzero.spi_registers.buf_texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00848_),
    .Q(\rbzero.spi_registers.buf_texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00849_),
    .Q(\rbzero.spi_registers.buf_texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00850_),
    .Q(\rbzero.spi_registers.buf_texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00851_),
    .Q(\rbzero.spi_registers.buf_texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00852_),
    .Q(\rbzero.spi_registers.buf_texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00853_),
    .Q(\rbzero.spi_registers.buf_texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00854_),
    .Q(\rbzero.spi_registers.buf_texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00855_),
    .Q(\rbzero.spi_registers.buf_texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00856_),
    .Q(\rbzero.spi_registers.buf_texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00857_),
    .Q(\rbzero.spi_registers.buf_texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00858_),
    .Q(\rbzero.spi_registers.buf_texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00859_),
    .Q(\rbzero.spi_registers.buf_texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00860_),
    .Q(\rbzero.spi_registers.buf_texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00861_),
    .Q(\rbzero.spi_registers.buf_texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00862_),
    .Q(\rbzero.spi_registers.buf_texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00863_),
    .Q(\rbzero.spi_registers.buf_texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00864_),
    .Q(\rbzero.spi_registers.buf_texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00865_),
    .Q(\rbzero.spi_registers.buf_texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00866_),
    .Q(\rbzero.spi_registers.buf_texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00867_),
    .Q(\rbzero.spi_registers.buf_texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00868_),
    .Q(\rbzero.spi_registers.buf_texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00869_),
    .Q(\rbzero.spi_registers.buf_texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00870_),
    .Q(\rbzero.spi_registers.buf_texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00871_),
    .Q(\rbzero.spi_registers.buf_texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00872_),
    .Q(\rbzero.spi_registers.buf_texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00873_),
    .Q(\rbzero.spi_registers.buf_texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00874_),
    .Q(\rbzero.spi_registers.buf_texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00875_),
    .Q(\rbzero.spi_registers.buf_texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21409_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00876_),
    .Q(\rbzero.spi_registers.buf_texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21410_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00877_),
    .Q(\rbzero.spi_registers.buf_texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21411_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00878_),
    .Q(\rbzero.spi_registers.buf_texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21412_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00879_),
    .Q(\rbzero.spi_registers.buf_texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21413_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00880_),
    .Q(\rbzero.spi_registers.buf_texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00881_),
    .Q(\rbzero.spi_registers.buf_texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00882_),
    .Q(\rbzero.spi_registers.buf_texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21416_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00883_),
    .Q(\rbzero.spi_registers.buf_texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00884_),
    .Q(\rbzero.spi_registers.buf_texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00885_),
    .Q(\rbzero.spi_registers.buf_texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21419_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00886_),
    .Q(\rbzero.spi_registers.buf_texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00887_),
    .Q(\rbzero.spi_registers.buf_texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00888_),
    .Q(\rbzero.spi_registers.buf_texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00889_),
    .Q(\rbzero.spi_registers.buf_texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00890_),
    .Q(\rbzero.spi_registers.buf_texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21424_ (.CLK(clknet_leaf_144_i_clk),
    .D(_00891_),
    .Q(\rbzero.spi_registers.buf_texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21425_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00892_),
    .Q(\rbzero.spi_registers.buf_texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(clknet_leaf_143_i_clk),
    .D(_00893_),
    .Q(\rbzero.spi_registers.buf_texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(clknet_leaf_143_i_clk),
    .D(_00894_),
    .Q(\rbzero.spi_registers.buf_texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(clknet_leaf_143_i_clk),
    .D(_00895_),
    .Q(\rbzero.spi_registers.buf_texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(clknet_leaf_143_i_clk),
    .D(_00896_),
    .Q(\rbzero.spi_registers.buf_texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(clknet_leaf_143_i_clk),
    .D(_00897_),
    .Q(\rbzero.spi_registers.buf_texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21431_ (.CLK(clknet_leaf_142_i_clk),
    .D(_00898_),
    .Q(\rbzero.spi_registers.buf_texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21432_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00899_),
    .Q(\rbzero.spi_registers.buf_texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21433_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00900_),
    .Q(\rbzero.spi_registers.buf_texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21434_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00901_),
    .Q(\rbzero.spi_registers.buf_texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00902_),
    .Q(\rbzero.spi_registers.buf_texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21436_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00903_),
    .Q(\rbzero.spi_registers.buf_texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21437_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00904_),
    .Q(\rbzero.spi_registers.buf_texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21438_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00905_),
    .Q(\rbzero.spi_registers.buf_texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00906_),
    .Q(\rbzero.spi_registers.buf_texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21440_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00907_),
    .Q(\rbzero.spi_registers.buf_texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21441_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00908_),
    .Q(\rbzero.spi_registers.buf_texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00909_),
    .Q(\rbzero.spi_registers.buf_texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00910_),
    .Q(\rbzero.spi_registers.buf_texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00911_),
    .Q(\rbzero.spi_registers.buf_texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00912_),
    .Q(\rbzero.spi_registers.buf_texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00913_),
    .Q(\rbzero.spi_registers.buf_texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21447_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00914_),
    .Q(\rbzero.spi_registers.buf_texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00915_),
    .Q(\rbzero.spi_registers.buf_texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00916_),
    .Q(\rbzero.spi_registers.buf_texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21450_ (.CLK(clknet_leaf_141_i_clk),
    .D(_00917_),
    .Q(\rbzero.spi_registers.buf_texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(clknet_leaf_142_i_clk),
    .D(_00918_),
    .Q(\rbzero.spi_registers.buf_texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00919_),
    .Q(\rbzero.spi_registers.buf_texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(clknet_leaf_142_i_clk),
    .D(_00920_),
    .Q(\rbzero.spi_registers.buf_texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00921_),
    .Q(\rbzero.spi_registers.buf_texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00922_),
    .Q(\rbzero.spi_registers.buf_texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00923_),
    .Q(\rbzero.spi_registers.buf_texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00924_),
    .Q(\rbzero.spi_registers.buf_texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00925_),
    .Q(\rbzero.spi_registers.buf_texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00926_),
    .Q(\rbzero.spi_registers.buf_texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_2 _21460_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00927_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21461_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00928_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21462_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00929_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21463_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00930_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00931_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21465_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00932_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00933_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00934_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21468_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00935_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21469_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00936_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21470_ (.CLK(clknet_4_5_0_i_clk),
    .D(_00937_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00938_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21472_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00939_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21473_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00940_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21474_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00941_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00942_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21476_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00943_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00944_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00945_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00946_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00947_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00948_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00949_),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_1 _21483_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00950_),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00951_),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00952_),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_2 _21486_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00953_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00954_),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21488_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00955_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_4 _21489_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00956_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21490_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00957_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21491_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00958_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21492_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00959_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21493_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00960_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00961_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21495_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00962_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _21496_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00963_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21497_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00964_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21498_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00965_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21499_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00966_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21500_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00967_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21501_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00968_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21502_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00969_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21503_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00970_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21504_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00971_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(clknet_leaf_106_i_clk),
    .D(_00972_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21506_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00973_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00974_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00975_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(clknet_leaf_109_i_clk),
    .D(_00976_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21510_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00977_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21511_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00978_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21512_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00979_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21513_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00980_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21514_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00981_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21515_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00982_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21516_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00983_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21517_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00984_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21518_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00985_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00986_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00987_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21521_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00988_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21522_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00989_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21523_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00990_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21524_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00991_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00992_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00993_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(clknet_leaf_108_i_clk),
    .D(_00994_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21528_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00995_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21529_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00996_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00997_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21531_ (.CLK(clknet_leaf_101_i_clk),
    .D(_00998_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21532_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00999_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01000_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _21534_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01001_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21535_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01002_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01003_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21537_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01004_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01005_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21539_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01006_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01007_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_4 _21541_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01008_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21542_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01009_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_4 _21543_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01010_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01011_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21545_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01012_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21546_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01013_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01014_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_4 _21548_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01015_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01016_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21550_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01017_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01018_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21552_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01019_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21553_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01020_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_2 _21554_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01021_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01022_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21556_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01023_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21557_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01024_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21558_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01025_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21559_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01026_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(clknet_leaf_102_i_clk),
    .D(_01027_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(clknet_leaf_102_i_clk),
    .D(_01028_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(clknet_leaf_139_i_clk),
    .D(_01029_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01030_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01031_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01032_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21566_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01033_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01034_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21568_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01035_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01036_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01037_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01038_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21572_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01039_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01040_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01041_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01042_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01043_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21577_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01044_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21578_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01045_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21579_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01046_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01047_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21581_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01048_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21582_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01049_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01050_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21584_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01051_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21585_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01052_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21586_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01053_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21587_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01054_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21588_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01055_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21589_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01056_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21590_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01057_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21591_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01058_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01059_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21593_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01060_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21594_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01061_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01062_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21596_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01063_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21597_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01064_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01065_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21599_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01066_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21600_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01067_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21601_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01068_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21602_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01069_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21603_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01070_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21604_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01071_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21605_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01072_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21606_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01073_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01074_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01075_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21609_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01076_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01077_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01078_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01079_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01080_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21614_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01081_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01082_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01083_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01084_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21618_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01085_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21619_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01086_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01087_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01088_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01089_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01090_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01091_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01092_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21626_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01093_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01094_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01095_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21629_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01096_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21630_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01097_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21631_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01098_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21632_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01099_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01100_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21634_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01101_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21635_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01102_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21636_ (.CLK(clknet_leaf_139_i_clk),
    .D(_01103_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21637_ (.CLK(clknet_leaf_139_i_clk),
    .D(_01104_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21638_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01105_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01106_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21640_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01107_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21641_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01108_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21642_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01109_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21643_ (.CLK(net154),
    .D(_01110_),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(net155),
    .D(_01111_),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21645_ (.CLK(net156),
    .D(_01112_),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21646_ (.CLK(net157),
    .D(_01113_),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21647_ (.CLK(net158),
    .D(_01114_),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21648_ (.CLK(net159),
    .D(_01115_),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21649_ (.CLK(net160),
    .D(_01116_),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21650_ (.CLK(net161),
    .D(_01117_),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21651_ (.CLK(net162),
    .D(_01118_),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(net163),
    .D(_01119_),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(net164),
    .D(_01120_),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(net165),
    .D(_01121_),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21655_ (.CLK(net166),
    .D(_01122_),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(net167),
    .D(_01123_),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(net168),
    .D(_01124_),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(net169),
    .D(_01125_),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21659_ (.CLK(net170),
    .D(_01126_),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(net171),
    .D(_01127_),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(net172),
    .D(_01128_),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(net173),
    .D(_01129_),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(net174),
    .D(_01130_),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(net175),
    .D(_01131_),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(net176),
    .D(_01132_),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(net177),
    .D(_01133_),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21667_ (.CLK(net178),
    .D(_01134_),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(net179),
    .D(_01135_),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21669_ (.CLK(net180),
    .D(_01136_),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21670_ (.CLK(net181),
    .D(_01137_),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21671_ (.CLK(net182),
    .D(_01138_),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21672_ (.CLK(net183),
    .D(_01139_),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21673_ (.CLK(net184),
    .D(_01140_),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21674_ (.CLK(net185),
    .D(_01141_),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21675_ (.CLK(net186),
    .D(_01142_),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(net187),
    .D(_01143_),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21677_ (.CLK(net188),
    .D(_01144_),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(net189),
    .D(_01145_),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(net190),
    .D(_01146_),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(net191),
    .D(_01147_),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(net192),
    .D(_01148_),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21682_ (.CLK(net193),
    .D(_01149_),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(net194),
    .D(_01150_),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(net195),
    .D(_01151_),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21685_ (.CLK(net196),
    .D(_01152_),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21686_ (.CLK(net197),
    .D(_01153_),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21687_ (.CLK(net198),
    .D(_01154_),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(net199),
    .D(_01155_),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21689_ (.CLK(net200),
    .D(_01156_),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21690_ (.CLK(net201),
    .D(_01157_),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21691_ (.CLK(net202),
    .D(_01158_),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(net203),
    .D(_01159_),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21693_ (.CLK(net204),
    .D(_01160_),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21694_ (.CLK(net205),
    .D(_01161_),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21695_ (.CLK(net206),
    .D(_01162_),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21696_ (.CLK(net207),
    .D(_01163_),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(net208),
    .D(_01164_),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21698_ (.CLK(net209),
    .D(_01165_),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21699_ (.CLK(net210),
    .D(_01166_),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(net211),
    .D(_01167_),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(net212),
    .D(_01168_),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21702_ (.CLK(net213),
    .D(_01169_),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21703_ (.CLK(net214),
    .D(_01170_),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21704_ (.CLK(net215),
    .D(_01171_),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21705_ (.CLK(net216),
    .D(_01172_),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21706_ (.CLK(net217),
    .D(_01173_),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21707_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01174_),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _21708_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01175_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21709_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01176_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21710_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01177_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21711_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01178_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21712_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01179_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21713_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01180_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21714_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01181_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21715_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01182_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21716_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01183_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21717_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01184_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21718_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01185_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21719_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01186_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21720_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01187_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21721_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01188_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21722_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01189_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21723_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01190_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21724_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01191_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21725_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01192_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21726_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01193_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21727_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01194_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01195_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01196_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01197_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21731_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01198_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21732_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01199_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21733_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01200_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21734_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01201_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21735_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01202_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21736_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01203_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21737_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01204_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21738_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01205_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21739_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01206_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21740_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01207_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21741_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01208_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21742_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01209_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21743_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01210_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21744_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01211_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21745_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01212_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21746_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01213_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21747_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01214_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21748_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01215_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21749_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01216_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21750_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01217_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21751_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01218_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21752_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01219_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21753_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01220_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21754_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01221_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21755_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01222_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21756_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01223_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21757_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01224_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21758_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01225_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21759_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01226_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01227_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01228_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21762_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01229_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21763_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01230_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21764_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01231_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21765_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01232_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21766_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01233_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21767_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01234_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21768_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01235_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21769_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01236_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21770_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01237_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21771_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01238_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21772_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01239_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21773_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01240_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01241_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21775_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01242_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21776_ (.CLK(clknet_leaf_139_i_clk),
    .D(_01243_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21777_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01244_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21778_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01245_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21779_ (.CLK(clknet_leaf_139_i_clk),
    .D(_01246_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01247_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21781_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01248_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21782_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01249_),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21783_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01250_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21784_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01251_),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01252_),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _21786_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01253_),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_2 _21787_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01254_),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21788_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01255_),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21789_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01256_),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21790_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01257_),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21791_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01258_),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21792_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01259_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21793_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01260_),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21794_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01261_),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21795_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01262_),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21796_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01263_),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01264_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21798_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01265_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21799_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01266_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21800_ (.CLK(net218),
    .D(_01267_),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(net219),
    .D(_01268_),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21802_ (.CLK(net220),
    .D(_01269_),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21803_ (.CLK(net221),
    .D(_01270_),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21804_ (.CLK(net222),
    .D(_01271_),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(net223),
    .D(_01272_),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(net224),
    .D(_01273_),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21807_ (.CLK(net225),
    .D(_01274_),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(net226),
    .D(_01275_),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(net227),
    .D(_01276_),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(net228),
    .D(_01277_),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(net229),
    .D(_01278_),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(net230),
    .D(_01279_),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(net231),
    .D(_01280_),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(net232),
    .D(_01281_),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21815_ (.CLK(net233),
    .D(_01282_),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21816_ (.CLK(net234),
    .D(_01283_),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21817_ (.CLK(net235),
    .D(_01284_),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(net236),
    .D(_01285_),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21819_ (.CLK(net237),
    .D(_01286_),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21820_ (.CLK(net238),
    .D(_01287_),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(net239),
    .D(_01288_),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21822_ (.CLK(net240),
    .D(_01289_),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21823_ (.CLK(net241),
    .D(_01290_),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21824_ (.CLK(net242),
    .D(_01291_),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21825_ (.CLK(net243),
    .D(_01292_),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21826_ (.CLK(net244),
    .D(_01293_),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21827_ (.CLK(net245),
    .D(_01294_),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21828_ (.CLK(net246),
    .D(_01295_),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21829_ (.CLK(net247),
    .D(_01296_),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21830_ (.CLK(net248),
    .D(_01297_),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21831_ (.CLK(net249),
    .D(_01298_),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21832_ (.CLK(net250),
    .D(_01299_),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21833_ (.CLK(net251),
    .D(_01300_),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(net252),
    .D(_01301_),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(net253),
    .D(_01302_),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(net254),
    .D(_01303_),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(net255),
    .D(_01304_),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(net256),
    .D(_01305_),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21839_ (.CLK(net257),
    .D(_01306_),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(net258),
    .D(_01307_),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21841_ (.CLK(net259),
    .D(_01308_),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21842_ (.CLK(net260),
    .D(_01309_),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21843_ (.CLK(net261),
    .D(_01310_),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21844_ (.CLK(net262),
    .D(_01311_),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(net263),
    .D(_01312_),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21846_ (.CLK(net264),
    .D(_01313_),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21847_ (.CLK(net265),
    .D(_01314_),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21848_ (.CLK(net266),
    .D(_01315_),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(net267),
    .D(_01316_),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(net268),
    .D(_01317_),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(net269),
    .D(_01318_),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(net270),
    .D(_01319_),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21853_ (.CLK(net271),
    .D(_01320_),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(net272),
    .D(_01321_),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(net273),
    .D(_01322_),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(net274),
    .D(_01323_),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(net275),
    .D(_01324_),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(net276),
    .D(_01325_),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(net277),
    .D(_01326_),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(net278),
    .D(_01327_),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(net279),
    .D(_01328_),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(net280),
    .D(_01329_),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21863_ (.CLK(net281),
    .D(_01330_),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(net282),
    .D(_01331_),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(net283),
    .D(_01332_),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(net284),
    .D(_01333_),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(net285),
    .D(_01334_),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(net286),
    .D(_01335_),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(net287),
    .D(_01336_),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(net288),
    .D(_01337_),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(net289),
    .D(_01338_),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(net290),
    .D(_01339_),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21873_ (.CLK(net291),
    .D(_01340_),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21874_ (.CLK(net292),
    .D(_01341_),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(net293),
    .D(_01342_),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(net294),
    .D(_01343_),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(net295),
    .D(_01344_),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21878_ (.CLK(net296),
    .D(_01345_),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21879_ (.CLK(net297),
    .D(_01346_),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21880_ (.CLK(net298),
    .D(_01347_),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(net299),
    .D(_01348_),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21882_ (.CLK(net300),
    .D(_01349_),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(net301),
    .D(_01350_),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(net302),
    .D(_01351_),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(net303),
    .D(_01352_),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(net304),
    .D(_01353_),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(net305),
    .D(_01354_),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(net306),
    .D(_01355_),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(net307),
    .D(_01356_),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(net308),
    .D(_01357_),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(net309),
    .D(_01358_),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(net310),
    .D(_01359_),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(net311),
    .D(_01360_),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(net312),
    .D(_01361_),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21895_ (.CLK(net313),
    .D(_01362_),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(net314),
    .D(_01363_),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(net315),
    .D(_01364_),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21898_ (.CLK(net316),
    .D(_01365_),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(net317),
    .D(_01366_),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(net318),
    .D(_01367_),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(net319),
    .D(_01368_),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(net320),
    .D(_01369_),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(net321),
    .D(_01370_),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(net322),
    .D(_01371_),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(net323),
    .D(_01372_),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(net324),
    .D(_01373_),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(net325),
    .D(_01374_),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(net326),
    .D(_01375_),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21909_ (.CLK(net327),
    .D(_01376_),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(net328),
    .D(_01377_),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21911_ (.CLK(net329),
    .D(_01378_),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(net330),
    .D(_01379_),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(net331),
    .D(_01380_),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(net332),
    .D(_01381_),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21915_ (.CLK(net333),
    .D(_01382_),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(net334),
    .D(_01383_),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(net335),
    .D(_01384_),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(net336),
    .D(_01385_),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(net337),
    .D(_01386_),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(net338),
    .D(_01387_),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(net339),
    .D(_01388_),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(net340),
    .D(_01389_),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(net341),
    .D(_01390_),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(net342),
    .D(_01391_),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(net343),
    .D(_01392_),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21926_ (.CLK(net344),
    .D(_01393_),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(net345),
    .D(_01394_),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(net346),
    .D(_01395_),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(net347),
    .D(_01396_),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21930_ (.CLK(net348),
    .D(_01397_),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21931_ (.CLK(net349),
    .D(_01398_),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(net350),
    .D(_01399_),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(net351),
    .D(_01400_),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(net352),
    .D(_01401_),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(net353),
    .D(_01402_),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(net354),
    .D(_01403_),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(net355),
    .D(_01404_),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(net356),
    .D(_01405_),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(net357),
    .D(_01406_),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(net358),
    .D(_01407_),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(net359),
    .D(_01408_),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(net360),
    .D(_01409_),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(net361),
    .D(_01410_),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21944_ (.CLK(net362),
    .D(_01411_),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(net363),
    .D(_01412_),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21946_ (.CLK(net364),
    .D(_01413_),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21947_ (.CLK(net365),
    .D(_01414_),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21948_ (.CLK(net366),
    .D(_01415_),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21949_ (.CLK(net367),
    .D(_01416_),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21950_ (.CLK(net368),
    .D(_01417_),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(net369),
    .D(_01418_),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(net370),
    .D(_01419_),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(net371),
    .D(_01420_),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(net372),
    .D(_01421_),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(net373),
    .D(_01422_),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(net374),
    .D(_01423_),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(net375),
    .D(_01424_),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21958_ (.CLK(net376),
    .D(_01425_),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(net377),
    .D(_01426_),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21960_ (.CLK(net378),
    .D(_01427_),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(net379),
    .D(_01428_),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(net380),
    .D(_01429_),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21963_ (.CLK(net381),
    .D(_01430_),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(net382),
    .D(_01431_),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(net383),
    .D(_01432_),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(net384),
    .D(_01433_),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21967_ (.CLK(net385),
    .D(_01434_),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(net386),
    .D(_01435_),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(net387),
    .D(_01436_),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(net388),
    .D(_01437_),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21971_ (.CLK(net389),
    .D(_01438_),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(net390),
    .D(_01439_),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(net391),
    .D(_01440_),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(net392),
    .D(_01441_),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(net393),
    .D(_01442_),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(net394),
    .D(_01443_),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(net395),
    .D(_01444_),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(net396),
    .D(_01445_),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(net397),
    .D(_01446_),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(net398),
    .D(_01447_),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(net399),
    .D(_01448_),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(net400),
    .D(_01449_),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(net401),
    .D(_01450_),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(net402),
    .D(_01451_),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(net403),
    .D(_01452_),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(net404),
    .D(_01453_),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(net405),
    .D(_01454_),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(net406),
    .D(_01455_),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(net407),
    .D(_01456_),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(net408),
    .D(_01457_),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21991_ (.CLK(net409),
    .D(_01458_),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21992_ (.CLK(net410),
    .D(_01459_),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(net411),
    .D(_01460_),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(net412),
    .D(_01461_),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(net413),
    .D(_01462_),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(net414),
    .D(_01463_),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(net415),
    .D(_01464_),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21998_ (.CLK(net416),
    .D(_01465_),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(net417),
    .D(_01466_),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(net418),
    .D(_01467_),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(net419),
    .D(_01468_),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(net420),
    .D(_01469_),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(net421),
    .D(_01470_),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(net422),
    .D(_01471_),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(net423),
    .D(_01472_),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(net424),
    .D(_01473_),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(net425),
    .D(_01474_),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(net426),
    .D(_01475_),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(net427),
    .D(_01476_),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(net428),
    .D(_01477_),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(net429),
    .D(_01478_),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22012_ (.CLK(net430),
    .D(_01479_),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22013_ (.CLK(net431),
    .D(_01480_),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(net432),
    .D(_01481_),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(net433),
    .D(_01482_),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(net434),
    .D(_01483_),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(net435),
    .D(_01484_),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(net436),
    .D(_01485_),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(net437),
    .D(_01486_),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(net438),
    .D(_01487_),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(net439),
    .D(_01488_),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22022_ (.CLK(net440),
    .D(_01489_),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(net441),
    .D(_01490_),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(net442),
    .D(_01491_),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(net443),
    .D(_01492_),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(net444),
    .D(_01493_),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(net445),
    .D(_01494_),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(net446),
    .D(_01495_),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(net447),
    .D(_01496_),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(net448),
    .D(_01497_),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(net449),
    .D(_01498_),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(net450),
    .D(_01499_),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22033_ (.CLK(net451),
    .D(_01500_),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(net452),
    .D(_01501_),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(net453),
    .D(_01502_),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22036_ (.CLK(net454),
    .D(_01503_),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(net455),
    .D(_01504_),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(net456),
    .D(_01505_),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(net457),
    .D(_01506_),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(net458),
    .D(_01507_),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(net459),
    .D(_01508_),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(net460),
    .D(_01509_),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(net461),
    .D(_01510_),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(net462),
    .D(_01511_),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(net463),
    .D(_01512_),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22046_ (.CLK(net464),
    .D(_01513_),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22047_ (.CLK(net465),
    .D(_01514_),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22048_ (.CLK(net466),
    .D(_01515_),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22049_ (.CLK(net467),
    .D(_01516_),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22050_ (.CLK(net468),
    .D(_01517_),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22051_ (.CLK(net469),
    .D(_01518_),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22052_ (.CLK(net470),
    .D(_01519_),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22053_ (.CLK(net471),
    .D(_01520_),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22054_ (.CLK(net472),
    .D(_01521_),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22055_ (.CLK(net473),
    .D(_01522_),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22056_ (.CLK(net474),
    .D(_01523_),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22057_ (.CLK(net475),
    .D(_01524_),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22058_ (.CLK(net476),
    .D(_01525_),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22059_ (.CLK(net477),
    .D(_01526_),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22060_ (.CLK(net478),
    .D(_01527_),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22061_ (.CLK(net479),
    .D(_01528_),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22062_ (.CLK(net480),
    .D(_01529_),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22063_ (.CLK(net481),
    .D(_01530_),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22064_ (.CLK(net482),
    .D(_01531_),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22065_ (.CLK(net483),
    .D(_01532_),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22066_ (.CLK(net484),
    .D(_01533_),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22067_ (.CLK(net485),
    .D(_01534_),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22068_ (.CLK(net486),
    .D(_01535_),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22069_ (.CLK(net487),
    .D(_01536_),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22070_ (.CLK(net488),
    .D(_01537_),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22071_ (.CLK(net489),
    .D(_01538_),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22072_ (.CLK(net490),
    .D(_01539_),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22073_ (.CLK(net491),
    .D(_01540_),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22074_ (.CLK(net492),
    .D(_01541_),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22075_ (.CLK(net493),
    .D(_01542_),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _22076_ (.CLK(net494),
    .D(_01543_),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22077_ (.CLK(net495),
    .D(_01544_),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22078_ (.CLK(net496),
    .D(_01545_),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22079_ (.CLK(net497),
    .D(_01546_),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22080_ (.CLK(net498),
    .D(_01547_),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22081_ (.CLK(net499),
    .D(_01548_),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22082_ (.CLK(net500),
    .D(_01549_),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22083_ (.CLK(net501),
    .D(_01550_),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22084_ (.CLK(net502),
    .D(_01551_),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _22085_ (.CLK(net503),
    .D(_01552_),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22086_ (.CLK(net504),
    .D(_01553_),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22087_ (.CLK(net505),
    .D(_01554_),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22088_ (.CLK(net506),
    .D(_01555_),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _22089_ (.CLK(net507),
    .D(_01556_),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _22090_ (.CLK(net508),
    .D(_01557_),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _22091_ (.CLK(net509),
    .D(_01558_),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _22092_ (.CLK(net510),
    .D(_01559_),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _22093_ (.CLK(net511),
    .D(_01560_),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _22094_ (.CLK(net512),
    .D(_01561_),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _22095_ (.CLK(net513),
    .D(_01562_),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _22096_ (.CLK(net134),
    .D(_01563_),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _22097_ (.CLK(net135),
    .D(_01564_),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _22098_ (.CLK(net136),
    .D(_01565_),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _22099_ (.CLK(net137),
    .D(_01566_),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _22100_ (.CLK(net138),
    .D(_01567_),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _22101_ (.CLK(net139),
    .D(_01568_),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _22102_ (.CLK(net140),
    .D(_01569_),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _22103_ (.CLK(net141),
    .D(_01570_),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _22104_ (.CLK(net142),
    .D(_01571_),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _22105_ (.CLK(net143),
    .D(_01572_),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22106_ (.CLK(net144),
    .D(_01573_),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22107_ (.CLK(net145),
    .D(_01574_),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22108_ (.CLK(net146),
    .D(_01575_),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22109_ (.CLK(net147),
    .D(_01576_),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22110_ (.CLK(net148),
    .D(_01577_),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22111_ (.CLK(net149),
    .D(_01578_),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22112_ (.CLK(net150),
    .D(_01579_),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22113_ (.CLK(net151),
    .D(_01580_),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22114_ (.CLK(net152),
    .D(_01581_),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22115_ (.CLK(net153),
    .D(_01582_),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22116_ (.CLK(net130),
    .D(_01583_),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22117_ (.CLK(net131),
    .D(_01584_),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22118_ (.CLK(net132),
    .D(_01585_),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22119_ (.CLK(net133),
    .D(_01586_),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22120_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01587_),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22121_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01588_),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22122_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01589_),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _22123_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01590_),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _22124_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01591_),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22125_ (.CLK(clknet_leaf_75_i_clk),
    .D(_01592_),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22126_ (.CLK(clknet_leaf_74_i_clk),
    .D(_01593_),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22127_ (.CLK(clknet_leaf_56_i_clk),
    .D(_01594_),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22128_ (.CLK(clknet_leaf_56_i_clk),
    .D(_01595_),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _22129_ (.CLK(clknet_leaf_57_i_clk),
    .D(_01596_),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _22130_ (.CLK(clknet_leaf_57_i_clk),
    .D(_01597_),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _22131_ (.CLK(clknet_leaf_57_i_clk),
    .D(_01598_),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _22132_ (.CLK(clknet_leaf_58_i_clk),
    .D(_01599_),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _22133_ (.CLK(clknet_leaf_58_i_clk),
    .D(_01600_),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22134_ (.CLK(clknet_leaf_61_i_clk),
    .D(_01601_),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22135_ (.CLK(clknet_leaf_61_i_clk),
    .D(_01602_),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22136_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01603_),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22137_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01604_),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22138_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01605_),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22139_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01606_),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22140_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01607_),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22141_ (.CLK(clknet_leaf_56_i_clk),
    .D(_01608_),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22142_ (.CLK(clknet_leaf_56_i_clk),
    .D(_01609_),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22143_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01610_),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_4 _22144_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01611_),
    .Q(\rbzero.trace_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22145_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01612_),
    .Q(\rbzero.trace_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _22146_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01613_),
    .Q(\rbzero.trace_state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _22147_ (.CLK(clknet_leaf_77_i_clk),
    .D(_01614_),
    .Q(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22148_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01615_),
    .Q(\reg_gpout[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22149_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01616_),
    .Q(\reg_gpout[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22150_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01617_),
    .Q(\reg_gpout[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22151_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01618_),
    .Q(\reg_gpout[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22152_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01619_),
    .Q(\reg_gpout[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22153_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01620_),
    .Q(\reg_gpout[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22154_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01621_),
    .Q(reg_hsync));
 sky130_fd_sc_hd__dfxtp_1 _22155_ (.CLK(clknet_leaf_56_i_clk),
    .D(_01622_),
    .Q(reg_vsync));
 sky130_fd_sc_hd__dfxtp_1 _22156_ (.CLK(clknet_leaf_57_i_clk),
    .D(_01623_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22157_ (.CLK(clknet_leaf_61_i_clk),
    .D(_01624_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22158_ (.CLK(clknet_leaf_61_i_clk),
    .D(_01625_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22159_ (.CLK(clknet_leaf_61_i_clk),
    .D(_01626_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22160_ (.CLK(clknet_leaf_60_i_clk),
    .D(_01627_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22161_ (.CLK(clknet_leaf_57_i_clk),
    .D(_01628_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22162_ (.CLK(clknet_leaf_59_i_clk),
    .D(_01629_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22163_ (.CLK(clknet_leaf_56_i_clk),
    .D(_01630_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22164_ (.CLK(clknet_leaf_59_i_clk),
    .D(_01631_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22165_ (.CLK(clknet_leaf_59_i_clk),
    .D(_01632_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22166_ (.CLK(clknet_leaf_59_i_clk),
    .D(_01633_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22167_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01634_),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22168_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01635_),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22169_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01636_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22170_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01637_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22171_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01638_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22172_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01639_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22173_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01640_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22174_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01641_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22175_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01642_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22176_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01643_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22177_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01644_),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22178_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01645_),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22179_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01646_),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22180_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01647_),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22181_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01648_),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22182_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01649_),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22183_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01650_),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22184_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01651_),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_122 (.HI(net122));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_124 (.HI(net124));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_125 (.HI(net125));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_126 (.HI(net126));
 sky130_fd_sc_hd__inv_2 _11494__1 (.A(clknet_leaf_51_i_clk),
    .Y(net127));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.HI(net111));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(i_debug_map_overlay),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(i_debug_trace_overlay),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(i_debug_vec_overlay),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(i_gpout0_sel[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(i_gpout0_sel[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(i_gpout0_sel[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(i_gpout0_sel[3]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(i_gpout0_sel[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(i_gpout0_sel[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(i_gpout1_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__buf_6 input11 (.A(i_gpout1_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(i_gpout1_sel[2]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(i_gpout1_sel[3]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 input14 (.A(i_gpout1_sel[4]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(i_gpout1_sel[5]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(i_gpout2_sel[0]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(i_gpout2_sel[1]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(i_gpout2_sel[2]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(i_gpout2_sel[3]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(i_gpout2_sel[4]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(i_gpout2_sel[5]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(i_gpout3_sel[0]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(i_gpout3_sel[1]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(i_gpout3_sel[2]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(i_gpout3_sel[3]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(i_gpout3_sel[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(i_gpout3_sel[5]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(i_gpout4_sel[0]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(i_gpout4_sel[1]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(i_gpout4_sel[2]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(i_gpout4_sel[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(i_gpout4_sel[4]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(i_gpout4_sel[5]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(i_gpout5_sel[0]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(i_gpout5_sel[1]),
    .X(net35));
 sky130_fd_sc_hd__buf_6 input36 (.A(i_gpout5_sel[2]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(i_gpout5_sel[3]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(i_gpout5_sel[4]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(i_gpout5_sel[5]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_16 input40 (.A(i_mode[0]),
    .X(net40));
 sky130_fd_sc_hd__buf_12 input41 (.A(i_mode[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input42 (.A(i_mode[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(i_reg_csb),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(i_reg_mosi),
    .X(net44));
 sky130_fd_sc_hd__buf_8 input45 (.A(i_reg_outs_enb),
    .X(net45));
 sky130_fd_sc_hd__buf_8 input46 (.A(i_reg_sclk),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(i_reset_lock_a),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(i_reset_lock_b),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(i_test_uc2),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(i_test_wci),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input51 (.A(i_tex_in[0]),
    .X(net51));
 sky130_fd_sc_hd__buf_6 input52 (.A(i_tex_in[1]),
    .X(net52));
 sky130_fd_sc_hd__buf_6 input53 (.A(i_tex_in[2]),
    .X(net53));
 sky130_fd_sc_hd__buf_4 input54 (.A(i_tex_in[3]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(i_vec_csb),
    .X(net55));
 sky130_fd_sc_hd__buf_4 input56 (.A(i_vec_mosi),
    .X(net56));
 sky130_fd_sc_hd__buf_6 input57 (.A(i_vec_sclk),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(o_hsync));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(o_reset));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(o_tex_csb));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(o_tex_out0));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net127),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(o_vsync));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_77 (.LO(net77));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_leaf_38_i_clk),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 net99_3 (.A(clknet_leaf_37_i_clk),
    .Y(net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_opt_6_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_opt_7_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_opt_5_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_opt_2_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_opt_3_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_opt_4_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_leaf_100_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_101_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_leaf_102_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_104_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_leaf_105_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_106_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_107_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_108_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_109_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_111_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_112_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_113_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_114_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_116_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_leaf_117_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_118_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_119_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_120_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_leaf_121_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_122_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_123_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_124_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_125_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_126_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_127_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_128_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_129_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_130_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_131_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_132_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_133_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_134_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_135_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_136_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_leaf_137_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_138_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_139_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_leaf_140_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_141_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_142_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_143_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_leaf_144_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_1_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_2_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_1_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_2_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_1_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_2_2_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_1_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_2_3_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_2_0_1_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_2_0_1_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_2_1_1_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_2_1_1_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_2_2_1_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_2_2_1_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_2_3_1_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_2_3_1_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_opt_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_opt_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_0_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_opt_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_0_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_opt_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_0_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_opt_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_0_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_opt_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_0_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_opt_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05731_ (.A(_05731_),
    .X(clknet_0__05731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05731_ (.A(clknet_0__05731_),
    .X(clknet_1_0__leaf__05731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05731_ (.A(clknet_0__05731_),
    .X(clknet_1_1__leaf__05731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05991_ (.A(_05991_),
    .X(clknet_0__05991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05991_ (.A(clknet_0__05991_),
    .X(clknet_1_0__leaf__05991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05991_ (.A(clknet_0__05991_),
    .X(clknet_1_1__leaf__05991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05762_ (.A(_05762_),
    .X(clknet_0__05762_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05762_ (.A(clknet_0__05762_),
    .X(clknet_1_0__leaf__05762_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05762_ (.A(clknet_0__05762_),
    .X(clknet_1_1__leaf__05762_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03849_ (.A(_03849_),
    .X(clknet_0__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03849_ (.A(clknet_0__03849_),
    .X(clknet_1_0__leaf__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03849_ (.A(clknet_0__03849_),
    .X(clknet_1_1__leaf__03849_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03848_ (.A(_03848_),
    .X(clknet_0__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03848_ (.A(clknet_0__03848_),
    .X(clknet_1_0__leaf__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03848_ (.A(clknet_0__03848_),
    .X(clknet_1_1__leaf__03848_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03837_ (.A(_03837_),
    .X(clknet_0__03837_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03837_ (.A(clknet_0__03837_),
    .X(clknet_1_0__leaf__03837_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03837_ (.A(clknet_0__03837_),
    .X(clknet_1_1__leaf__03837_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03847_ (.A(_03847_),
    .X(clknet_0__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03847_ (.A(clknet_0__03847_),
    .X(clknet_1_0__leaf__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03847_ (.A(clknet_0__03847_),
    .X(clknet_1_1__leaf__03847_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03846_ (.A(_03846_),
    .X(clknet_0__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03846_ (.A(clknet_0__03846_),
    .X(clknet_1_0__leaf__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03846_ (.A(clknet_0__03846_),
    .X(clknet_1_1__leaf__03846_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03845_ (.A(_03845_),
    .X(clknet_0__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03845_ (.A(clknet_0__03845_),
    .X(clknet_1_0__leaf__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03845_ (.A(clknet_0__03845_),
    .X(clknet_1_1__leaf__03845_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03844_ (.A(_03844_),
    .X(clknet_0__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03844_ (.A(clknet_0__03844_),
    .X(clknet_1_0__leaf__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03844_ (.A(clknet_0__03844_),
    .X(clknet_1_1__leaf__03844_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03843_ (.A(_03843_),
    .X(clknet_0__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03843_ (.A(clknet_0__03843_),
    .X(clknet_1_0__leaf__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03843_ (.A(clknet_0__03843_),
    .X(clknet_1_1__leaf__03843_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03842_ (.A(_03842_),
    .X(clknet_0__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03842_ (.A(clknet_0__03842_),
    .X(clknet_1_0__leaf__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03842_ (.A(clknet_0__03842_),
    .X(clknet_1_1__leaf__03842_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03841_ (.A(_03841_),
    .X(clknet_0__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03841_ (.A(clknet_0__03841_),
    .X(clknet_1_0__leaf__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03841_ (.A(clknet_0__03841_),
    .X(clknet_1_1__leaf__03841_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03840_ (.A(_03840_),
    .X(clknet_0__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03840_ (.A(clknet_0__03840_),
    .X(clknet_1_0__leaf__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03840_ (.A(clknet_0__03840_),
    .X(clknet_1_1__leaf__03840_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03839_ (.A(_03839_),
    .X(clknet_0__03839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03839_ (.A(clknet_0__03839_),
    .X(clknet_1_0__leaf__03839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03839_ (.A(clknet_0__03839_),
    .X(clknet_1_1__leaf__03839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03838_ (.A(_03838_),
    .X(clknet_0__03838_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03838_ (.A(clknet_0__03838_),
    .X(clknet_1_0__leaf__03838_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03838_ (.A(clknet_0__03838_),
    .X(clknet_1_1__leaf__03838_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03826_ (.A(_03826_),
    .X(clknet_0__03826_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03826_ (.A(clknet_0__03826_),
    .X(clknet_1_0__leaf__03826_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03826_ (.A(clknet_0__03826_),
    .X(clknet_1_1__leaf__03826_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03836_ (.A(_03836_),
    .X(clknet_0__03836_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03836_ (.A(clknet_0__03836_),
    .X(clknet_1_0__leaf__03836_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03836_ (.A(clknet_0__03836_),
    .X(clknet_1_1__leaf__03836_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03835_ (.A(_03835_),
    .X(clknet_0__03835_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03835_ (.A(clknet_0__03835_),
    .X(clknet_1_0__leaf__03835_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03835_ (.A(clknet_0__03835_),
    .X(clknet_1_1__leaf__03835_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03834_ (.A(_03834_),
    .X(clknet_0__03834_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03834_ (.A(clknet_0__03834_),
    .X(clknet_1_0__leaf__03834_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03834_ (.A(clknet_0__03834_),
    .X(clknet_1_1__leaf__03834_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03833_ (.A(_03833_),
    .X(clknet_0__03833_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03833_ (.A(clknet_0__03833_),
    .X(clknet_1_0__leaf__03833_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03833_ (.A(clknet_0__03833_),
    .X(clknet_1_1__leaf__03833_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03832_ (.A(_03832_),
    .X(clknet_0__03832_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03832_ (.A(clknet_0__03832_),
    .X(clknet_1_0__leaf__03832_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03832_ (.A(clknet_0__03832_),
    .X(clknet_1_1__leaf__03832_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03831_ (.A(_03831_),
    .X(clknet_0__03831_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03831_ (.A(clknet_0__03831_),
    .X(clknet_1_0__leaf__03831_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03831_ (.A(clknet_0__03831_),
    .X(clknet_1_1__leaf__03831_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03830_ (.A(_03830_),
    .X(clknet_0__03830_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03830_ (.A(clknet_0__03830_),
    .X(clknet_1_0__leaf__03830_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03830_ (.A(clknet_0__03830_),
    .X(clknet_1_1__leaf__03830_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03829_ (.A(_03829_),
    .X(clknet_0__03829_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03829_ (.A(clknet_0__03829_),
    .X(clknet_1_0__leaf__03829_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03829_ (.A(clknet_0__03829_),
    .X(clknet_1_1__leaf__03829_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03828_ (.A(_03828_),
    .X(clknet_0__03828_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03828_ (.A(clknet_0__03828_),
    .X(clknet_1_0__leaf__03828_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03828_ (.A(clknet_0__03828_),
    .X(clknet_1_1__leaf__03828_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03827_ (.A(_03827_),
    .X(clknet_0__03827_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03827_ (.A(clknet_0__03827_),
    .X(clknet_1_0__leaf__03827_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03827_ (.A(clknet_0__03827_),
    .X(clknet_1_1__leaf__03827_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03616_ (.A(_03616_),
    .X(clknet_0__03616_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03616_ (.A(clknet_0__03616_),
    .X(clknet_1_0__leaf__03616_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03616_ (.A(clknet_0__03616_),
    .X(clknet_1_1__leaf__03616_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03825_ (.A(_03825_),
    .X(clknet_0__03825_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03825_ (.A(clknet_0__03825_),
    .X(clknet_1_0__leaf__03825_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03825_ (.A(clknet_0__03825_),
    .X(clknet_1_1__leaf__03825_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03824_ (.A(_03824_),
    .X(clknet_0__03824_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03824_ (.A(clknet_0__03824_),
    .X(clknet_1_0__leaf__03824_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03824_ (.A(clknet_0__03824_),
    .X(clknet_1_1__leaf__03824_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03823_ (.A(_03823_),
    .X(clknet_0__03823_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03823_ (.A(clknet_0__03823_),
    .X(clknet_1_0__leaf__03823_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03823_ (.A(clknet_0__03823_),
    .X(clknet_1_1__leaf__03823_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03822_ (.A(_03822_),
    .X(clknet_0__03822_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03822_ (.A(clknet_0__03822_),
    .X(clknet_1_0__leaf__03822_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03822_ (.A(clknet_0__03822_),
    .X(clknet_1_1__leaf__03822_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03821_ (.A(_03821_),
    .X(clknet_0__03821_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03821_ (.A(clknet_0__03821_),
    .X(clknet_1_0__leaf__03821_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03821_ (.A(clknet_0__03821_),
    .X(clknet_1_1__leaf__03821_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03820_ (.A(_03820_),
    .X(clknet_0__03820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03820_ (.A(clknet_0__03820_),
    .X(clknet_1_0__leaf__03820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03820_ (.A(clknet_0__03820_),
    .X(clknet_1_1__leaf__03820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03819_ (.A(_03819_),
    .X(clknet_0__03819_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03819_ (.A(clknet_0__03819_),
    .X(clknet_1_0__leaf__03819_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03819_ (.A(clknet_0__03819_),
    .X(clknet_1_1__leaf__03819_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03818_ (.A(_03818_),
    .X(clknet_0__03818_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03818_ (.A(clknet_0__03818_),
    .X(clknet_1_0__leaf__03818_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03818_ (.A(clknet_0__03818_),
    .X(clknet_1_1__leaf__03818_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03817_ (.A(_03817_),
    .X(clknet_0__03817_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03817_ (.A(clknet_0__03817_),
    .X(clknet_1_0__leaf__03817_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03817_ (.A(clknet_0__03817_),
    .X(clknet_1_1__leaf__03817_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03617_ (.A(_03617_),
    .X(clknet_0__03617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03617_ (.A(clknet_0__03617_),
    .X(clknet_1_0__leaf__03617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03617_ (.A(clknet_0__03617_),
    .X(clknet_1_1__leaf__03617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03609_ (.A(_03609_),
    .X(clknet_0__03609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03609_ (.A(clknet_0__03609_),
    .X(clknet_1_0__leaf__03609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03609_ (.A(clknet_0__03609_),
    .X(clknet_1_1__leaf__03609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03615_ (.A(_03615_),
    .X(clknet_0__03615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03615_ (.A(clknet_0__03615_),
    .X(clknet_1_0__leaf__03615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03615_ (.A(clknet_0__03615_),
    .X(clknet_1_1__leaf__03615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03614_ (.A(_03614_),
    .X(clknet_0__03614_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03614_ (.A(clknet_0__03614_),
    .X(clknet_1_0__leaf__03614_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03614_ (.A(clknet_0__03614_),
    .X(clknet_1_1__leaf__03614_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03613_ (.A(_03613_),
    .X(clknet_0__03613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03613_ (.A(clknet_0__03613_),
    .X(clknet_1_0__leaf__03613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03613_ (.A(clknet_0__03613_),
    .X(clknet_1_1__leaf__03613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03612_ (.A(_03612_),
    .X(clknet_0__03612_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03612_ (.A(clknet_0__03612_),
    .X(clknet_1_0__leaf__03612_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03612_ (.A(clknet_0__03612_),
    .X(clknet_1_1__leaf__03612_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03611_ (.A(_03611_),
    .X(clknet_0__03611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03611_ (.A(clknet_0__03611_),
    .X(clknet_1_0__leaf__03611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03611_ (.A(clknet_0__03611_),
    .X(clknet_1_1__leaf__03611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03610_ (.A(_03610_),
    .X(clknet_0__03610_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03610_ (.A(clknet_0__03610_),
    .X(clknet_1_0__leaf__03610_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03610_ (.A(clknet_0__03610_),
    .X(clknet_1_1__leaf__03610_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05944_ (.A(_05944_),
    .X(clknet_0__05944_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05944_ (.A(clknet_0__05944_),
    .X(clknet_1_0__leaf__05944_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05944_ (.A(clknet_0__05944_),
    .X(clknet_1_1__leaf__05944_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05893_ (.A(_05893_),
    .X(clknet_0__05893_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05893_ (.A(clknet_0__05893_),
    .X(clknet_1_0__leaf__05893_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05893_ (.A(clknet_0__05893_),
    .X(clknet_1_1__leaf__05893_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05839_ (.A(_05839_),
    .X(clknet_0__05839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05839_ (.A(clknet_0__05839_),
    .X(clknet_1_0__leaf__05839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05839_ (.A(clknet_0__05839_),
    .X(clknet_1_1__leaf__05839_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05786_ (.A(_05786_),
    .X(clknet_0__05786_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05786_ (.A(clknet_0__05786_),
    .X(clknet_1_0__leaf__05786_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05786_ (.A(clknet_0__05786_),
    .X(clknet_1_1__leaf__05786_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rbzero.tex_r1[40] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\rbzero.pov.ready_buffer[40] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02653_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_04687_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_04925_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_06155_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_07042_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_08113_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_08120_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_08191_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_08191_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_08219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_08798_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_09221_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_09589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_09702_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_09732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_09784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\rbzero.trace_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_02235_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_04898_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_04982_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_05672_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_06163_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_09570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_09732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_04847_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_05089_));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1163 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1171 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1243 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1250 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1151 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1094 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1245 ();
 assign o_rgb[0] = net77;
 assign o_rgb[10] = net85;
 assign o_rgb[11] = net86;
 assign o_rgb[12] = net87;
 assign o_rgb[13] = net88;
 assign o_rgb[16] = net89;
 assign o_rgb[17] = net90;
 assign o_rgb[18] = net91;
 assign o_rgb[19] = net92;
 assign o_rgb[1] = net78;
 assign o_rgb[20] = net93;
 assign o_rgb[21] = net94;
 assign o_rgb[2] = net79;
 assign o_rgb[3] = net80;
 assign o_rgb[4] = net81;
 assign o_rgb[5] = net82;
 assign o_rgb[8] = net83;
 assign o_rgb[9] = net84;
 assign ones[0] = net111;
 assign ones[10] = net121;
 assign ones[11] = net122;
 assign ones[12] = net123;
 assign ones[13] = net124;
 assign ones[14] = net125;
 assign ones[15] = net126;
 assign ones[1] = net112;
 assign ones[2] = net113;
 assign ones[3] = net114;
 assign ones[4] = net115;
 assign ones[5] = net116;
 assign ones[6] = net117;
 assign ones[7] = net118;
 assign ones[8] = net119;
 assign ones[9] = net120;
 assign zeros[0] = net95;
 assign zeros[10] = net105;
 assign zeros[11] = net106;
 assign zeros[12] = net107;
 assign zeros[13] = net108;
 assign zeros[14] = net109;
 assign zeros[15] = net110;
 assign zeros[1] = net96;
 assign zeros[2] = net97;
 assign zeros[3] = net98;
 assign zeros[4] = net99;
 assign zeros[5] = net100;
 assign zeros[6] = net101;
 assign zeros[7] = net102;
 assign zeros[8] = net103;
 assign zeros[9] = net104;
endmodule

